
module register_file ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8735, n8737, n8739, n8741, n8743, n8745, n8747, n8749, n8751, n8753,
         n8755, n8757, n8759, n8761, n8763, n8765, n8767, n8769, n8771, n8773,
         n8775, n8777, n8779, n8781, n8783, n8785, n8787, n8789, n8791, n8793,
         n8795, n8797, n8799, n8801, n8803, n8805, n8807, n8809, n8811, n8813,
         n8815, n8817, n8819, n8821, n8823, n8825, n8827, n8829, n8831, n8833,
         n8835, n8837, n8839, n8841, n8843, n8845, n8847, n8849, n8851, n8853,
         n8855, n8857, n8859, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8992, n8994, n8996, n8998, n9000, n9002, n9004,
         n9006, n9008, n9010, n9012, n9014, n9016, n9018, n9020, n9022, n9024,
         n9026, n9028, n9030, n9032, n9034, n9036, n9038, n9040, n9042, n9044,
         n9046, n9048, n9050, n9052, n9054, n9056, n9058, n9060, n9062, n9064,
         n9066, n9068, n9070, n9072, n9074, n9076, n9078, n9080, n9082, n9084,
         n9086, n9088, n9090, n9092, n9094, n9096, n9098, n9100, n9102, n9104,
         n9106, n9108, n9110, n9112, n9114, n9116, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n17221, n17224, n17227, n17230, n17233,
         n17236, n17239, n17242, n17245, n17248, n17251, n17254, n17257,
         n17260, n17263, n17266, n17269, n17272, n17275, n17278, n17281,
         n17284, n17287, n17290, n17293, n17296, n17299, n17302, n17305,
         n17308, n17311, n17314, n17317, n17320, n17323, n17326, n17329,
         n17332, n17335, n17338, n17341, n17344, n17347, n17350, n17353,
         n17356, n17359, n17362, n17365, n17368, n17371, n17374, n17377,
         n17380, n17383, n17386, n17389, n17392, n17395, n17398, n17401,
         n17404, n17407, n17410, n17471, n17472, n17474, n17475, n17477,
         n17478, n17480, n17481, n17483, n17484, n17486, n17487, n17489,
         n17490, n17492, n17493, n17495, n17496, n17498, n17499, n17501,
         n17502, n17504, n17505, n17507, n17508, n17510, n17511, n17513,
         n17514, n17516, n17517, n17519, n17520, n17522, n17523, n17525,
         n17526, n17528, n17529, n17531, n17532, n17534, n17535, n17537,
         n17538, n17540, n17541, n17543, n17544, n17546, n17547, n17549,
         n17550, n17552, n17553, n17555, n17556, n17558, n17559, n17561,
         n17562, n17564, n17565, n17567, n17568, n17570, n17571, n17573,
         n17574, n17576, n17577, n17579, n17580, n17582, n17583, n17585,
         n17586, n17588, n17589, n17591, n17592, n17594, n17595, n17597,
         n17598, n17600, n17601, n17603, n17604, n17606, n17607, n17609,
         n17610, n17612, n17613, n17615, n17616, n17618, n17619, n17621,
         n17622, n17624, n17625, n17627, n17628, n17630, n17631, n17633,
         n17634, n17636, n17637, n17639, n17640, n17642, n17643, n17645,
         n17646, n17648, n17649, n17651, n17652, n17654, n17655, n17657,
         n17658, n17660, n17661, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23856, n23858, n23860, n23862, n23864, n23866,
         n23868, n23870, n23872, n23874, n23876, n23878, n23880, n23882,
         n23884, n23886, n23888, n23890, n23892, n23894, n23896, n23898,
         n23900, n23902, n23904, n23906, n23908, n23910, n23912, n23914,
         n23916, n23918, n23920, n23922, n23924, n23926, n23928, n23930,
         n23932, n23934, n23936, n23938, n23940, n23942, n23944, n23946,
         n23948, n23950, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564;

  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6403), .CK(CLK), .Q(n19396), .QN(n9118)
         );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6402), .CK(CLK), .Q(n19397), .QN(n9120)
         );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6401), .CK(CLK), .Q(n19398), .QN(n9122)
         );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6400), .CK(CLK), .Q(n19399), .QN(n9124)
         );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6399), .CK(CLK), .Q(n24331), .QN(n9126)
         );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6398), .CK(CLK), .Q(n24330), .QN(n9128)
         );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6397), .CK(CLK), .Q(n24329), .QN(n9130)
         );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6396), .CK(CLK), .Q(n24328), .QN(n9132)
         );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6395), .CK(CLK), .Q(n24327), .QN(n9134)
         );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6394), .CK(CLK), .Q(n24326), .QN(n9136)
         );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6393), .CK(CLK), .Q(n24325), .QN(n9138)
         );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6392), .CK(CLK), .Q(n24324), .QN(n9140)
         );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6391), .CK(CLK), .Q(n24323), .QN(n9142)
         );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6390), .CK(CLK), .Q(n24322), .QN(n9144)
         );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6389), .CK(CLK), .Q(n24321), .QN(n9146)
         );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6388), .CK(CLK), .Q(n24320), .QN(n9148)
         );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6387), .CK(CLK), .Q(n24319), .QN(n9150)
         );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6386), .CK(CLK), .Q(n24318), .QN(n9152)
         );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6385), .CK(CLK), .Q(n24317), .QN(n9154)
         );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6384), .CK(CLK), .Q(n24316), .QN(n9156)
         );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6383), .CK(CLK), .Q(n24315), .QN(n9158)
         );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6382), .CK(CLK), .Q(n24314), .QN(n9160)
         );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6381), .CK(CLK), .Q(n24313), .QN(n9162)
         );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6380), .CK(CLK), .Q(n24312), .QN(n9164)
         );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6379), .CK(CLK), .Q(n24311), .QN(n9166)
         );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6378), .CK(CLK), .Q(n24310), .QN(n9168)
         );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6377), .CK(CLK), .Q(n24309), .QN(n9170)
         );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6376), .CK(CLK), .Q(n24308), .QN(n9172)
         );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6375), .CK(CLK), .Q(n24307), .QN(n9174)
         );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6374), .CK(CLK), .Q(n24306), .QN(n9176)
         );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6373), .CK(CLK), .Q(n24305), .QN(n9178)
         );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6372), .CK(CLK), .Q(n24304), .QN(n9180)
         );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6371), .CK(CLK), .Q(n24303), .QN(n9182)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6370), .CK(CLK), .Q(n24302), .QN(n9184)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6369), .CK(CLK), .Q(n24301), .QN(n9186)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6368), .CK(CLK), .Q(n24300), .QN(n9188)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6367), .CK(CLK), .Q(n24299), .QN(n9190)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6366), .CK(CLK), .Q(n24298), .QN(n9192)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6365), .CK(CLK), .Q(n24297), .QN(n9194)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6364), .CK(CLK), .Q(n24296), .QN(n9196)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6363), .CK(CLK), .Q(n24295), .QN(n9198)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6362), .CK(CLK), .Q(n24294), .QN(n9200)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6361), .CK(CLK), .Q(n24293), .QN(n9202)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6360), .CK(CLK), .Q(n24292), .QN(n9204)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6359), .CK(CLK), .Q(n24291), .QN(n9206)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6358), .CK(CLK), .Q(n24290), .QN(n9208)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6357), .CK(CLK), .Q(n24289), .QN(n9210)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6356), .CK(CLK), .Q(n24288), .QN(n9212)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6355), .CK(CLK), .Q(n24287), .QN(n9214)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6354), .CK(CLK), .Q(n24286), .QN(n9216)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6353), .CK(CLK), .Q(n24285), .QN(n9218)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6352), .CK(CLK), .Q(n24284), .QN(n9220)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6351), .CK(CLK), .Q(n24283), .QN(n9222)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6350), .CK(CLK), .Q(n24282), .QN(n9224)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6349), .CK(CLK), .Q(n24281), .QN(n9226)
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6348), .CK(CLK), .Q(n24280), .QN(n9228)
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6347), .CK(CLK), .Q(n24279), .QN(n9230)
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6346), .CK(CLK), .Q(n24278), .QN(n9232)
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6345), .CK(CLK), .Q(n24277), .QN(n9234)
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6344), .CK(CLK), .Q(n24276), .QN(n9236)
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6343), .CK(CLK), .Q(n24275), .QN(n9238)
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6342), .CK(CLK), .Q(n24274), .QN(n9240)
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6341), .CK(CLK), .Q(n24273), .QN(n9242)
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6340), .CK(CLK), .Q(n24272), .QN(n9244)
         );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6275), .CK(CLK), .QN(n833) );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6274), .CK(CLK), .QN(n834) );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6273), .CK(CLK), .QN(n835) );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6272), .CK(CLK), .QN(n836) );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6271), .CK(CLK), .QN(n837) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6270), .CK(CLK), .QN(n838) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6269), .CK(CLK), .QN(n839) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6268), .CK(CLK), .QN(n840) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6267), .CK(CLK), .QN(n841) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6266), .CK(CLK), .QN(n842) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6265), .CK(CLK), .QN(n843) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6264), .CK(CLK), .QN(n844) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6263), .CK(CLK), .QN(n845) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6262), .CK(CLK), .QN(n846) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6261), .CK(CLK), .QN(n847) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6260), .CK(CLK), .QN(n848) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6259), .CK(CLK), .QN(n849) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6258), .CK(CLK), .QN(n850) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6257), .CK(CLK), .QN(n851) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6256), .CK(CLK), .QN(n852) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6255), .CK(CLK), .QN(n853) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6254), .CK(CLK), .QN(n854) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6253), .CK(CLK), .QN(n855) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6252), .CK(CLK), .QN(n856) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6251), .CK(CLK), .QN(n857) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6250), .CK(CLK), .QN(n858) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6249), .CK(CLK), .QN(n859) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6248), .CK(CLK), .QN(n860) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6247), .CK(CLK), .QN(n861) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6246), .CK(CLK), .QN(n862) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6245), .CK(CLK), .QN(n863) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6244), .CK(CLK), .QN(n864) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6243), .CK(CLK), .QN(n865) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6242), .CK(CLK), .QN(n866) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6241), .CK(CLK), .QN(n867) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6240), .CK(CLK), .QN(n868) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6239), .CK(CLK), .QN(n869) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6238), .CK(CLK), .QN(n870) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6237), .CK(CLK), .QN(n871) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6236), .CK(CLK), .QN(n872) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6235), .CK(CLK), .QN(n873) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6234), .CK(CLK), .QN(n874) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6233), .CK(CLK), .QN(n875) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6232), .CK(CLK), .QN(n876) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6231), .CK(CLK), .QN(n877) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6230), .CK(CLK), .QN(n878) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6229), .CK(CLK), .QN(n879) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6228), .CK(CLK), .QN(n880) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6227), .CK(CLK), .QN(n881) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6226), .CK(CLK), .QN(n882) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6225), .CK(CLK), .QN(n883) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6224), .CK(CLK), .QN(n884) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6223), .CK(CLK), .QN(n885) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6222), .CK(CLK), .QN(n886) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6221), .CK(CLK), .QN(n887) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6220), .CK(CLK), .QN(n888) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6219), .CK(CLK), .QN(n889) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6218), .CK(CLK), .QN(n890) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6217), .CK(CLK), .QN(n891) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6216), .CK(CLK), .QN(n892) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6215), .CK(CLK), .QN(n893) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6214), .CK(CLK), .QN(n894) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6213), .CK(CLK), .QN(n895) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6212), .CK(CLK), .QN(n896) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n5631), .CK(CLK), .Q(n19588), .QN(n9127)
         );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n5630), .CK(CLK), .Q(n19589), .QN(n9129)
         );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n5629), .CK(CLK), .Q(n19590), .QN(n9131)
         );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n5628), .CK(CLK), .Q(n19591), .QN(n9133)
         );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n5627), .CK(CLK), .Q(n19592), .QN(n9135)
         );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n5626), .CK(CLK), .Q(n19593), .QN(n9137)
         );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n5625), .CK(CLK), .Q(n19594), .QN(n9139)
         );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n5624), .CK(CLK), .Q(n19595), .QN(n9141)
         );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n5623), .CK(CLK), .Q(n19596), .QN(n9143)
         );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n5622), .CK(CLK), .Q(n19597), .QN(n9145)
         );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n5621), .CK(CLK), .Q(n19598), .QN(n9147)
         );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5620), .CK(CLK), .Q(n19599), .QN(n9149)
         );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5619), .CK(CLK), .Q(n19600), .QN(n9151)
         );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5618), .CK(CLK), .Q(n19601), .QN(n9153)
         );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5617), .CK(CLK), .Q(n19602), .QN(n9155)
         );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5616), .CK(CLK), .Q(n19603), .QN(n9157)
         );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5615), .CK(CLK), .Q(n19604), .QN(n9159)
         );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5614), .CK(CLK), .Q(n19605), .QN(n9161)
         );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5613), .CK(CLK), .Q(n19606), .QN(n9163)
         );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5612), .CK(CLK), .Q(n19607), .QN(n9165)
         );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5611), .CK(CLK), .Q(n19608), .QN(n9167)
         );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5610), .CK(CLK), .Q(n19609), .QN(n9169)
         );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5609), .CK(CLK), .Q(n19610), .QN(n9171)
         );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5608), .CK(CLK), .Q(n19611), .QN(n9173)
         );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5607), .CK(CLK), .Q(n19612), .QN(n9175)
         );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5606), .CK(CLK), .Q(n19613), .QN(n9177)
         );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5605), .CK(CLK), .Q(n19614), .QN(n9179)
         );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5604), .CK(CLK), .Q(n19615), .QN(n9181)
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5603), .CK(CLK), .Q(n19616), .QN(n9183)
         );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5602), .CK(CLK), .Q(n19617), .QN(n9185)
         );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5601), .CK(CLK), .Q(n19618), .QN(n9187)
         );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5600), .CK(CLK), .Q(n19619), .QN(n9189)
         );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5599), .CK(CLK), .Q(n19620), .QN(n9191)
         );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5598), .CK(CLK), .Q(n19621), .QN(n9193)
         );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5597), .CK(CLK), .Q(n19622), .QN(n9195)
         );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5596), .CK(CLK), .Q(n19623), .QN(n9197)
         );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5595), .CK(CLK), .Q(n19624), .QN(n9199)
         );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5594), .CK(CLK), .Q(n19625), .QN(n9201)
         );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5593), .CK(CLK), .Q(n19626), .QN(n9203)
         );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5592), .CK(CLK), .Q(n19627), .QN(n9205)
         );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5591), .CK(CLK), .Q(n19628), .QN(n9207)
         );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5590), .CK(CLK), .Q(n19629), .QN(n9209)
         );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5589), .CK(CLK), .Q(n19630), .QN(n9211)
         );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5588), .CK(CLK), .Q(n19631), .QN(n9213)
         );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5587), .CK(CLK), .Q(n19632), .QN(n9215)
         );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5586), .CK(CLK), .Q(n19633), .QN(n9217)
         );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5585), .CK(CLK), .Q(n19634), .QN(n9219)
         );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5584), .CK(CLK), .Q(n19635), .QN(n9221)
         );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5583), .CK(CLK), .Q(n19636), .QN(n9223)
         );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5582), .CK(CLK), .Q(n19637), .QN(n9225)
         );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5581), .CK(CLK), .Q(n19638), .QN(n9227)
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5580), .CK(CLK), .Q(n19639), .QN(n9229)
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5579), .CK(CLK), .Q(n19640), .QN(n9231)
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5578), .CK(CLK), .Q(n19641), .QN(n9233)
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5577), .CK(CLK), .Q(n19642), .QN(n9235)
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5576), .CK(CLK), .Q(n19643), .QN(n9237)
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5575), .CK(CLK), .Q(n19644), .QN(n9239)
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5574), .CK(CLK), .Q(n19645), .QN(n9241)
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5573), .CK(CLK), .Q(n19646), .QN(n9243)
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5572), .CK(CLK), .Q(n19647), .QN(n9245)
         );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5506), .CK(CLK), .QN(n7303) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5505), .CK(CLK), .QN(n7305) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5504), .CK(CLK), .QN(n7307) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5503), .CK(CLK), .QN(n7309) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5502), .CK(CLK), .QN(n7311) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5501), .CK(CLK), .QN(n7313) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5500), .CK(CLK), .QN(n7315) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5499), .CK(CLK), .QN(n7317) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5498), .CK(CLK), .QN(n7319) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5497), .CK(CLK), .QN(n7321) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5496), .CK(CLK), .QN(n7323) );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5495), .CK(CLK), .QN(n7325) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5494), .CK(CLK), .QN(n7327) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5493), .CK(CLK), .QN(n7329) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5492), .CK(CLK), .QN(n7331) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5491), .CK(CLK), .QN(n7333) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5490), .CK(CLK), .QN(n7335) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5489), .CK(CLK), .QN(n7337) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5488), .CK(CLK), .QN(n7339) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5487), .CK(CLK), .QN(n7341) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5486), .CK(CLK), .QN(n7343) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5485), .CK(CLK), .QN(n7345) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5484), .CK(CLK), .QN(n7347) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5483), .CK(CLK), .QN(n7349) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5482), .CK(CLK), .QN(n7351) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5481), .CK(CLK), .QN(n7353) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5480), .CK(CLK), .QN(n7355) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5479), .CK(CLK), .QN(n7357) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5478), .CK(CLK), .QN(n7359) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5477), .CK(CLK), .QN(n7361) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5476), .CK(CLK), .QN(n7363) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5475), .CK(CLK), .QN(n7365) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5474), .CK(CLK), .QN(n7367) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5473), .CK(CLK), .QN(n7369) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5472), .CK(CLK), .QN(n7371) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5471), .CK(CLK), .QN(n7373) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5470), .CK(CLK), .QN(n7375) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5469), .CK(CLK), .QN(n7377) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5468), .CK(CLK), .QN(n7379) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5467), .CK(CLK), .QN(n7381) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5466), .CK(CLK), .QN(n7383) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5465), .CK(CLK), .QN(n7385) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5464), .CK(CLK), .QN(n7387) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5463), .CK(CLK), .QN(n7389) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5462), .CK(CLK), .QN(n7391) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5461), .CK(CLK), .QN(n7393) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5460), .CK(CLK), .QN(n7395) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5459), .CK(CLK), .QN(n7397) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5458), .CK(CLK), .QN(n7399) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5457), .CK(CLK), .QN(n7401) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5456), .CK(CLK), .QN(n7403) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5455), .CK(CLK), .QN(n7405) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5454), .CK(CLK), .QN(n7407) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5453), .CK(CLK), .QN(n7409) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5452), .CK(CLK), .QN(n7411) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5451), .CK(CLK), .QN(n7413) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5450), .CK(CLK), .QN(n7415) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5449), .CK(CLK), .QN(n7417) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5448), .CK(CLK), .QN(n7419) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5447), .CK(CLK), .QN(n7421) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5446), .CK(CLK), .QN(n7423) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5445), .CK(CLK), .QN(n7425) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5444), .CK(CLK), .QN(n7427) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5251), .CK(CLK), .Q(n24355), .QN(n8862)
         );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5250), .CK(CLK), .Q(n24354), .QN(n8864)
         );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5249), .CK(CLK), .Q(n24353), .QN(n8866)
         );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5248), .CK(CLK), .Q(n24352), .QN(n8868)
         );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5247), .CK(CLK), .Q(n24351), .QN(n8870)
         );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5246), .CK(CLK), .Q(n24350), .QN(n8872)
         );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5245), .CK(CLK), .Q(n24349), .QN(n8874)
         );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5244), .CK(CLK), .Q(n24348), .QN(n8876)
         );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5243), .CK(CLK), .Q(n24347), .QN(n8878)
         );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5242), .CK(CLK), .Q(n24346), .QN(n8880)
         );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5241), .CK(CLK), .Q(n24345), .QN(n8882)
         );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5240), .CK(CLK), .Q(n24344), .QN(n8884)
         );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5239), .CK(CLK), .Q(n24343), .QN(n8886)
         );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5238), .CK(CLK), .Q(n24342), .QN(n8888)
         );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5237), .CK(CLK), .Q(n24341), .QN(n8890)
         );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5236), .CK(CLK), .Q(n24340), .QN(n8892)
         );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5235), .CK(CLK), .Q(n24339), .QN(n8894)
         );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5234), .CK(CLK), .Q(n24338), .QN(n8896)
         );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5233), .CK(CLK), .Q(n24337), .QN(n8898)
         );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5232), .CK(CLK), .Q(n24336), .QN(n8900)
         );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5231), .CK(CLK), .Q(n24335), .QN(n8902)
         );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5230), .CK(CLK), .Q(n24334), .QN(n8904)
         );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5229), .CK(CLK), .Q(n24333), .QN(n8906)
         );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5228), .CK(CLK), .Q(n24332), .QN(n8908)
         );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5227), .CK(CLK), .Q(n24395), .QN(n8910)
         );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5226), .CK(CLK), .Q(n24394), .QN(n8912)
         );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5225), .CK(CLK), .Q(n24393), .QN(n8914)
         );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5224), .CK(CLK), .Q(n24392), .QN(n8916)
         );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5223), .CK(CLK), .Q(n24391), .QN(n8918)
         );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5222), .CK(CLK), .Q(n24390), .QN(n8920)
         );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5221), .CK(CLK), .Q(n24389), .QN(n8922)
         );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5220), .CK(CLK), .Q(n24388), .QN(n8924)
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5219), .CK(CLK), .Q(n24387), .QN(n8926)
         );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5218), .CK(CLK), .Q(n24386), .QN(n8928)
         );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5217), .CK(CLK), .Q(n24385), .QN(n8930)
         );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5216), .CK(CLK), .Q(n24384), .QN(n8932)
         );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5215), .CK(CLK), .Q(n24383), .QN(n8934)
         );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5214), .CK(CLK), .Q(n24382), .QN(n8936)
         );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5213), .CK(CLK), .Q(n24381), .QN(n8938)
         );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5212), .CK(CLK), .Q(n24380), .QN(n8940)
         );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5211), .CK(CLK), .Q(n24379), .QN(n8942)
         );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5210), .CK(CLK), .Q(n24378), .QN(n8944)
         );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5209), .CK(CLK), .Q(n24377), .QN(n8946)
         );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5208), .CK(CLK), .Q(n24376), .QN(n8948)
         );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5207), .CK(CLK), .Q(n24375), .QN(n8950)
         );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5206), .CK(CLK), .Q(n24374), .QN(n8952)
         );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5205), .CK(CLK), .Q(n24373), .QN(n8954)
         );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5204), .CK(CLK), .Q(n24372), .QN(n8956)
         );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5203), .CK(CLK), .Q(n24371), .QN(n8958)
         );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5202), .CK(CLK), .Q(n24370), .QN(n8960)
         );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5201), .CK(CLK), .Q(n24369), .QN(n8962)
         );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5200), .CK(CLK), .Q(n24368), .QN(n8964)
         );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5199), .CK(CLK), .Q(n24367), .QN(n8966)
         );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5198), .CK(CLK), .Q(n24366), .QN(n8968)
         );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5197), .CK(CLK), .Q(n24365), .QN(n8970)
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5196), .CK(CLK), .Q(n24364), .QN(n8972)
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5195), .CK(CLK), .Q(n24363), .QN(n8974)
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5194), .CK(CLK), .Q(n24362), .QN(n8976)
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5193), .CK(CLK), .Q(n24361), .QN(n8978)
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5192), .CK(CLK), .Q(n24360), .QN(n8980)
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5191), .CK(CLK), .Q(n24359), .QN(n8982)
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5190), .CK(CLK), .Q(n24358), .QN(n8984)
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5189), .CK(CLK), .Q(n24357), .QN(n8986)
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5188), .CK(CLK), .Q(n24356), .QN(n8988)
         );
  DFF_X1 \OUT1_reg[63]  ( .D(n5059), .CK(CLK), .Q(OUT1[63]), .QN(n11846) );
  DFF_X1 \OUT1_reg[62]  ( .D(n5058), .CK(CLK), .Q(OUT1[62]), .QN(n11845) );
  DFF_X1 \OUT1_reg[61]  ( .D(n5057), .CK(CLK), .Q(OUT1[61]), .QN(n11844) );
  DFF_X1 \OUT1_reg[60]  ( .D(n5056), .CK(CLK), .Q(OUT1[60]), .QN(n11843) );
  DFF_X1 \OUT1_reg[59]  ( .D(n5055), .CK(CLK), .Q(OUT1[59]), .QN(n11842) );
  DFF_X1 \OUT1_reg[58]  ( .D(n5054), .CK(CLK), .Q(OUT1[58]), .QN(n11841) );
  DFF_X1 \OUT1_reg[57]  ( .D(n5053), .CK(CLK), .Q(OUT1[57]), .QN(n11840) );
  DFF_X1 \OUT1_reg[56]  ( .D(n5052), .CK(CLK), .Q(OUT1[56]), .QN(n11839) );
  DFF_X1 \OUT1_reg[55]  ( .D(n5051), .CK(CLK), .Q(OUT1[55]), .QN(n11838) );
  DFF_X1 \OUT1_reg[54]  ( .D(n5050), .CK(CLK), .Q(OUT1[54]), .QN(n11837) );
  DFF_X1 \OUT1_reg[53]  ( .D(n5049), .CK(CLK), .Q(OUT1[53]), .QN(n11836) );
  DFF_X1 \OUT1_reg[52]  ( .D(n5048), .CK(CLK), .Q(OUT1[52]), .QN(n11835) );
  DFF_X1 \OUT1_reg[51]  ( .D(n5047), .CK(CLK), .Q(OUT1[51]), .QN(n11834) );
  DFF_X1 \OUT1_reg[50]  ( .D(n5046), .CK(CLK), .Q(OUT1[50]), .QN(n11833) );
  DFF_X1 \OUT1_reg[49]  ( .D(n5045), .CK(CLK), .Q(OUT1[49]), .QN(n11832) );
  DFF_X1 \OUT1_reg[48]  ( .D(n5044), .CK(CLK), .Q(OUT1[48]), .QN(n11831) );
  DFF_X1 \OUT1_reg[47]  ( .D(n5043), .CK(CLK), .Q(OUT1[47]), .QN(n11830) );
  DFF_X1 \OUT1_reg[46]  ( .D(n5042), .CK(CLK), .Q(OUT1[46]), .QN(n11829) );
  DFF_X1 \OUT1_reg[45]  ( .D(n5041), .CK(CLK), .Q(OUT1[45]), .QN(n11828) );
  DFF_X1 \OUT1_reg[44]  ( .D(n5040), .CK(CLK), .Q(OUT1[44]), .QN(n11827) );
  DFF_X1 \OUT1_reg[43]  ( .D(n5039), .CK(CLK), .Q(OUT1[43]), .QN(n11826) );
  DFF_X1 \OUT1_reg[42]  ( .D(n5038), .CK(CLK), .Q(OUT1[42]), .QN(n11825) );
  DFF_X1 \OUT1_reg[41]  ( .D(n5037), .CK(CLK), .Q(OUT1[41]), .QN(n11824) );
  DFF_X1 \OUT1_reg[40]  ( .D(n5036), .CK(CLK), .Q(OUT1[40]), .QN(n11823) );
  DFF_X1 \OUT1_reg[39]  ( .D(n5035), .CK(CLK), .Q(OUT1[39]), .QN(n11822) );
  DFF_X1 \OUT1_reg[38]  ( .D(n5034), .CK(CLK), .Q(OUT1[38]), .QN(n11821) );
  DFF_X1 \OUT1_reg[37]  ( .D(n5033), .CK(CLK), .Q(OUT1[37]), .QN(n11820) );
  DFF_X1 \OUT1_reg[36]  ( .D(n5032), .CK(CLK), .Q(OUT1[36]), .QN(n11819) );
  DFF_X1 \OUT1_reg[35]  ( .D(n5031), .CK(CLK), .Q(OUT1[35]), .QN(n11818) );
  DFF_X1 \OUT1_reg[34]  ( .D(n5030), .CK(CLK), .Q(OUT1[34]), .QN(n11817) );
  DFF_X1 \OUT1_reg[33]  ( .D(n5029), .CK(CLK), .Q(OUT1[33]), .QN(n11816) );
  DFF_X1 \OUT1_reg[32]  ( .D(n5028), .CK(CLK), .Q(OUT1[32]), .QN(n11815) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5027), .CK(CLK), .Q(OUT1[31]), .QN(n11814) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5026), .CK(CLK), .Q(OUT1[30]), .QN(n11813) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5025), .CK(CLK), .Q(OUT1[29]), .QN(n11812) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5024), .CK(CLK), .Q(OUT1[28]), .QN(n11811) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5023), .CK(CLK), .Q(OUT1[27]), .QN(n11810) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5022), .CK(CLK), .Q(OUT1[26]), .QN(n11809) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5021), .CK(CLK), .Q(OUT1[25]), .QN(n11808) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5020), .CK(CLK), .Q(OUT1[24]), .QN(n11807) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5019), .CK(CLK), .Q(OUT1[23]), .QN(n11806) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5018), .CK(CLK), .Q(OUT1[22]), .QN(n11805) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5017), .CK(CLK), .Q(OUT1[21]), .QN(n11804) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5016), .CK(CLK), .Q(OUT1[20]), .QN(n11803) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5015), .CK(CLK), .Q(OUT1[19]), .QN(n11802) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5014), .CK(CLK), .Q(OUT1[18]), .QN(n11801) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5013), .CK(CLK), .Q(OUT1[17]), .QN(n11800) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5012), .CK(CLK), .Q(OUT1[16]), .QN(n11799) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5011), .CK(CLK), .Q(OUT1[15]), .QN(n11798) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5010), .CK(CLK), .Q(OUT1[14]), .QN(n11797) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5009), .CK(CLK), .Q(OUT1[13]), .QN(n11796) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5008), .CK(CLK), .Q(OUT1[12]), .QN(n11795) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5007), .CK(CLK), .Q(OUT1[11]), .QN(n11794) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5006), .CK(CLK), .Q(OUT1[10]), .QN(n11793) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5005), .CK(CLK), .Q(OUT1[9]), .QN(n11792) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5004), .CK(CLK), .Q(OUT1[8]), .QN(n11791) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5003), .CK(CLK), .Q(OUT1[7]), .QN(n11790) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5002), .CK(CLK), .Q(OUT1[6]), .QN(n11789) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5001), .CK(CLK), .Q(OUT1[5]), .QN(n11788) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5000), .CK(CLK), .Q(OUT1[4]), .QN(n11787) );
  DFF_X1 \OUT1_reg[3]  ( .D(n4999), .CK(CLK), .Q(OUT1[3]), .QN(n11786) );
  DFF_X1 \OUT1_reg[2]  ( .D(n4998), .CK(CLK), .Q(OUT1[2]), .QN(n11785) );
  DFF_X1 \OUT1_reg[1]  ( .D(n4997), .CK(CLK), .Q(OUT1[1]), .QN(n11784) );
  DFF_X1 \OUT1_reg[0]  ( .D(n4996), .CK(CLK), .Q(OUT1[0]), .QN(n11783) );
  DFF_X1 \OUT2_reg[39]  ( .D(n4971), .CK(CLK), .Q(OUT2[39]) );
  DFF_X1 \OUT2_reg[38]  ( .D(n4970), .CK(CLK), .Q(OUT2[38]) );
  DFF_X1 \OUT2_reg[37]  ( .D(n4969), .CK(CLK), .Q(OUT2[37]) );
  DFF_X1 \OUT2_reg[36]  ( .D(n4968), .CK(CLK), .Q(OUT2[36]) );
  DFF_X1 \OUT2_reg[35]  ( .D(n4967), .CK(CLK), .Q(OUT2[35]) );
  DFF_X1 \OUT2_reg[34]  ( .D(n4966), .CK(CLK), .Q(OUT2[34]) );
  DFF_X1 \OUT2_reg[33]  ( .D(n4965), .CK(CLK), .Q(OUT2[33]) );
  DFF_X1 \OUT2_reg[32]  ( .D(n4964), .CK(CLK), .Q(OUT2[32]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n4963), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n4962), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n4961), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n4960), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n4959), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n4958), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n4957), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n4956), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n4955), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n4954), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n4953), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n4952), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n4951), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n4950), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n4949), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n4948), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n4947), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n4946), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n4945), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n4944), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n4943), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n4942), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n4941), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n4940), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n4939), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n4938), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n4937), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n4936), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n4935), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n4934), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n4933), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n4932), .CK(CLK), .Q(OUT2[0]) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n5891), .CK(CLK), .Q(n19802), .QN(n8863)
         );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n5890), .CK(CLK), .Q(n19803), .QN(n8865)
         );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n5889), .CK(CLK), .Q(n19804), .QN(n8867)
         );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n5888), .CK(CLK), .Q(n19805), .QN(n8869)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6147), .CK(CLK), .Q(n19810), .QN(n7300)
         );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6146), .CK(CLK), .Q(n19811), .QN(n7302)
         );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6145), .CK(CLK), .Q(n19812), .QN(n7304)
         );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6144), .CK(CLK), .Q(n19813), .QN(n7306)
         );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6467), .CK(CLK), .Q(n19814), .QN(n7428)
         );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6466), .CK(CLK), .Q(n19815), .QN(n7430)
         );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6465), .CK(CLK), .Q(n19816), .QN(n7432)
         );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6464), .CK(CLK), .Q(n19817), .QN(n7434)
         );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n6787), .CK(CLK), .Q(n24211), .QN(n17221)
         );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n6786), .CK(CLK), .Q(n24210), .QN(n17224)
         );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n6785), .CK(CLK), .Q(n24209), .QN(n17227)
         );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n6784), .CK(CLK), .Q(n24208), .QN(n17230)
         );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n5887), .CK(CLK), .Q(n19822), .QN(n8871)
         );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n5886), .CK(CLK), .Q(n19823), .QN(n8873)
         );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n5885), .CK(CLK), .Q(n19824), .QN(n8875)
         );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n5884), .CK(CLK), .Q(n19825), .QN(n8877)
         );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n5883), .CK(CLK), .Q(n19826), .QN(n8879)
         );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n5882), .CK(CLK), .Q(n19827), .QN(n8881)
         );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n5881), .CK(CLK), .Q(n19828), .QN(n8883)
         );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n5880), .CK(CLK), .Q(n19829), .QN(n8885)
         );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n5879), .CK(CLK), .Q(n19830), .QN(n8887)
         );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n5878), .CK(CLK), .Q(n19831), .QN(n8889)
         );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n5877), .CK(CLK), .Q(n19832), .QN(n8891)
         );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n5876), .CK(CLK), .Q(n19833), .QN(n8893)
         );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n5875), .CK(CLK), .Q(n19834), .QN(n8895)
         );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n5874), .CK(CLK), .Q(n19835), .QN(n8897)
         );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n5873), .CK(CLK), .Q(n19836), .QN(n8899)
         );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n5872), .CK(CLK), .Q(n19837), .QN(n8901)
         );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n5871), .CK(CLK), .Q(n19838), .QN(n8903)
         );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n5870), .CK(CLK), .Q(n19839), .QN(n8905)
         );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n5869), .CK(CLK), .Q(n19840), .QN(n8907)
         );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n5868), .CK(CLK), .Q(n19841), .QN(n8909)
         );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n5867), .CK(CLK), .Q(n19842), .QN(n8911)
         );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n5866), .CK(CLK), .Q(n19843), .QN(n8913)
         );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n5865), .CK(CLK), .Q(n19844), .QN(n8915)
         );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n5864), .CK(CLK), .Q(n19845), .QN(n8917)
         );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n5863), .CK(CLK), .Q(n19846), .QN(n8919)
         );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n5862), .CK(CLK), .Q(n19847), .QN(n8921)
         );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n5861), .CK(CLK), .Q(n19848), .QN(n8923)
         );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n5860), .CK(CLK), .Q(n19849), .QN(n8925)
         );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n5859), .CK(CLK), .Q(n19850), .QN(n8927)
         );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n5858), .CK(CLK), .Q(n19851), .QN(n8929)
         );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n5857), .CK(CLK), .Q(n19852), .QN(n8931)
         );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n5856), .CK(CLK), .Q(n19853), .QN(n8933)
         );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n5855), .CK(CLK), .Q(n19854), .QN(n8935)
         );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n5854), .CK(CLK), .Q(n19855), .QN(n8937)
         );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n5853), .CK(CLK), .Q(n19856), .QN(n8939)
         );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n5852), .CK(CLK), .Q(n19857), .QN(n8941)
         );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6143), .CK(CLK), .Q(n19894), .QN(n7308)
         );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6142), .CK(CLK), .Q(n19895), .QN(n7310)
         );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6141), .CK(CLK), .Q(n19896), .QN(n7312)
         );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6140), .CK(CLK), .Q(n19897), .QN(n7314)
         );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6139), .CK(CLK), .Q(n19898), .QN(n7316)
         );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6138), .CK(CLK), .Q(n19899), .QN(n7318)
         );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6137), .CK(CLK), .Q(n19900), .QN(n7320)
         );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6136), .CK(CLK), .Q(n19901), .QN(n7322)
         );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6135), .CK(CLK), .Q(n19902), .QN(n7324)
         );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6134), .CK(CLK), .Q(n19903), .QN(n7326)
         );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6133), .CK(CLK), .Q(n19904), .QN(n7328)
         );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6132), .CK(CLK), .Q(n19905), .QN(n7330)
         );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6131), .CK(CLK), .Q(n19906), .QN(n7332)
         );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6130), .CK(CLK), .Q(n19907), .QN(n7334)
         );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6129), .CK(CLK), .Q(n19908), .QN(n7336)
         );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6128), .CK(CLK), .Q(n19909), .QN(n7338)
         );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6127), .CK(CLK), .Q(n19910), .QN(n7340)
         );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6126), .CK(CLK), .Q(n19911), .QN(n7342)
         );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6125), .CK(CLK), .Q(n19912), .QN(n7344)
         );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6124), .CK(CLK), .Q(n19913), .QN(n7346)
         );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6123), .CK(CLK), .Q(n19914), .QN(n7348)
         );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6122), .CK(CLK), .Q(n19915), .QN(n7350)
         );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6121), .CK(CLK), .Q(n19916), .QN(n7352)
         );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6120), .CK(CLK), .Q(n19917), .QN(n7354)
         );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6119), .CK(CLK), .Q(n19918), .QN(n7356)
         );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6118), .CK(CLK), .Q(n19919), .QN(n7358)
         );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6117), .CK(CLK), .Q(n19920), .QN(n7360)
         );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6116), .CK(CLK), .Q(n19921), .QN(n7362)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6115), .CK(CLK), .Q(n19922), .QN(n7364)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6114), .CK(CLK), .Q(n19923), .QN(n7366)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6113), .CK(CLK), .Q(n19924), .QN(n7368)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6112), .CK(CLK), .Q(n19925), .QN(n7370)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6111), .CK(CLK), .Q(n19926), .QN(n7372)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6110), .CK(CLK), .Q(n19927), .QN(n7374)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6109), .CK(CLK), .Q(n19928), .QN(n7376)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6108), .CK(CLK), .Q(n19929), .QN(n7378)
         );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6463), .CK(CLK), .Q(n24207), .QN(n7436)
         );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6462), .CK(CLK), .Q(n24206), .QN(n7438)
         );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6461), .CK(CLK), .Q(n24205), .QN(n7440)
         );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6460), .CK(CLK), .Q(n24204), .QN(n7442)
         );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6459), .CK(CLK), .Q(n24203), .QN(n7444)
         );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6458), .CK(CLK), .Q(n24202), .QN(n7446)
         );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6457), .CK(CLK), .Q(n24201), .QN(n7448)
         );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6456), .CK(CLK), .Q(n24200), .QN(n7450)
         );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6455), .CK(CLK), .Q(n24199), .QN(n7452)
         );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6454), .CK(CLK), .Q(n24198), .QN(n7454)
         );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6453), .CK(CLK), .Q(n24197), .QN(n7456)
         );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6452), .CK(CLK), .Q(n24196), .QN(n7458)
         );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6451), .CK(CLK), .Q(n24195), .QN(n7460)
         );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6450), .CK(CLK), .Q(n24194), .QN(n7462)
         );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6449), .CK(CLK), .Q(n24193), .QN(n7464)
         );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6448), .CK(CLK), .Q(n24192), .QN(n7466)
         );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6447), .CK(CLK), .Q(n24191), .QN(n7468)
         );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6446), .CK(CLK), .Q(n24190), .QN(n7470)
         );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6445), .CK(CLK), .Q(n24189), .QN(n7472)
         );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6444), .CK(CLK), .Q(n24188), .QN(n7474)
         );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6443), .CK(CLK), .Q(n24187), .QN(n7476)
         );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6442), .CK(CLK), .Q(n24186), .QN(n7478)
         );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6441), .CK(CLK), .Q(n24185), .QN(n7480)
         );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6440), .CK(CLK), .Q(n24184), .QN(n7482)
         );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6439), .CK(CLK), .Q(n24183), .QN(n7484)
         );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6438), .CK(CLK), .Q(n24182), .QN(n7486)
         );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6437), .CK(CLK), .Q(n24181), .QN(n7488)
         );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6436), .CK(CLK), .Q(n24180), .QN(n7490)
         );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6435), .CK(CLK), .Q(n24179), .QN(n7492)
         );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6434), .CK(CLK), .Q(n24178), .QN(n7494)
         );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6433), .CK(CLK), .Q(n24177), .QN(n7496)
         );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6432), .CK(CLK), .Q(n24176), .QN(n7498)
         );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6431), .CK(CLK), .Q(n24175), .QN(n7500)
         );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6430), .CK(CLK), .Q(n24174), .QN(n7502)
         );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6429), .CK(CLK), .Q(n24173), .QN(n7504)
         );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6428), .CK(CLK), .Q(n24172), .QN(n7506)
         );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n6783), .CK(CLK), .Q(n24271), .QN(n17233)
         );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n6782), .CK(CLK), .Q(n24270), .QN(n17236)
         );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n6781), .CK(CLK), .Q(n24269), .QN(n17239)
         );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n6780), .CK(CLK), .Q(n24268), .QN(n17242)
         );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n6779), .CK(CLK), .Q(n24267), .QN(n17245)
         );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n6778), .CK(CLK), .Q(n24266), .QN(n17248)
         );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n6777), .CK(CLK), .Q(n24265), .QN(n17251)
         );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n6776), .CK(CLK), .Q(n24264), .QN(n17254)
         );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n6775), .CK(CLK), .Q(n24263), .QN(n17257)
         );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n6774), .CK(CLK), .Q(n24262), .QN(n17260)
         );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n6773), .CK(CLK), .Q(n24261), .QN(n17263)
         );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n6772), .CK(CLK), .Q(n24260), .QN(n17266)
         );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n6771), .CK(CLK), .Q(n24259), .QN(n17269)
         );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n6770), .CK(CLK), .Q(n24258), .QN(n17272)
         );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n6769), .CK(CLK), .Q(n24257), .QN(n17275)
         );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n6768), .CK(CLK), .Q(n24256), .QN(n17278)
         );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n6767), .CK(CLK), .Q(n24255), .QN(n17281)
         );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n6766), .CK(CLK), .Q(n24254), .QN(n17284)
         );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n6765), .CK(CLK), .Q(n24253), .QN(n17287)
         );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n6764), .CK(CLK), .Q(n24252), .QN(n17290)
         );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n6763), .CK(CLK), .Q(n24251), .QN(n17293)
         );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n6762), .CK(CLK), .Q(n24250), .QN(n17296)
         );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n6761), .CK(CLK), .Q(n24249), .QN(n17299)
         );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n6760), .CK(CLK), .Q(n24248), .QN(n17302)
         );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n6759), .CK(CLK), .Q(n24247), .QN(n17305)
         );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n6758), .CK(CLK), .Q(n24246), .QN(n17308)
         );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n6757), .CK(CLK), .Q(n24245), .QN(n17311)
         );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n6756), .CK(CLK), .Q(n24244), .QN(n17314)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n6755), .CK(CLK), .Q(n24243), .QN(n17317)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n6754), .CK(CLK), .Q(n24242), .QN(n17320)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n6753), .CK(CLK), .Q(n24241), .QN(n17323)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n6752), .CK(CLK), .Q(n24240), .QN(n17326)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n6751), .CK(CLK), .Q(n24239), .QN(n17329)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n6750), .CK(CLK), .Q(n24238), .QN(n17332)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n6749), .CK(CLK), .Q(n24237), .QN(n17335)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n6748), .CK(CLK), .Q(n24236), .QN(n17338)
         );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n5851), .CK(CLK), .Q(n20002), .QN(n8943)
         );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n5850), .CK(CLK), .Q(n20003), .QN(n8945)
         );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n5849), .CK(CLK), .Q(n20004), .QN(n8947)
         );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n5848), .CK(CLK), .Q(n20005), .QN(n8949)
         );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n5847), .CK(CLK), .Q(n20006), .QN(n8951)
         );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n5846), .CK(CLK), .Q(n20007), .QN(n8953)
         );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n5845), .CK(CLK), .Q(n20008), .QN(n8955)
         );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n5844), .CK(CLK), .Q(n20009), .QN(n8957)
         );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n5843), .CK(CLK), .Q(n20010), .QN(n8959)
         );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n5842), .CK(CLK), .Q(n20011), .QN(n8961)
         );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n5841), .CK(CLK), .Q(n20012), .QN(n8963)
         );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n5840), .CK(CLK), .Q(n20013), .QN(n8965)
         );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n5839), .CK(CLK), .Q(n20014), .QN(n8967)
         );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n5838), .CK(CLK), .Q(n20015), .QN(n8969)
         );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n5837), .CK(CLK), .Q(n20016), .QN(n8971)
         );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n5836), .CK(CLK), .Q(n20017), .QN(n8973)
         );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n5835), .CK(CLK), .Q(n20018), .QN(n8975)
         );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n5834), .CK(CLK), .Q(n20019), .QN(n8977)
         );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n5833), .CK(CLK), .Q(n20020), .QN(n8979)
         );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n5832), .CK(CLK), .Q(n20021), .QN(n8981)
         );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n5831), .CK(CLK), .Q(n20022), .QN(n8983)
         );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n5830), .CK(CLK), .Q(n20023), .QN(n8985)
         );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n5829), .CK(CLK), .Q(n20024), .QN(n8987)
         );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n5828), .CK(CLK), .Q(n20025), .QN(n8989)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6107), .CK(CLK), .Q(n20050), .QN(n7380)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6106), .CK(CLK), .Q(n20051), .QN(n7382)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6105), .CK(CLK), .Q(n20052), .QN(n7384)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6104), .CK(CLK), .Q(n20053), .QN(n7386)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6103), .CK(CLK), .Q(n20054), .QN(n7388)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6102), .CK(CLK), .Q(n20055), .QN(n7390)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6101), .CK(CLK), .Q(n20056), .QN(n7392)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6100), .CK(CLK), .Q(n20057), .QN(n7394)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6099), .CK(CLK), .Q(n20058), .QN(n7396)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6098), .CK(CLK), .Q(n20059), .QN(n7398)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6097), .CK(CLK), .Q(n20060), .QN(n7400)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6096), .CK(CLK), .Q(n20061), .QN(n7402)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6095), .CK(CLK), .Q(n20062), .QN(n7404)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6094), .CK(CLK), .Q(n20063), .QN(n7406)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6093), .CK(CLK), .Q(n20064), .QN(n7408)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6092), .CK(CLK), .Q(n20065), .QN(n7410)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6091), .CK(CLK), .Q(n20066), .QN(n7412)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6090), .CK(CLK), .Q(n20067), .QN(n7414)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6089), .CK(CLK), .Q(n20068), .QN(n7416)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6088), .CK(CLK), .Q(n20069), .QN(n7418)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6087), .CK(CLK), .Q(n20070), .QN(n7420)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6086), .CK(CLK), .Q(n20071), .QN(n7422)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6085), .CK(CLK), .Q(n20072), .QN(n7424)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6084), .CK(CLK), .Q(n20073), .QN(n7426)
         );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6427), .CK(CLK), .Q(n24171), .QN(n7508)
         );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6426), .CK(CLK), .Q(n24170), .QN(n7510)
         );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6425), .CK(CLK), .Q(n24169), .QN(n7512)
         );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6424), .CK(CLK), .Q(n24168), .QN(n7514)
         );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6423), .CK(CLK), .Q(n24167), .QN(n7516)
         );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6422), .CK(CLK), .Q(n24166), .QN(n7518)
         );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6421), .CK(CLK), .Q(n24165), .QN(n7520)
         );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6420), .CK(CLK), .Q(n24164), .QN(n7522)
         );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6419), .CK(CLK), .Q(n24163), .QN(n7524)
         );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6418), .CK(CLK), .Q(n24162), .QN(n7526)
         );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6417), .CK(CLK), .Q(n24161), .QN(n7528)
         );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6416), .CK(CLK), .Q(n24160), .QN(n7530)
         );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6415), .CK(CLK), .Q(n24159), .QN(n7532)
         );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6414), .CK(CLK), .Q(n24158), .QN(n7534)
         );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6413), .CK(CLK), .Q(n24157), .QN(n7536)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6412), .CK(CLK), .Q(n24156), .QN(n7538)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6411), .CK(CLK), .Q(n24155), .QN(n7540)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6410), .CK(CLK), .Q(n24154), .QN(n7542)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6409), .CK(CLK), .Q(n24153), .QN(n7544)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6408), .CK(CLK), .Q(n24152), .QN(n7546)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6407), .CK(CLK), .Q(n24151), .QN(n7548)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6406), .CK(CLK), .Q(n24150), .QN(n7550)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6405), .CK(CLK), .Q(n24149), .QN(n7552)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6404), .CK(CLK), .Q(n24148), .QN(n7554)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n6747), .CK(CLK), .Q(n24235), .QN(n17341)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n6746), .CK(CLK), .Q(n24234), .QN(n17344)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n6745), .CK(CLK), .Q(n24233), .QN(n17347)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n6744), .CK(CLK), .Q(n24232), .QN(n17350)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n6743), .CK(CLK), .Q(n24231), .QN(n17353)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n6742), .CK(CLK), .Q(n24230), .QN(n17356)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n6741), .CK(CLK), .Q(n24229), .QN(n17359)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n6740), .CK(CLK), .Q(n24228), .QN(n17362)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n6739), .CK(CLK), .Q(n24227), .QN(n17365)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n6738), .CK(CLK), .Q(n24226), .QN(n17368)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n6737), .CK(CLK), .Q(n24225), .QN(n17371)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n6736), .CK(CLK), .Q(n24224), .QN(n17374)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n6735), .CK(CLK), .Q(n24223), .QN(n17377)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n6734), .CK(CLK), .Q(n24222), .QN(n17380)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n6733), .CK(CLK), .Q(n24221), .QN(n17383)
         );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n6732), .CK(CLK), .Q(n24220), .QN(n17386)
         );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n6731), .CK(CLK), .Q(n24219), .QN(n17389)
         );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n6730), .CK(CLK), .Q(n24218), .QN(n17392)
         );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n6729), .CK(CLK), .Q(n24217), .QN(n17395)
         );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n6728), .CK(CLK), .Q(n24216), .QN(n17398)
         );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n6727), .CK(CLK), .Q(n24215), .QN(n17401)
         );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n6726), .CK(CLK), .Q(n24214), .QN(n17404)
         );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n6725), .CK(CLK), .Q(n24213), .QN(n17407)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n6724), .CK(CLK), .Q(n24212), .QN(n17410)
         );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7031), .CK(CLK), .Q(n20122), .QN(n77) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7030), .CK(CLK), .Q(n20123), .QN(n78) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7029), .CK(CLK), .Q(n20124), .QN(n79) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7028), .CK(CLK), .Q(n20125), .QN(n80) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7027), .CK(CLK), .Q(n20126), .QN(n81) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7026), .CK(CLK), .Q(n20127), .QN(n82) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7025), .CK(CLK), .Q(n20128), .QN(n83) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7024), .CK(CLK), .Q(n20129), .QN(n84) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7023), .CK(CLK), .Q(n20130), .QN(n85) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7021), .CK(CLK), .Q(n20131), .QN(n87) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7019), .CK(CLK), .Q(n20132), .QN(n89) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7015), .CK(CLK), .Q(n20133), .QN(n93) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7022), .CK(CLK), .Q(n20134), .QN(n86) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7020), .CK(CLK), .Q(n20135), .QN(n88) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7018), .CK(CLK), .Q(n20136), .QN(n90) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7017), .CK(CLK), .Q(n20137), .QN(n91) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7016), .CK(CLK), .Q(n20138), .QN(n92) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7014), .CK(CLK), .Q(n20139), .QN(n94) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7013), .CK(CLK), .Q(n20140), .QN(n95) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7012), .CK(CLK), .Q(n20141), .QN(n96) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7011), .CK(CLK), .Q(n20142), .QN(n97) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7010), .CK(CLK), .Q(n20143), .QN(n98) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7009), .CK(CLK), .Q(n20144), .QN(n99) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n5635), .CK(CLK), .Q(n20153), .QN(n9119)
         );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n5634), .CK(CLK), .Q(n20154), .QN(n9121)
         );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n5633), .CK(CLK), .Q(n20155), .QN(n9123)
         );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n5632), .CK(CLK), .Q(n20156), .QN(n9125)
         );
  NAND3_X1 U18613 ( .A1(n19192), .A2(n19191), .A3(n21269), .ZN(n21253) );
  NAND3_X1 U18614 ( .A1(n21269), .A2(n19191), .A3(ADD_WR[3]), .ZN(n21271) );
  NAND3_X1 U18615 ( .A1(n21269), .A2(n19192), .A3(ADD_WR[4]), .ZN(n21280) );
  NAND3_X1 U18616 ( .A1(n19194), .A2(n19193), .A3(n19195), .ZN(n21254) );
  NAND3_X1 U18617 ( .A1(n19194), .A2(n19193), .A3(ADD_WR[0]), .ZN(n21256) );
  NAND3_X1 U18618 ( .A1(n19195), .A2(n19193), .A3(ADD_WR[1]), .ZN(n21258) );
  NAND3_X1 U18619 ( .A1(ADD_WR[0]), .A2(n19193), .A3(ADD_WR[1]), .ZN(n21260)
         );
  NAND3_X1 U18620 ( .A1(n19195), .A2(n19194), .A3(ADD_WR[2]), .ZN(n21262) );
  NAND3_X1 U18621 ( .A1(ADD_WR[0]), .A2(n19194), .A3(ADD_WR[2]), .ZN(n21264)
         );
  NAND3_X1 U18622 ( .A1(ADD_WR[1]), .A2(n19195), .A3(ADD_WR[2]), .ZN(n21266)
         );
  NAND3_X1 U18623 ( .A1(ADD_WR[3]), .A2(n21269), .A3(ADD_WR[4]), .ZN(n21289)
         );
  NAND3_X1 U18624 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n21268) );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n5699), .CK(CLK), .Q(n19524), .QN(n7429)
         );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n5698), .CK(CLK), .Q(n19525), .QN(n7431)
         );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n5697), .CK(CLK), .Q(n19526), .QN(n7433)
         );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n5696), .CK(CLK), .Q(n19527), .QN(n7435)
         );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n5955), .CK(CLK), .Q(n19806), .QN(n8735)
         );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n5954), .CK(CLK), .Q(n19807), .QN(n8737)
         );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n5953), .CK(CLK), .Q(n19808), .QN(n8739)
         );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n5952), .CK(CLK), .Q(n19809), .QN(n8741)
         );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6211), .CK(CLK), .Q(n19460), .QN(n8990)
         );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6210), .CK(CLK), .Q(n19461), .QN(n8992)
         );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6209), .CK(CLK), .Q(n19462), .QN(n8994)
         );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6208), .CK(CLK), .Q(n19463), .QN(n8996)
         );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n5695), .CK(CLK), .Q(n19528), .QN(n7437)
         );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n5694), .CK(CLK), .Q(n19529), .QN(n7439)
         );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n5693), .CK(CLK), .Q(n19530), .QN(n7441)
         );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n5692), .CK(CLK), .Q(n19531), .QN(n7443)
         );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n5691), .CK(CLK), .Q(n19532), .QN(n7445)
         );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n5690), .CK(CLK), .Q(n19533), .QN(n7447)
         );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n5689), .CK(CLK), .Q(n19534), .QN(n7449)
         );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n5688), .CK(CLK), .Q(n19535), .QN(n7451)
         );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n5687), .CK(CLK), .Q(n19536), .QN(n7453)
         );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n5686), .CK(CLK), .Q(n19537), .QN(n7455)
         );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n5685), .CK(CLK), .Q(n19538), .QN(n7457)
         );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n5684), .CK(CLK), .Q(n19539), .QN(n7459)
         );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n5683), .CK(CLK), .Q(n19540), .QN(n7461)
         );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n5682), .CK(CLK), .Q(n19541), .QN(n7463)
         );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n5681), .CK(CLK), .Q(n19542), .QN(n7465)
         );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n5680), .CK(CLK), .Q(n19543), .QN(n7467)
         );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n5679), .CK(CLK), .Q(n19544), .QN(n7469)
         );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n5678), .CK(CLK), .Q(n19545), .QN(n7471)
         );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n5677), .CK(CLK), .Q(n19546), .QN(n7473)
         );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n5676), .CK(CLK), .Q(n19547), .QN(n7475)
         );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n5675), .CK(CLK), .Q(n19548), .QN(n7477)
         );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n5674), .CK(CLK), .Q(n19549), .QN(n7479)
         );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n5673), .CK(CLK), .Q(n19550), .QN(n7481)
         );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n5672), .CK(CLK), .Q(n19551), .QN(n7483)
         );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n5671), .CK(CLK), .Q(n19552), .QN(n7485)
         );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n5670), .CK(CLK), .Q(n19553), .QN(n7487)
         );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n5669), .CK(CLK), .Q(n19554), .QN(n7489)
         );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n5668), .CK(CLK), .Q(n19555), .QN(n7491)
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n5667), .CK(CLK), .Q(n19556), .QN(n7493)
         );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n5666), .CK(CLK), .Q(n19557), .QN(n7495)
         );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n5665), .CK(CLK), .Q(n19558), .QN(n7497)
         );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n5664), .CK(CLK), .Q(n19559), .QN(n7499)
         );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n5663), .CK(CLK), .Q(n19560), .QN(n7501)
         );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n5662), .CK(CLK), .Q(n19561), .QN(n7503)
         );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n5661), .CK(CLK), .Q(n19562), .QN(n7505)
         );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n5660), .CK(CLK), .Q(n19563), .QN(n7507)
         );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n5951), .CK(CLK), .Q(n19858), .QN(n8743)
         );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n5950), .CK(CLK), .Q(n19859), .QN(n8745)
         );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n5949), .CK(CLK), .Q(n19860), .QN(n8747)
         );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n5948), .CK(CLK), .Q(n19861), .QN(n8749)
         );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n5947), .CK(CLK), .Q(n19862), .QN(n8751)
         );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n5946), .CK(CLK), .Q(n19863), .QN(n8753)
         );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n5945), .CK(CLK), .Q(n19864), .QN(n8755)
         );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n5944), .CK(CLK), .Q(n19865), .QN(n8757)
         );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n5943), .CK(CLK), .Q(n19866), .QN(n8759)
         );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n5942), .CK(CLK), .Q(n19867), .QN(n8761)
         );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n5941), .CK(CLK), .Q(n19868), .QN(n8763)
         );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n5940), .CK(CLK), .Q(n19869), .QN(n8765)
         );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n5939), .CK(CLK), .Q(n19870), .QN(n8767)
         );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n5938), .CK(CLK), .Q(n19871), .QN(n8769)
         );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n5937), .CK(CLK), .Q(n19872), .QN(n8771)
         );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n5936), .CK(CLK), .Q(n19873), .QN(n8773)
         );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n5935), .CK(CLK), .Q(n19874), .QN(n8775)
         );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n5934), .CK(CLK), .Q(n19875), .QN(n8777)
         );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n5933), .CK(CLK), .Q(n19876), .QN(n8779)
         );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n5932), .CK(CLK), .Q(n19877), .QN(n8781)
         );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n5931), .CK(CLK), .Q(n19878), .QN(n8783)
         );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n5930), .CK(CLK), .Q(n19879), .QN(n8785)
         );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n5929), .CK(CLK), .Q(n19880), .QN(n8787)
         );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n5928), .CK(CLK), .Q(n19881), .QN(n8789)
         );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n5927), .CK(CLK), .Q(n19882), .QN(n8791)
         );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n5926), .CK(CLK), .Q(n19883), .QN(n8793)
         );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n5925), .CK(CLK), .Q(n19884), .QN(n8795)
         );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n5924), .CK(CLK), .Q(n19885), .QN(n8797)
         );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n5923), .CK(CLK), .Q(n19886), .QN(n8799)
         );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n5922), .CK(CLK), .Q(n19887), .QN(n8801)
         );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n5921), .CK(CLK), .Q(n19888), .QN(n8803)
         );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n5920), .CK(CLK), .Q(n19889), .QN(n8805)
         );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n5919), .CK(CLK), .Q(n19890), .QN(n8807)
         );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n5918), .CK(CLK), .Q(n19891), .QN(n8809)
         );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n5917), .CK(CLK), .Q(n19892), .QN(n8811)
         );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n5916), .CK(CLK), .Q(n19893), .QN(n8813)
         );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6207), .CK(CLK), .Q(n19464), .QN(n8998)
         );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6206), .CK(CLK), .Q(n19465), .QN(n9000)
         );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6205), .CK(CLK), .Q(n19466), .QN(n9002)
         );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6204), .CK(CLK), .Q(n19467), .QN(n9004)
         );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6203), .CK(CLK), .Q(n19468), .QN(n9006)
         );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6202), .CK(CLK), .Q(n19469), .QN(n9008)
         );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6201), .CK(CLK), .Q(n19470), .QN(n9010)
         );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6200), .CK(CLK), .Q(n19471), .QN(n9012)
         );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6199), .CK(CLK), .Q(n19472), .QN(n9014)
         );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6198), .CK(CLK), .Q(n19473), .QN(n9016)
         );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6197), .CK(CLK), .Q(n19474), .QN(n9018)
         );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6196), .CK(CLK), .Q(n19475), .QN(n9020)
         );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6195), .CK(CLK), .Q(n19476), .QN(n9022)
         );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6194), .CK(CLK), .Q(n19477), .QN(n9024)
         );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6193), .CK(CLK), .Q(n19478), .QN(n9026)
         );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6192), .CK(CLK), .Q(n19479), .QN(n9028)
         );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6191), .CK(CLK), .Q(n19480), .QN(n9030)
         );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6190), .CK(CLK), .Q(n19481), .QN(n9032)
         );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6189), .CK(CLK), .Q(n19482), .QN(n9034)
         );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6188), .CK(CLK), .Q(n19483), .QN(n9036)
         );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6187), .CK(CLK), .Q(n19484), .QN(n9038)
         );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6186), .CK(CLK), .Q(n19485), .QN(n9040)
         );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6185), .CK(CLK), .Q(n19486), .QN(n9042)
         );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6184), .CK(CLK), .Q(n19487), .QN(n9044)
         );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6183), .CK(CLK), .Q(n19488), .QN(n9046)
         );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6182), .CK(CLK), .Q(n19489), .QN(n9048)
         );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6181), .CK(CLK), .Q(n19490), .QN(n9050)
         );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6180), .CK(CLK), .Q(n19491), .QN(n9052)
         );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6179), .CK(CLK), .Q(n19492), .QN(n9054)
         );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6178), .CK(CLK), .Q(n19493), .QN(n9056)
         );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6177), .CK(CLK), .Q(n19494), .QN(n9058)
         );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6176), .CK(CLK), .Q(n19495), .QN(n9060)
         );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6175), .CK(CLK), .Q(n19496), .QN(n9062)
         );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6174), .CK(CLK), .Q(n19497), .QN(n9064)
         );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6173), .CK(CLK), .Q(n19498), .QN(n9066)
         );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6172), .CK(CLK), .Q(n19499), .QN(n9068)
         );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n5659), .CK(CLK), .Q(n19564), .QN(n7509)
         );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n5658), .CK(CLK), .Q(n19565), .QN(n7511)
         );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n5657), .CK(CLK), .Q(n19566), .QN(n7513)
         );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n5656), .CK(CLK), .Q(n19567), .QN(n7515)
         );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n5655), .CK(CLK), .Q(n19568), .QN(n7517)
         );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n5654), .CK(CLK), .Q(n19569), .QN(n7519)
         );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n5653), .CK(CLK), .Q(n19570), .QN(n7521)
         );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n5652), .CK(CLK), .Q(n19571), .QN(n7523)
         );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n5651), .CK(CLK), .Q(n19572), .QN(n7525)
         );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n5650), .CK(CLK), .Q(n19573), .QN(n7527)
         );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n5649), .CK(CLK), .Q(n19574), .QN(n7529)
         );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n5648), .CK(CLK), .Q(n19575), .QN(n7531)
         );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n5647), .CK(CLK), .Q(n19576), .QN(n7533)
         );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n5646), .CK(CLK), .Q(n19577), .QN(n7535)
         );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n5645), .CK(CLK), .Q(n19578), .QN(n7537)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n5644), .CK(CLK), .Q(n19579), .QN(n7539)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n5643), .CK(CLK), .Q(n19580), .QN(n7541)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n5642), .CK(CLK), .Q(n19581), .QN(n7543)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n5641), .CK(CLK), .Q(n19582), .QN(n7545)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n5640), .CK(CLK), .Q(n19583), .QN(n7547)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n5639), .CK(CLK), .Q(n19584), .QN(n7549)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n5638), .CK(CLK), .Q(n19585), .QN(n7551)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n5637), .CK(CLK), .Q(n19586), .QN(n7553)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n5636), .CK(CLK), .Q(n19587), .QN(n7555)
         );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n5915), .CK(CLK), .Q(n20026), .QN(n8815)
         );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n5914), .CK(CLK), .Q(n20027), .QN(n8817)
         );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n5913), .CK(CLK), .Q(n20028), .QN(n8819)
         );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n5912), .CK(CLK), .Q(n20029), .QN(n8821)
         );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n5911), .CK(CLK), .Q(n20030), .QN(n8823)
         );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n5910), .CK(CLK), .Q(n20031), .QN(n8825)
         );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n5909), .CK(CLK), .Q(n20032), .QN(n8827)
         );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n5908), .CK(CLK), .Q(n20033), .QN(n8829)
         );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n5907), .CK(CLK), .Q(n20034), .QN(n8831)
         );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n5906), .CK(CLK), .Q(n20035), .QN(n8833)
         );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n5905), .CK(CLK), .Q(n20036), .QN(n8835)
         );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n5904), .CK(CLK), .Q(n20037), .QN(n8837)
         );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n5903), .CK(CLK), .Q(n20038), .QN(n8839)
         );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n5902), .CK(CLK), .Q(n20039), .QN(n8841)
         );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n5901), .CK(CLK), .Q(n20040), .QN(n8843)
         );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n5900), .CK(CLK), .Q(n20041), .QN(n8845)
         );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n5899), .CK(CLK), .Q(n20042), .QN(n8847)
         );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n5898), .CK(CLK), .Q(n20043), .QN(n8849)
         );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n5897), .CK(CLK), .Q(n20044), .QN(n8851)
         );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n5896), .CK(CLK), .Q(n20045), .QN(n8853)
         );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n5895), .CK(CLK), .Q(n20046), .QN(n8855)
         );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n5894), .CK(CLK), .Q(n20047), .QN(n8857)
         );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n5893), .CK(CLK), .Q(n20048), .QN(n8859)
         );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n5892), .CK(CLK), .Q(n20049), .QN(n8861)
         );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6171), .CK(CLK), .Q(n19500), .QN(n9070)
         );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6170), .CK(CLK), .Q(n19501), .QN(n9072)
         );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6169), .CK(CLK), .Q(n19502), .QN(n9074)
         );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6168), .CK(CLK), .Q(n19503), .QN(n9076)
         );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6167), .CK(CLK), .Q(n19504), .QN(n9078)
         );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6166), .CK(CLK), .Q(n19505), .QN(n9080)
         );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6165), .CK(CLK), .Q(n19506), .QN(n9082)
         );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6164), .CK(CLK), .Q(n19507), .QN(n9084)
         );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6163), .CK(CLK), .Q(n19508), .QN(n9086)
         );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6162), .CK(CLK), .Q(n19509), .QN(n9088)
         );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6161), .CK(CLK), .Q(n19510), .QN(n9090)
         );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6160), .CK(CLK), .Q(n19511), .QN(n9092)
         );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6159), .CK(CLK), .Q(n19512), .QN(n9094)
         );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6158), .CK(CLK), .Q(n19513), .QN(n9096)
         );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6157), .CK(CLK), .Q(n19514), .QN(n9098)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6156), .CK(CLK), .Q(n19515), .QN(n9100)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6155), .CK(CLK), .Q(n19516), .QN(n9102)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6154), .CK(CLK), .Q(n19517), .QN(n9104)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6153), .CK(CLK), .Q(n19518), .QN(n9106)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6152), .CK(CLK), .Q(n19519), .QN(n9108)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6151), .CK(CLK), .Q(n19520), .QN(n9110)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6150), .CK(CLK), .Q(n19521), .QN(n9112)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6149), .CK(CLK), .Q(n19522), .QN(n9114)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6148), .CK(CLK), .Q(n19523), .QN(n9116)
         );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5507), .CK(CLK), .QN(n7301) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5063), .CK(CLK), .Q(n8282), .QN(n20187)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5062), .CK(CLK), .Q(n8283), .QN(n20188)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5061), .CK(CLK), .Q(n8284), .QN(n20189)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5060), .CK(CLK), .Q(n8285), .QN(n20526)
         );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5099), .CK(CLK), .Q(n8246), .QN(n20214)
         );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5098), .CK(CLK), .Q(n8247), .QN(n20215)
         );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5097), .CK(CLK), .Q(n8248), .QN(n20216)
         );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5096), .CK(CLK), .Q(n8249), .QN(n20217)
         );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5095), .CK(CLK), .Q(n8250), .QN(n20218)
         );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5094), .CK(CLK), .Q(n8251), .QN(n20219)
         );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5093), .CK(CLK), .Q(n8252), .QN(n20220)
         );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5092), .CK(CLK), .Q(n8253), .QN(n20221)
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5091), .CK(CLK), .Q(n8254), .QN(n20222)
         );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5090), .CK(CLK), .Q(n8255), .QN(n20223)
         );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5089), .CK(CLK), .Q(n8256), .QN(n20224)
         );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5088), .CK(CLK), .Q(n8257), .QN(n20225)
         );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5087), .CK(CLK), .Q(n8258), .QN(n20226)
         );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5086), .CK(CLK), .Q(n8259), .QN(n20227)
         );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5085), .CK(CLK), .Q(n8260), .QN(n20228)
         );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5084), .CK(CLK), .Q(n8261), .QN(n20229)
         );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5083), .CK(CLK), .Q(n8262), .QN(n20230)
         );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5082), .CK(CLK), .Q(n8263), .QN(n20231)
         );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5081), .CK(CLK), .Q(n8264), .QN(n20232)
         );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5080), .CK(CLK), .Q(n8265), .QN(n20233)
         );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5079), .CK(CLK), .Q(n8266), .QN(n20234)
         );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5078), .CK(CLK), .Q(n8267), .QN(n20235)
         );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5077), .CK(CLK), .Q(n8268), .QN(n20236)
         );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5076), .CK(CLK), .Q(n8269), .QN(n20237)
         );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5075), .CK(CLK), .Q(n8270), .QN(n20238)
         );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5074), .CK(CLK), .Q(n8271), .QN(n20239)
         );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5073), .CK(CLK), .Q(n8272), .QN(n20240)
         );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5072), .CK(CLK), .Q(n8273), .QN(n20241)
         );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5071), .CK(CLK), .Q(n8274), .QN(n20242)
         );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5070), .CK(CLK), .Q(n8275), .QN(n20243)
         );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5069), .CK(CLK), .Q(n8276), .QN(n20244)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5068), .CK(CLK), .Q(n8277), .QN(n20245)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5067), .CK(CLK), .Q(n8278), .QN(n20246)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5066), .CK(CLK), .Q(n8279), .QN(n20247)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5065), .CK(CLK), .Q(n8280), .QN(n20248)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5064), .CK(CLK), .Q(n8281), .QN(n20249)
         );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5123), .CK(CLK), .Q(n8222), .QN(n20190)
         );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5122), .CK(CLK), .Q(n8223), .QN(n20191)
         );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5121), .CK(CLK), .Q(n8224), .QN(n20192)
         );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5120), .CK(CLK), .Q(n8225), .QN(n20193)
         );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5119), .CK(CLK), .Q(n8226), .QN(n20194)
         );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5118), .CK(CLK), .Q(n8227), .QN(n20195)
         );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5117), .CK(CLK), .Q(n8228), .QN(n20196)
         );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5116), .CK(CLK), .Q(n8229), .QN(n20197)
         );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5115), .CK(CLK), .Q(n8230), .QN(n20198)
         );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5114), .CK(CLK), .Q(n8231), .QN(n20199)
         );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5113), .CK(CLK), .Q(n8232), .QN(n20200)
         );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5112), .CK(CLK), .Q(n8233), .QN(n20201)
         );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5111), .CK(CLK), .Q(n8234), .QN(n20202)
         );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5110), .CK(CLK), .Q(n8235), .QN(n20203)
         );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5109), .CK(CLK), .Q(n8236), .QN(n20204)
         );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5108), .CK(CLK), .Q(n8237), .QN(n20205)
         );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5107), .CK(CLK), .Q(n8238), .QN(n20206)
         );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5106), .CK(CLK), .Q(n8239), .QN(n20207)
         );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5105), .CK(CLK), .Q(n8240), .QN(n20208)
         );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5104), .CK(CLK), .Q(n8241), .QN(n20209)
         );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5103), .CK(CLK), .Q(n8242), .QN(n20210)
         );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5102), .CK(CLK), .Q(n8243), .QN(n20211)
         );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5101), .CK(CLK), .Q(n8244), .QN(n20212)
         );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5100), .CK(CLK), .Q(n8245), .QN(n20213)
         );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n5827), .CK(CLK), .QN(n20514) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n5826), .CK(CLK), .QN(n20515) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n5825), .CK(CLK), .QN(n20516) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n5824), .CK(CLK), .QN(n20517) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n6915), .CK(CLK), .QN(n20250) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n6914), .CK(CLK), .QN(n20251) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n6913), .CK(CLK), .QN(n20252) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n6912), .CK(CLK), .QN(n20253) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n6019), .CK(CLK), .QN(n20262) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n6018), .CK(CLK), .QN(n20263) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n6017), .CK(CLK), .QN(n20264) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n6016), .CK(CLK), .QN(n20265) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5571), .CK(CLK), .QN(n20149) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5570), .CK(CLK), .QN(n20150) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5569), .CK(CLK), .QN(n20151) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5568), .CK(CLK), .QN(n20152) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n6659), .CK(CLK), .QN(n20539) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n6658), .CK(CLK), .QN(n20540) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n6657), .CK(CLK), .QN(n20541) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n6656), .CK(CLK), .QN(n20542) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n6723), .CK(CLK), .QN(n20522) );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n6722), .CK(CLK), .QN(n20523) );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n6721), .CK(CLK), .QN(n20524) );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n6720), .CK(CLK), .QN(n20525) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n6979), .CK(CLK), .QN(n20258) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n6978), .CK(CLK), .QN(n20259) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n6977), .CK(CLK), .QN(n20260) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n6976), .CK(CLK), .QN(n20261) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n5823), .CK(CLK), .QN(n20619) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n5822), .CK(CLK), .QN(n20620) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n5821), .CK(CLK), .QN(n20621) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n5820), .CK(CLK), .QN(n20622) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n5819), .CK(CLK), .QN(n20623) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n5818), .CK(CLK), .QN(n20624) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n5817), .CK(CLK), .QN(n20625) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n5816), .CK(CLK), .QN(n20626) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n5815), .CK(CLK), .QN(n20627) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n5814), .CK(CLK), .QN(n20628) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n5813), .CK(CLK), .QN(n20629) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n5812), .CK(CLK), .QN(n20630) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n5811), .CK(CLK), .QN(n20631) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n5810), .CK(CLK), .QN(n20632) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n5809), .CK(CLK), .QN(n20633) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n5808), .CK(CLK), .QN(n20634) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n5807), .CK(CLK), .QN(n20635) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n5806), .CK(CLK), .QN(n20636) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n5805), .CK(CLK), .QN(n20637) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n5804), .CK(CLK), .QN(n20638) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n5803), .CK(CLK), .QN(n20639) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n5802), .CK(CLK), .QN(n20640) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n5801), .CK(CLK), .QN(n20641) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n5800), .CK(CLK), .QN(n20642) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n5799), .CK(CLK), .QN(n20643) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n5798), .CK(CLK), .QN(n20644) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n5797), .CK(CLK), .QN(n20645) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n5796), .CK(CLK), .QN(n20646) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n5795), .CK(CLK), .QN(n20647) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n5794), .CK(CLK), .QN(n20648) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n5793), .CK(CLK), .QN(n20649) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n5792), .CK(CLK), .QN(n20650) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n5791), .CK(CLK), .QN(n20651) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n5790), .CK(CLK), .QN(n20652) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n5789), .CK(CLK), .QN(n20653) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n5788), .CK(CLK), .QN(n20654) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n6911), .CK(CLK), .QN(n20266) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n6910), .CK(CLK), .QN(n20267) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n6909), .CK(CLK), .QN(n20268) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n6908), .CK(CLK), .QN(n20269) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n6907), .CK(CLK), .QN(n20270) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n6906), .CK(CLK), .QN(n20271) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n6905), .CK(CLK), .QN(n20272) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n6904), .CK(CLK), .QN(n20273) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n6903), .CK(CLK), .QN(n20274) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n6902), .CK(CLK), .QN(n20275) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n6901), .CK(CLK), .QN(n20276) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n6900), .CK(CLK), .QN(n20277) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n6899), .CK(CLK), .QN(n20278) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n6898), .CK(CLK), .QN(n20279) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n6897), .CK(CLK), .QN(n20280) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n6896), .CK(CLK), .QN(n20281) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n6895), .CK(CLK), .QN(n20282) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n6894), .CK(CLK), .QN(n20283) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n6893), .CK(CLK), .QN(n20284) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n6892), .CK(CLK), .QN(n20285) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n6891), .CK(CLK), .QN(n20286) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n6890), .CK(CLK), .QN(n20287) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n6889), .CK(CLK), .QN(n20288) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n6888), .CK(CLK), .QN(n20289) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n6887), .CK(CLK), .QN(n20290) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n6886), .CK(CLK), .QN(n20291) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n6885), .CK(CLK), .QN(n20292) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n6884), .CK(CLK), .QN(n20293) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n6883), .CK(CLK), .QN(n20294) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n6882), .CK(CLK), .QN(n20295) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n6881), .CK(CLK), .QN(n20296) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n6880), .CK(CLK), .QN(n20297) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n6879), .CK(CLK), .QN(n20298) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n6878), .CK(CLK), .QN(n20299) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n6877), .CK(CLK), .QN(n20300) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n6876), .CK(CLK), .QN(n20301) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n5787), .CK(CLK), .QN(n20775) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n5786), .CK(CLK), .QN(n20776) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n5785), .CK(CLK), .QN(n20777) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n5784), .CK(CLK), .QN(n20778) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n5783), .CK(CLK), .QN(n20779) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n5782), .CK(CLK), .QN(n20780) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n5781), .CK(CLK), .QN(n20781) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n5780), .CK(CLK), .QN(n20782) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n5779), .CK(CLK), .QN(n20783) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n5778), .CK(CLK), .QN(n20784) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n5777), .CK(CLK), .QN(n20785) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n5776), .CK(CLK), .QN(n20786) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n5775), .CK(CLK), .QN(n20787) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n5774), .CK(CLK), .QN(n20788) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n5773), .CK(CLK), .QN(n20789) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n5772), .CK(CLK), .QN(n20790) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n5771), .CK(CLK), .QN(n20791) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n5770), .CK(CLK), .QN(n20792) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n5769), .CK(CLK), .QN(n20793) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n5768), .CK(CLK), .QN(n20794) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n5767), .CK(CLK), .QN(n20795) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n5766), .CK(CLK), .QN(n20796) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n5765), .CK(CLK), .QN(n20797) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n5764), .CK(CLK), .QN(n20798) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n6875), .CK(CLK), .QN(n20374) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n6874), .CK(CLK), .QN(n20375) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n6873), .CK(CLK), .QN(n20376) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n6872), .CK(CLK), .QN(n20377) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n6871), .CK(CLK), .QN(n20378) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n6870), .CK(CLK), .QN(n20379) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n6869), .CK(CLK), .QN(n20380) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n6868), .CK(CLK), .QN(n20381) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n6867), .CK(CLK), .QN(n20382) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n6866), .CK(CLK), .QN(n20383) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n6865), .CK(CLK), .QN(n20384) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n6864), .CK(CLK), .QN(n20385) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n6863), .CK(CLK), .QN(n20386) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n6862), .CK(CLK), .QN(n20387) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n6861), .CK(CLK), .QN(n20388) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n6860), .CK(CLK), .QN(n20389) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n6859), .CK(CLK), .QN(n20390) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n6858), .CK(CLK), .QN(n20391) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n6857), .CK(CLK), .QN(n20392) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n6856), .CK(CLK), .QN(n20393) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n6855), .CK(CLK), .QN(n20394) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n6854), .CK(CLK), .QN(n20395) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n6853), .CK(CLK), .QN(n20396) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n6852), .CK(CLK), .QN(n20397) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n6015), .CK(CLK), .QN(n20446) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n6014), .CK(CLK), .QN(n20447) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n6013), .CK(CLK), .QN(n20448) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n6012), .CK(CLK), .QN(n20449) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n6011), .CK(CLK), .QN(n20450) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n6010), .CK(CLK), .QN(n20451) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n6009), .CK(CLK), .QN(n20452) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n6008), .CK(CLK), .QN(n20453) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n6007), .CK(CLK), .QN(n20454) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n6006), .CK(CLK), .QN(n20455) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n6005), .CK(CLK), .QN(n20456) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n6004), .CK(CLK), .QN(n20457) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n6003), .CK(CLK), .QN(n20458) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n6002), .CK(CLK), .QN(n20459) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n6001), .CK(CLK), .QN(n20460) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n6000), .CK(CLK), .QN(n20461) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n5999), .CK(CLK), .QN(n20462) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n5998), .CK(CLK), .QN(n20463) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n5997), .CK(CLK), .QN(n20464) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n5996), .CK(CLK), .QN(n20465) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n5995), .CK(CLK), .QN(n20466) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n5994), .CK(CLK), .QN(n20467) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n5993), .CK(CLK), .QN(n20468) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n5992), .CK(CLK), .QN(n20469) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n5991), .CK(CLK), .QN(n20470) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n5990), .CK(CLK), .QN(n20471) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n5989), .CK(CLK), .QN(n20472) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n5988), .CK(CLK), .QN(n20473) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n5987), .CK(CLK), .QN(n20474) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n5986), .CK(CLK), .QN(n20475) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n5985), .CK(CLK), .QN(n20476) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n5984), .CK(CLK), .QN(n20477) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n5983), .CK(CLK), .QN(n20478) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n5982), .CK(CLK), .QN(n20479) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n5981), .CK(CLK), .QN(n20480) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n5980), .CK(CLK), .QN(n20481) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5567), .CK(CLK), .QN(n19648) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5566), .CK(CLK), .QN(n19649) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5565), .CK(CLK), .QN(n19650) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5564), .CK(CLK), .QN(n19651) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5563), .CK(CLK), .QN(n19652) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5562), .CK(CLK), .QN(n19653) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5561), .CK(CLK), .QN(n19654) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5560), .CK(CLK), .QN(n19655) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5559), .CK(CLK), .QN(n19656) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5558), .CK(CLK), .QN(n19657) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5557), .CK(CLK), .QN(n19658) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5556), .CK(CLK), .QN(n19659) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5555), .CK(CLK), .QN(n19660) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5554), .CK(CLK), .QN(n19661) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5553), .CK(CLK), .QN(n19662) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5552), .CK(CLK), .QN(n19663) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5551), .CK(CLK), .QN(n19664) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5550), .CK(CLK), .QN(n19665) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5549), .CK(CLK), .QN(n19666) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5548), .CK(CLK), .QN(n19667) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5547), .CK(CLK), .QN(n19668) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5546), .CK(CLK), .QN(n19669) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5545), .CK(CLK), .QN(n19670) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5544), .CK(CLK), .QN(n19671) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5543), .CK(CLK), .QN(n19672) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5542), .CK(CLK), .QN(n19673) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5541), .CK(CLK), .QN(n19674) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5540), .CK(CLK), .QN(n19675) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5539), .CK(CLK), .QN(n19676) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5538), .CK(CLK), .QN(n19677) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5537), .CK(CLK), .QN(n19678) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5536), .CK(CLK), .QN(n19679) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5535), .CK(CLK), .QN(n19680) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5534), .CK(CLK), .QN(n19681) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5533), .CK(CLK), .QN(n19682) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5532), .CK(CLK), .QN(n19683) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n6655), .CK(CLK), .QN(n20979) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n6654), .CK(CLK), .QN(n20980) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n6653), .CK(CLK), .QN(n20981) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n6652), .CK(CLK), .QN(n20982) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n6651), .CK(CLK), .QN(n20983) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n6650), .CK(CLK), .QN(n20984) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n6649), .CK(CLK), .QN(n20985) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n6648), .CK(CLK), .QN(n20986) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n6647), .CK(CLK), .QN(n20987) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n6646), .CK(CLK), .QN(n20988) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n6645), .CK(CLK), .QN(n20989) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n6644), .CK(CLK), .QN(n20990) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n6643), .CK(CLK), .QN(n20991) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n6642), .CK(CLK), .QN(n20992) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n6641), .CK(CLK), .QN(n20993) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n6640), .CK(CLK), .QN(n20994) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n6639), .CK(CLK), .QN(n20995) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n6638), .CK(CLK), .QN(n20996) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n6637), .CK(CLK), .QN(n20997) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n6636), .CK(CLK), .QN(n20998) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n6635), .CK(CLK), .QN(n20999) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n6634), .CK(CLK), .QN(n21000) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n6633), .CK(CLK), .QN(n21001) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n6632), .CK(CLK), .QN(n21002) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n6631), .CK(CLK), .QN(n21003) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n6630), .CK(CLK), .QN(n21004) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n6629), .CK(CLK), .QN(n21005) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n6628), .CK(CLK), .QN(n21006) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n6627), .CK(CLK), .QN(n21007) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n6626), .CK(CLK), .QN(n21008) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n6625), .CK(CLK), .QN(n21009) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n6624), .CK(CLK), .QN(n21010) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n6623), .CK(CLK), .QN(n21011) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n6622), .CK(CLK), .QN(n21012) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n6621), .CK(CLK), .QN(n21013) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6620), .CK(CLK), .QN(n21014) );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n6719), .CK(CLK), .QN(n20691) );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n6718), .CK(CLK), .QN(n20692) );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n6717), .CK(CLK), .QN(n20693) );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n6716), .CK(CLK), .QN(n20694) );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n6715), .CK(CLK), .QN(n20695) );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n6714), .CK(CLK), .QN(n20696) );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n6713), .CK(CLK), .QN(n20697) );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n6712), .CK(CLK), .QN(n20698) );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n6711), .CK(CLK), .QN(n20699) );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n6710), .CK(CLK), .QN(n20700) );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n6709), .CK(CLK), .QN(n20701) );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n6708), .CK(CLK), .QN(n20702) );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n6707), .CK(CLK), .QN(n20703) );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n6706), .CK(CLK), .QN(n20704) );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n6705), .CK(CLK), .QN(n20705) );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n6704), .CK(CLK), .QN(n20706) );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n6703), .CK(CLK), .QN(n20707) );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n6702), .CK(CLK), .QN(n20708) );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n6701), .CK(CLK), .QN(n20709) );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n6700), .CK(CLK), .QN(n20710) );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n6699), .CK(CLK), .QN(n20711) );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n6698), .CK(CLK), .QN(n20712) );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n6697), .CK(CLK), .QN(n20713) );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n6696), .CK(CLK), .QN(n20714) );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n6695), .CK(CLK), .QN(n20715) );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n6694), .CK(CLK), .QN(n20716) );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n6693), .CK(CLK), .QN(n20717) );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n6692), .CK(CLK), .QN(n20718) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n6691), .CK(CLK), .QN(n20719) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n6690), .CK(CLK), .QN(n20720) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n6689), .CK(CLK), .QN(n20721) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n6688), .CK(CLK), .QN(n20722) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n6687), .CK(CLK), .QN(n20723) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n6686), .CK(CLK), .QN(n20724) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n6685), .CK(CLK), .QN(n20725) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n6684), .CK(CLK), .QN(n20726) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n6975), .CK(CLK), .QN(n20338) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n6974), .CK(CLK), .QN(n20339) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n6973), .CK(CLK), .QN(n20340) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n6972), .CK(CLK), .QN(n20341) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n6971), .CK(CLK), .QN(n20342) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n6970), .CK(CLK), .QN(n20343) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n6969), .CK(CLK), .QN(n20344) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n6968), .CK(CLK), .QN(n20345) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n6967), .CK(CLK), .QN(n20346) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n6966), .CK(CLK), .QN(n20347) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n6965), .CK(CLK), .QN(n20348) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n6964), .CK(CLK), .QN(n20349) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n6963), .CK(CLK), .QN(n20350) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n6962), .CK(CLK), .QN(n20351) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n6961), .CK(CLK), .QN(n20352) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n6960), .CK(CLK), .QN(n20353) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n6959), .CK(CLK), .QN(n20354) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n6958), .CK(CLK), .QN(n20355) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n6957), .CK(CLK), .QN(n20356) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n6956), .CK(CLK), .QN(n20357) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n6955), .CK(CLK), .QN(n20358) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n6954), .CK(CLK), .QN(n20359) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n6953), .CK(CLK), .QN(n20360) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n6952), .CK(CLK), .QN(n20361) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n6951), .CK(CLK), .QN(n20362) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n6950), .CK(CLK), .QN(n20363) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n6949), .CK(CLK), .QN(n20364) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n6948), .CK(CLK), .QN(n20365) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n6947), .CK(CLK), .QN(n20366) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n6946), .CK(CLK), .QN(n20367) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n6945), .CK(CLK), .QN(n20368) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n6944), .CK(CLK), .QN(n20369) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n6943), .CK(CLK), .QN(n20370) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n6942), .CK(CLK), .QN(n20371) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n6941), .CK(CLK), .QN(n20372) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n6940), .CK(CLK), .QN(n20373) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n5979), .CK(CLK), .QN(n20482) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n5978), .CK(CLK), .QN(n20483) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n5977), .CK(CLK), .QN(n20484) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n5976), .CK(CLK), .QN(n20485) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n5975), .CK(CLK), .QN(n20486) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n5974), .CK(CLK), .QN(n20487) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n5973), .CK(CLK), .QN(n20488) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n5972), .CK(CLK), .QN(n20489) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n5971), .CK(CLK), .QN(n20490) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n5970), .CK(CLK), .QN(n20491) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n5969), .CK(CLK), .QN(n20492) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n5968), .CK(CLK), .QN(n20493) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n5967), .CK(CLK), .QN(n20494) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n5966), .CK(CLK), .QN(n20495) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n5965), .CK(CLK), .QN(n20496) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n5964), .CK(CLK), .QN(n20497) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n5963), .CK(CLK), .QN(n20498) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n5962), .CK(CLK), .QN(n20499) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n5961), .CK(CLK), .QN(n20500) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n5960), .CK(CLK), .QN(n20501) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n5959), .CK(CLK), .QN(n20502) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n5958), .CK(CLK), .QN(n20503) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n5957), .CK(CLK), .QN(n20504) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n5956), .CK(CLK), .QN(n20505) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5531), .CK(CLK), .QN(n19684) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5530), .CK(CLK), .QN(n19685) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5529), .CK(CLK), .QN(n19686) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5528), .CK(CLK), .QN(n19687) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5527), .CK(CLK), .QN(n19688) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5526), .CK(CLK), .QN(n19689) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5525), .CK(CLK), .QN(n19690) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5524), .CK(CLK), .QN(n19691) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5523), .CK(CLK), .QN(n19692) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5522), .CK(CLK), .QN(n19693) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5521), .CK(CLK), .QN(n19694) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5520), .CK(CLK), .QN(n19695) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5519), .CK(CLK), .QN(n19696) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5518), .CK(CLK), .QN(n19697) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5517), .CK(CLK), .QN(n19698) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5516), .CK(CLK), .QN(n19699) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5515), .CK(CLK), .QN(n19700) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5514), .CK(CLK), .QN(n19701) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5513), .CK(CLK), .QN(n19702) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5512), .CK(CLK), .QN(n19703) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5511), .CK(CLK), .QN(n19704) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5510), .CK(CLK), .QN(n19705) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5509), .CK(CLK), .QN(n19706) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5508), .CK(CLK), .QN(n19707) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6619), .CK(CLK), .QN(n21099) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6618), .CK(CLK), .QN(n21100) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6617), .CK(CLK), .QN(n21101) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6616), .CK(CLK), .QN(n21102) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6615), .CK(CLK), .QN(n21103) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6614), .CK(CLK), .QN(n21104) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6613), .CK(CLK), .QN(n21105) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6612), .CK(CLK), .QN(n21106) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6611), .CK(CLK), .QN(n21107) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6610), .CK(CLK), .QN(n21108) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6609), .CK(CLK), .QN(n21109) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6608), .CK(CLK), .QN(n21110) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6607), .CK(CLK), .QN(n21111) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6606), .CK(CLK), .QN(n21112) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6605), .CK(CLK), .QN(n21113) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6604), .CK(CLK), .QN(n21114) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6603), .CK(CLK), .QN(n21115) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6602), .CK(CLK), .QN(n21116) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6601), .CK(CLK), .QN(n21117) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6600), .CK(CLK), .QN(n21118) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6599), .CK(CLK), .QN(n21119) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6598), .CK(CLK), .QN(n21120) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6597), .CK(CLK), .QN(n21121) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6596), .CK(CLK), .QN(n21122) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n6683), .CK(CLK), .QN(n20823) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n6682), .CK(CLK), .QN(n20824) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n6681), .CK(CLK), .QN(n20825) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n6680), .CK(CLK), .QN(n20826) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n6679), .CK(CLK), .QN(n20827) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n6678), .CK(CLK), .QN(n20828) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n6677), .CK(CLK), .QN(n20829) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n6676), .CK(CLK), .QN(n20830) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n6675), .CK(CLK), .QN(n20831) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n6674), .CK(CLK), .QN(n20832) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n6673), .CK(CLK), .QN(n20833) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n6672), .CK(CLK), .QN(n20834) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n6671), .CK(CLK), .QN(n20835) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n6670), .CK(CLK), .QN(n20836) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n6669), .CK(CLK), .QN(n20837) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n6668), .CK(CLK), .QN(n20838) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n6667), .CK(CLK), .QN(n20839) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n6666), .CK(CLK), .QN(n20840) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n6665), .CK(CLK), .QN(n20841) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n6664), .CK(CLK), .QN(n20842) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n6663), .CK(CLK), .QN(n20843) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n6662), .CK(CLK), .QN(n20844) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n6661), .CK(CLK), .QN(n20845) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n6660), .CK(CLK), .QN(n20846) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n6939), .CK(CLK), .QN(n20422) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n6938), .CK(CLK), .QN(n20423) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n6937), .CK(CLK), .QN(n20424) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n6936), .CK(CLK), .QN(n20425) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n6935), .CK(CLK), .QN(n20426) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n6934), .CK(CLK), .QN(n20427) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n6933), .CK(CLK), .QN(n20428) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n6932), .CK(CLK), .QN(n20429) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n6931), .CK(CLK), .QN(n20430) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n6930), .CK(CLK), .QN(n20431) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n6929), .CK(CLK), .QN(n20432) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n6928), .CK(CLK), .QN(n20433) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n6927), .CK(CLK), .QN(n20434) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n6926), .CK(CLK), .QN(n20435) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n6925), .CK(CLK), .QN(n20436) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n6924), .CK(CLK), .QN(n20437) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n6923), .CK(CLK), .QN(n20438) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n6922), .CK(CLK), .QN(n20439) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n6921), .CK(CLK), .QN(n20440) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n6920), .CK(CLK), .QN(n20441) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n6919), .CK(CLK), .QN(n20442) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n6918), .CK(CLK), .QN(n20443) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n6917), .CK(CLK), .QN(n20444) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n6916), .CK(CLK), .QN(n20445) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n6851), .CK(CLK), .Q(n17661), .QN(n19332)
         );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n6850), .CK(CLK), .Q(n17658), .QN(n19333)
         );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n6849), .CK(CLK), .Q(n17655), .QN(n19334)
         );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n6848), .CK(CLK), .Q(n17652), .QN(n19335)
         );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n5763), .CK(CLK), .Q(n8478), .QN(n20543)
         );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n5762), .CK(CLK), .Q(n8479), .QN(n20544)
         );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n5761), .CK(CLK), .Q(n8480), .QN(n20545)
         );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n5760), .CK(CLK), .Q(n8481), .QN(n20546)
         );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6083), .CK(CLK), .Q(n8606), .QN(n20518)
         );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6082), .CK(CLK), .Q(n8607), .QN(n20519)
         );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6081), .CK(CLK), .Q(n8608), .QN(n20520)
         );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6080), .CK(CLK), .Q(n8609), .QN(n20521)
         );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6531), .CK(CLK), .Q(n23967), .QN(n20254)
         );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6530), .CK(CLK), .Q(n23966), .QN(n20255)
         );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6529), .CK(CLK), .Q(n23965), .QN(n20256)
         );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6528), .CK(CLK), .Q(n23964), .QN(n20257)
         );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7107), .CK(CLK), .Q(n17660), .QN(n19268)
         );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7106), .CK(CLK), .Q(n17657), .QN(n19269)
         );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7105), .CK(CLK), .Q(n17654), .QN(n19270)
         );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7104), .CK(CLK), .Q(n17651), .QN(n19271)
         );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n6847), .CK(CLK), .Q(n17649), .QN(n19336)
         );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n6846), .CK(CLK), .Q(n17646), .QN(n19337)
         );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n6845), .CK(CLK), .Q(n17643), .QN(n19338)
         );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n6844), .CK(CLK), .Q(n17640), .QN(n19339)
         );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n6843), .CK(CLK), .Q(n17637), .QN(n19340)
         );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n6842), .CK(CLK), .Q(n17634), .QN(n19341)
         );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n6841), .CK(CLK), .Q(n17631), .QN(n19342)
         );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n6840), .CK(CLK), .Q(n17628), .QN(n19343)
         );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n6839), .CK(CLK), .Q(n17538), .QN(n19344)
         );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n6838), .CK(CLK), .Q(n17535), .QN(n19345)
         );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n6837), .CK(CLK), .Q(n17532), .QN(n19346)
         );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n6836), .CK(CLK), .Q(n17529), .QN(n19347)
         );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n6835), .CK(CLK), .Q(n17526), .QN(n19348)
         );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n6834), .CK(CLK), .Q(n17523), .QN(n19349)
         );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n6833), .CK(CLK), .Q(n17520), .QN(n19350)
         );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n6832), .CK(CLK), .Q(n17517), .QN(n19351)
         );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n6831), .CK(CLK), .Q(n17514), .QN(n19352)
         );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n6830), .CK(CLK), .Q(n17511), .QN(n19353)
         );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n6829), .CK(CLK), .Q(n17508), .QN(n19354)
         );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n6828), .CK(CLK), .Q(n17505), .QN(n19355)
         );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n6827), .CK(CLK), .Q(n17502), .QN(n19356)
         );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n6826), .CK(CLK), .Q(n17499), .QN(n19357)
         );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n6825), .CK(CLK), .Q(n17496), .QN(n19358)
         );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n6824), .CK(CLK), .Q(n17493), .QN(n19359)
         );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n6823), .CK(CLK), .Q(n17490), .QN(n19360)
         );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n6822), .CK(CLK), .Q(n17487), .QN(n19361)
         );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n6821), .CK(CLK), .Q(n17484), .QN(n19362)
         );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n6820), .CK(CLK), .Q(n17481), .QN(n19363)
         );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n6819), .CK(CLK), .Q(n17478), .QN(n19364)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n6818), .CK(CLK), .Q(n17475), .QN(n19365)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n6817), .CK(CLK), .Q(n17472), .QN(n19366)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n6816), .CK(CLK), .Q(n17625), .QN(n19367)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n6815), .CK(CLK), .Q(n17622), .QN(n19368)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n6814), .CK(CLK), .Q(n17619), .QN(n19369)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n6813), .CK(CLK), .Q(n17616), .QN(n19370)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n6812), .CK(CLK), .Q(n17613), .QN(n19371)
         );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n5759), .CK(CLK), .Q(n8482), .QN(n21015)
         );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n5758), .CK(CLK), .Q(n8483), .QN(n21016)
         );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n5757), .CK(CLK), .Q(n8484), .QN(n21017)
         );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n5756), .CK(CLK), .Q(n8485), .QN(n21018)
         );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n5755), .CK(CLK), .Q(n8486), .QN(n21019)
         );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n5754), .CK(CLK), .Q(n8487), .QN(n21020)
         );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n5753), .CK(CLK), .Q(n8488), .QN(n21021)
         );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n5752), .CK(CLK), .Q(n8489), .QN(n21022)
         );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n5751), .CK(CLK), .Q(n8490), .QN(n21023)
         );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n5750), .CK(CLK), .Q(n8491), .QN(n21024)
         );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n5749), .CK(CLK), .Q(n8492), .QN(n21025)
         );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n5748), .CK(CLK), .Q(n8493), .QN(n21026)
         );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n5747), .CK(CLK), .Q(n8494), .QN(n21027)
         );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n5746), .CK(CLK), .Q(n8495), .QN(n21028)
         );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n5745), .CK(CLK), .Q(n8496), .QN(n21029)
         );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n5744), .CK(CLK), .Q(n8497), .QN(n21030)
         );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n5743), .CK(CLK), .Q(n8498), .QN(n21031)
         );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n5742), .CK(CLK), .Q(n8499), .QN(n21032)
         );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n5741), .CK(CLK), .Q(n8500), .QN(n21033)
         );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n5740), .CK(CLK), .Q(n8501), .QN(n21034)
         );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n5739), .CK(CLK), .Q(n8502), .QN(n21035)
         );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n5738), .CK(CLK), .Q(n8503), .QN(n21036)
         );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n5737), .CK(CLK), .Q(n8504), .QN(n21037)
         );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n5736), .CK(CLK), .Q(n8505), .QN(n21038)
         );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n5735), .CK(CLK), .Q(n8506), .QN(n21039)
         );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n5734), .CK(CLK), .Q(n8507), .QN(n21040)
         );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n5733), .CK(CLK), .Q(n8508), .QN(n21041)
         );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n5732), .CK(CLK), .Q(n8509), .QN(n21042)
         );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n5731), .CK(CLK), .Q(n8510), .QN(n21043)
         );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n5730), .CK(CLK), .Q(n8511), .QN(n21044)
         );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n5729), .CK(CLK), .Q(n8512), .QN(n21045)
         );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n5728), .CK(CLK), .Q(n8513), .QN(n21046)
         );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n5727), .CK(CLK), .Q(n8514), .QN(n21047)
         );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n5726), .CK(CLK), .Q(n8515), .QN(n21048)
         );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n5725), .CK(CLK), .Q(n8516), .QN(n21049)
         );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n5724), .CK(CLK), .Q(n8517), .QN(n21050)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n6811), .CK(CLK), .Q(n17610), .QN(n19372)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n6810), .CK(CLK), .Q(n17607), .QN(n19373)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n6809), .CK(CLK), .Q(n17604), .QN(n19374)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n6808), .CK(CLK), .Q(n17601), .QN(n19375)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n6807), .CK(CLK), .Q(n17598), .QN(n19376)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n6806), .CK(CLK), .Q(n17595), .QN(n19377)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n6805), .CK(CLK), .Q(n17592), .QN(n19378)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n6804), .CK(CLK), .Q(n17589), .QN(n19379)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n6803), .CK(CLK), .Q(n17586), .QN(n19380)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n6802), .CK(CLK), .Q(n17583), .QN(n19381)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n6801), .CK(CLK), .Q(n17580), .QN(n19382)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n6800), .CK(CLK), .Q(n17577), .QN(n19383)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n6799), .CK(CLK), .Q(n17574), .QN(n19384)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n6798), .CK(CLK), .Q(n17571), .QN(n19385)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n6797), .CK(CLK), .Q(n17568), .QN(n19386)
         );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n6796), .CK(CLK), .Q(n17565), .QN(n19387)
         );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n6795), .CK(CLK), .Q(n17562), .QN(n19388)
         );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n6794), .CK(CLK), .Q(n17559), .QN(n19389)
         );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n6793), .CK(CLK), .Q(n17556), .QN(n19390)
         );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n6792), .CK(CLK), .Q(n17553), .QN(n19391)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n6791), .CK(CLK), .Q(n17550), .QN(n19392)
         );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n6790), .CK(CLK), .Q(n17547), .QN(n19393)
         );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n6789), .CK(CLK), .Q(n17544), .QN(n19394)
         );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n6788), .CK(CLK), .Q(n17541), .QN(n19395)
         );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6339), .CK(CLK), .Q(n8286), .QN(n20531)
         );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6338), .CK(CLK), .Q(n8287), .QN(n20532)
         );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6337), .CK(CLK), .Q(n8288), .QN(n20533)
         );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6336), .CK(CLK), .Q(n8289), .QN(n20534)
         );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6595), .CK(CLK), .Q(n8030), .QN(n20535)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6594), .CK(CLK), .Q(n8031), .QN(n20536)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6593), .CK(CLK), .Q(n8032), .QN(n20537)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6592), .CK(CLK), .Q(n8033), .QN(n20538)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n5723), .CK(CLK), .Q(n8518), .QN(n21123)
         );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n5722), .CK(CLK), .Q(n8519), .QN(n21124)
         );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n5721), .CK(CLK), .Q(n8520), .QN(n21125)
         );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n5720), .CK(CLK), .Q(n8521), .QN(n21126)
         );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n5719), .CK(CLK), .Q(n8522), .QN(n21127)
         );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n5718), .CK(CLK), .Q(n8523), .QN(n21128)
         );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n5717), .CK(CLK), .Q(n8524), .QN(n21129)
         );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n5716), .CK(CLK), .Q(n8525), .QN(n21130)
         );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n5715), .CK(CLK), .Q(n8526), .QN(n21131)
         );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n5714), .CK(CLK), .Q(n8527), .QN(n21132)
         );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n5713), .CK(CLK), .Q(n8528), .QN(n21133)
         );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n5712), .CK(CLK), .Q(n8529), .QN(n21134)
         );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n5711), .CK(CLK), .Q(n8530), .QN(n21135)
         );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n5710), .CK(CLK), .Q(n8531), .QN(n21136)
         );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n5709), .CK(CLK), .Q(n8532), .QN(n21137)
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n5708), .CK(CLK), .Q(n8533), .QN(n21138)
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n5707), .CK(CLK), .Q(n8534), .QN(n21139)
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n5706), .CK(CLK), .Q(n8535), .QN(n21140)
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n5705), .CK(CLK), .Q(n8536), .QN(n21141)
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n5704), .CK(CLK), .Q(n8537), .QN(n21142)
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n5703), .CK(CLK), .Q(n8538), .QN(n21143)
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n5702), .CK(CLK), .Q(n8539), .QN(n21144)
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n5701), .CK(CLK), .Q(n8540), .QN(n21145)
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n5700), .CK(CLK), .Q(n8541), .QN(n21146)
         );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5315), .CK(CLK), .Q(n24031), .QN(n20145) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5314), .CK(CLK), .Q(n24030), .QN(n20146) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5313), .CK(CLK), .Q(n24029), .QN(n20147) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5312), .CK(CLK), .Q(n24028), .QN(n20148) );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5187), .CK(CLK), .Q(n8670), .QN(n20506)
         );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5186), .CK(CLK), .Q(n8671), .QN(n20507)
         );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5185), .CK(CLK), .Q(n8672), .QN(n20508)
         );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5184), .CK(CLK), .Q(n8673), .QN(n20509)
         );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5443), .CK(CLK), .Q(n8350), .QN(n20510)
         );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5442), .CK(CLK), .Q(n8351), .QN(n20511)
         );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5441), .CK(CLK), .Q(n8352), .QN(n20512)
         );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5440), .CK(CLK), .Q(n8353), .QN(n20513)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n6981), .CK(CLK), .Q(n7708), .QN(n21147)
         );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6079), .CK(CLK), .Q(n8610), .QN(n20655)
         );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6078), .CK(CLK), .Q(n8611), .QN(n20656)
         );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6077), .CK(CLK), .Q(n8612), .QN(n20657)
         );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6076), .CK(CLK), .Q(n8613), .QN(n20658)
         );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6075), .CK(CLK), .Q(n8614), .QN(n20659)
         );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6074), .CK(CLK), .Q(n8615), .QN(n20660)
         );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6073), .CK(CLK), .Q(n8616), .QN(n20661)
         );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6072), .CK(CLK), .Q(n8617), .QN(n20662)
         );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6071), .CK(CLK), .Q(n8618), .QN(n20663)
         );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6070), .CK(CLK), .Q(n8619), .QN(n20664)
         );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n6069), .CK(CLK), .Q(n8620), .QN(n20665)
         );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n6068), .CK(CLK), .Q(n8621), .QN(n20666)
         );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n6067), .CK(CLK), .Q(n8622), .QN(n20667)
         );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n6066), .CK(CLK), .Q(n8623), .QN(n20668)
         );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n6065), .CK(CLK), .Q(n8624), .QN(n20669)
         );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n6064), .CK(CLK), .Q(n8625), .QN(n20670)
         );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n6063), .CK(CLK), .Q(n8626), .QN(n20671)
         );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n6062), .CK(CLK), .Q(n8627), .QN(n20672)
         );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n6061), .CK(CLK), .Q(n8628), .QN(n20673)
         );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n6060), .CK(CLK), .Q(n8629), .QN(n20674)
         );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n6059), .CK(CLK), .Q(n8630), .QN(n20675)
         );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n6058), .CK(CLK), .Q(n8631), .QN(n20676)
         );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n6057), .CK(CLK), .Q(n8632), .QN(n20677)
         );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n6056), .CK(CLK), .Q(n8633), .QN(n20678)
         );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n6055), .CK(CLK), .Q(n8634), .QN(n20679)
         );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n6054), .CK(CLK), .Q(n8635), .QN(n20680)
         );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n6053), .CK(CLK), .Q(n8636), .QN(n20681)
         );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n6052), .CK(CLK), .Q(n8637), .QN(n20682)
         );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n6051), .CK(CLK), .Q(n8638), .QN(n20683)
         );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n6050), .CK(CLK), .Q(n8639), .QN(n20684)
         );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n6049), .CK(CLK), .Q(n8640), .QN(n20685)
         );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n6048), .CK(CLK), .Q(n8641), .QN(n20686)
         );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n6047), .CK(CLK), .Q(n8642), .QN(n20687)
         );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n6046), .CK(CLK), .Q(n8643), .QN(n20688)
         );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n6045), .CK(CLK), .Q(n8644), .QN(n20689)
         );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n6044), .CK(CLK), .Q(n8645), .QN(n20690)
         );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6527), .CK(CLK), .Q(n23963), .QN(n20302)
         );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6526), .CK(CLK), .Q(n23962), .QN(n20303)
         );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6525), .CK(CLK), .Q(n23961), .QN(n20304)
         );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6524), .CK(CLK), .Q(n23960), .QN(n20305)
         );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6523), .CK(CLK), .Q(n23959), .QN(n20306)
         );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6522), .CK(CLK), .Q(n23958), .QN(n20307)
         );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6521), .CK(CLK), .Q(n23957), .QN(n20308)
         );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6520), .CK(CLK), .Q(n23956), .QN(n20309)
         );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6519), .CK(CLK), .Q(n23955), .QN(n20310)
         );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6518), .CK(CLK), .Q(n23954), .QN(n20311)
         );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6517), .CK(CLK), .Q(n23953), .QN(n20312)
         );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6516), .CK(CLK), .Q(n23952), .QN(n20313)
         );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6515), .CK(CLK), .Q(n23950), .QN(n20314)
         );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6514), .CK(CLK), .Q(n23948), .QN(n20315)
         );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6513), .CK(CLK), .Q(n23946), .QN(n20316)
         );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6512), .CK(CLK), .Q(n23944), .QN(n20317)
         );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6511), .CK(CLK), .Q(n23942), .QN(n20318)
         );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6510), .CK(CLK), .Q(n23940), .QN(n20319)
         );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6509), .CK(CLK), .Q(n23938), .QN(n20320)
         );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6508), .CK(CLK), .Q(n23936), .QN(n20321)
         );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6507), .CK(CLK), .Q(n23934), .QN(n20322)
         );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6506), .CK(CLK), .Q(n23932), .QN(n20323)
         );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6505), .CK(CLK), .Q(n23930), .QN(n20324)
         );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6504), .CK(CLK), .Q(n23928), .QN(n20325)
         );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6503), .CK(CLK), .Q(n23926), .QN(n20326)
         );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6502), .CK(CLK), .Q(n23924), .QN(n20327)
         );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6501), .CK(CLK), .Q(n23922), .QN(n20328)
         );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6500), .CK(CLK), .Q(n23920), .QN(n20329)
         );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6499), .CK(CLK), .Q(n23918), .QN(n20330)
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6498), .CK(CLK), .Q(n23916), .QN(n20331)
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6497), .CK(CLK), .Q(n23914), .QN(n20332)
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6496), .CK(CLK), .Q(n23912), .QN(n20333)
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6495), .CK(CLK), .Q(n23910), .QN(n20334)
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6494), .CK(CLK), .Q(n23908), .QN(n20335)
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6493), .CK(CLK), .Q(n23906), .QN(n20336)
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6492), .CK(CLK), .Q(n23904), .QN(n20337)
         );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n6043), .CK(CLK), .Q(n8646), .QN(n20799)
         );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n6042), .CK(CLK), .Q(n8647), .QN(n20800)
         );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n6041), .CK(CLK), .Q(n8648), .QN(n20801)
         );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n6040), .CK(CLK), .Q(n8649), .QN(n20802)
         );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n6039), .CK(CLK), .Q(n8650), .QN(n20803)
         );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n6038), .CK(CLK), .Q(n8651), .QN(n20804)
         );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n6037), .CK(CLK), .Q(n8652), .QN(n20805)
         );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n6036), .CK(CLK), .Q(n8653), .QN(n20806)
         );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n6035), .CK(CLK), .Q(n8654), .QN(n20807)
         );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n6034), .CK(CLK), .Q(n8655), .QN(n20808)
         );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n6033), .CK(CLK), .Q(n8656), .QN(n20809)
         );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n6032), .CK(CLK), .Q(n8657), .QN(n20810)
         );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n6031), .CK(CLK), .Q(n8658), .QN(n20811)
         );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n6030), .CK(CLK), .Q(n8659), .QN(n20812)
         );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n6029), .CK(CLK), .Q(n8660), .QN(n20813)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n6028), .CK(CLK), .Q(n8661), .QN(n20814)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n6027), .CK(CLK), .Q(n8662), .QN(n20815)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n6026), .CK(CLK), .Q(n8663), .QN(n20816)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n6025), .CK(CLK), .Q(n8664), .QN(n20817)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n6024), .CK(CLK), .Q(n8665), .QN(n20818)
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n6023), .CK(CLK), .Q(n8666), .QN(n20819)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n6022), .CK(CLK), .Q(n8667), .QN(n20820)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n6021), .CK(CLK), .Q(n8668), .QN(n20821)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n6020), .CK(CLK), .Q(n8669), .QN(n20822)
         );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7103), .CK(CLK), .Q(n17648), .QN(n19272)
         );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7102), .CK(CLK), .Q(n17645), .QN(n19273)
         );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7101), .CK(CLK), .Q(n17642), .QN(n19274)
         );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7100), .CK(CLK), .Q(n17639), .QN(n19275)
         );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7099), .CK(CLK), .Q(n17636), .QN(n19276)
         );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7098), .CK(CLK), .Q(n17633), .QN(n19277)
         );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7097), .CK(CLK), .Q(n17630), .QN(n19278)
         );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7096), .CK(CLK), .Q(n17627), .QN(n19279)
         );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7095), .CK(CLK), .Q(n17537), .QN(n19280)
         );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7094), .CK(CLK), .Q(n17534), .QN(n19281)
         );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7093), .CK(CLK), .Q(n17531), .QN(n19282)
         );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7092), .CK(CLK), .Q(n17528), .QN(n19283)
         );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7091), .CK(CLK), .Q(n17525), .QN(n19284)
         );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7090), .CK(CLK), .Q(n17522), .QN(n19285)
         );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7089), .CK(CLK), .Q(n17519), .QN(n19286)
         );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7088), .CK(CLK), .Q(n17516), .QN(n19287)
         );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7087), .CK(CLK), .Q(n17513), .QN(n19288)
         );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7086), .CK(CLK), .Q(n17510), .QN(n19289)
         );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7085), .CK(CLK), .Q(n17507), .QN(n19290)
         );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7084), .CK(CLK), .Q(n17504), .QN(n19291)
         );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7083), .CK(CLK), .Q(n17501), .QN(n19292)
         );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7082), .CK(CLK), .Q(n17498), .QN(n19293)
         );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7081), .CK(CLK), .Q(n17495), .QN(n19294)
         );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7080), .CK(CLK), .Q(n17492), .QN(n19295)
         );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7079), .CK(CLK), .Q(n17489), .QN(n19296)
         );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7078), .CK(CLK), .Q(n17486), .QN(n19297)
         );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7077), .CK(CLK), .Q(n17483), .QN(n19298)
         );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7076), .CK(CLK), .Q(n17480), .QN(n19299)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7075), .CK(CLK), .Q(n17477), .QN(n19300)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7074), .CK(CLK), .Q(n17474), .QN(n19301)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7073), .CK(CLK), .Q(n17471), .QN(n19302)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7072), .CK(CLK), .Q(n17624), .QN(n19303)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7071), .CK(CLK), .Q(n17621), .QN(n19304)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7070), .CK(CLK), .Q(n17618), .QN(n19305)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7069), .CK(CLK), .Q(n17615), .QN(n19306)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7068), .CK(CLK), .Q(n17612), .QN(n19307)
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6491), .CK(CLK), .Q(n23902), .QN(n20398)
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6490), .CK(CLK), .Q(n23900), .QN(n20399)
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6489), .CK(CLK), .Q(n23898), .QN(n20400)
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6488), .CK(CLK), .Q(n23896), .QN(n20401)
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6487), .CK(CLK), .Q(n23894), .QN(n20402)
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6486), .CK(CLK), .Q(n23892), .QN(n20403)
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6485), .CK(CLK), .Q(n23890), .QN(n20404)
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6484), .CK(CLK), .Q(n23888), .QN(n20405)
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6483), .CK(CLK), .Q(n23886), .QN(n20406)
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6482), .CK(CLK), .Q(n23884), .QN(n20407)
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6481), .CK(CLK), .Q(n23882), .QN(n20408)
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6480), .CK(CLK), .Q(n23880), .QN(n20409)
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6479), .CK(CLK), .Q(n23878), .QN(n20410)
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6478), .CK(CLK), .Q(n23876), .QN(n20411)
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6477), .CK(CLK), .Q(n23874), .QN(n20412)
         );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6476), .CK(CLK), .Q(n23872), .QN(n20413)
         );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6475), .CK(CLK), .Q(n23870), .QN(n20414)
         );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6474), .CK(CLK), .Q(n23868), .QN(n20415)
         );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6473), .CK(CLK), .Q(n23866), .QN(n20416)
         );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6472), .CK(CLK), .Q(n23864), .QN(n20417)
         );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6471), .CK(CLK), .Q(n23862), .QN(n20418)
         );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6470), .CK(CLK), .Q(n23860), .QN(n20419)
         );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6469), .CK(CLK), .Q(n23858), .QN(n20420)
         );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6468), .CK(CLK), .Q(n23856), .QN(n20421)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7067), .CK(CLK), .Q(n17609), .QN(n19308)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7066), .CK(CLK), .Q(n17606), .QN(n19309)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7065), .CK(CLK), .Q(n17603), .QN(n19310)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7064), .CK(CLK), .Q(n17600), .QN(n19311)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7063), .CK(CLK), .Q(n17597), .QN(n19312)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7062), .CK(CLK), .Q(n17594), .QN(n19313)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7061), .CK(CLK), .Q(n17591), .QN(n19314)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7060), .CK(CLK), .Q(n17588), .QN(n19315)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7059), .CK(CLK), .Q(n17585), .QN(n19316)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7058), .CK(CLK), .Q(n17582), .QN(n19317)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7057), .CK(CLK), .Q(n17579), .QN(n19318)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7056), .CK(CLK), .Q(n17576), .QN(n19319)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n7055), .CK(CLK), .Q(n17573), .QN(n19320)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n7054), .CK(CLK), .Q(n17570), .QN(n19321)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n7053), .CK(CLK), .Q(n17567), .QN(n19322)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n7052), .CK(CLK), .Q(n17564), .QN(n19323)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n7051), .CK(CLK), .Q(n17561), .QN(n19324)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n7050), .CK(CLK), .Q(n17558), .QN(n19325)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n7049), .CK(CLK), .Q(n17555), .QN(n19326)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n7048), .CK(CLK), .Q(n17552), .QN(n19327)
         );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n7047), .CK(CLK), .Q(n17549), .QN(n19328)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n7046), .CK(CLK), .Q(n17546), .QN(n19329)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n7045), .CK(CLK), .Q(n17543), .QN(n19330)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n7044), .CK(CLK), .Q(n17540), .QN(n19331)
         );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6335), .CK(CLK), .Q(n8290), .QN(n20907)
         );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6334), .CK(CLK), .Q(n8291), .QN(n20908)
         );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6333), .CK(CLK), .Q(n8292), .QN(n20909)
         );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6332), .CK(CLK), .Q(n8293), .QN(n20910)
         );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6331), .CK(CLK), .Q(n8294), .QN(n20911)
         );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6330), .CK(CLK), .Q(n8295), .QN(n20912)
         );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6329), .CK(CLK), .Q(n8296), .QN(n20913)
         );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6328), .CK(CLK), .Q(n8297), .QN(n20914)
         );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6327), .CK(CLK), .Q(n8298), .QN(n20915)
         );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6326), .CK(CLK), .Q(n8299), .QN(n20916)
         );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6325), .CK(CLK), .Q(n8300), .QN(n20917)
         );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6324), .CK(CLK), .Q(n8301), .QN(n20918)
         );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6323), .CK(CLK), .Q(n8302), .QN(n20919)
         );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6322), .CK(CLK), .Q(n8303), .QN(n20920)
         );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6321), .CK(CLK), .Q(n8304), .QN(n20921)
         );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6320), .CK(CLK), .Q(n8305), .QN(n20922)
         );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6319), .CK(CLK), .Q(n8306), .QN(n20923)
         );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6318), .CK(CLK), .Q(n8307), .QN(n20924)
         );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6317), .CK(CLK), .Q(n8308), .QN(n20925)
         );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6316), .CK(CLK), .Q(n8309), .QN(n20926)
         );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6315), .CK(CLK), .Q(n8310), .QN(n20927)
         );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6314), .CK(CLK), .Q(n8311), .QN(n20928)
         );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6313), .CK(CLK), .Q(n8312), .QN(n20929)
         );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6312), .CK(CLK), .Q(n8313), .QN(n20930)
         );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6311), .CK(CLK), .Q(n8314), .QN(n20931)
         );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6310), .CK(CLK), .Q(n8315), .QN(n20932)
         );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6309), .CK(CLK), .Q(n8316), .QN(n20933)
         );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6308), .CK(CLK), .Q(n8317), .QN(n20934)
         );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6307), .CK(CLK), .Q(n8318), .QN(n20935)
         );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6306), .CK(CLK), .Q(n8319), .QN(n20936)
         );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6305), .CK(CLK), .Q(n8320), .QN(n20937)
         );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6304), .CK(CLK), .Q(n8321), .QN(n20938)
         );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6303), .CK(CLK), .Q(n8322), .QN(n20939)
         );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6302), .CK(CLK), .Q(n8323), .QN(n20940)
         );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6301), .CK(CLK), .Q(n8324), .QN(n20941)
         );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6300), .CK(CLK), .Q(n8325), .QN(n20942)
         );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6591), .CK(CLK), .Q(n8034), .QN(n20943)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6590), .CK(CLK), .Q(n8035), .QN(n20944)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6589), .CK(CLK), .Q(n8036), .QN(n20945)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6588), .CK(CLK), .Q(n8037), .QN(n20946)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6587), .CK(CLK), .Q(n8038), .QN(n20947)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6586), .CK(CLK), .Q(n8039), .QN(n20948)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6585), .CK(CLK), .Q(n8040), .QN(n20949)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6584), .CK(CLK), .Q(n8041), .QN(n20950)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6583), .CK(CLK), .Q(n8042), .QN(n20951)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6582), .CK(CLK), .Q(n8043), .QN(n20952)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6581), .CK(CLK), .Q(n8044), .QN(n20953)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6580), .CK(CLK), .Q(n8045), .QN(n20954)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6579), .CK(CLK), .Q(n8046), .QN(n20955)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6578), .CK(CLK), .Q(n8047), .QN(n20956)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6577), .CK(CLK), .Q(n8048), .QN(n20957)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6576), .CK(CLK), .Q(n8049), .QN(n20958)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6575), .CK(CLK), .Q(n8050), .QN(n20959)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6574), .CK(CLK), .Q(n8051), .QN(n20960)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6573), .CK(CLK), .Q(n8052), .QN(n20961)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6572), .CK(CLK), .Q(n8053), .QN(n20962)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6571), .CK(CLK), .Q(n8054), .QN(n20963)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6570), .CK(CLK), .Q(n8055), .QN(n20964)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6569), .CK(CLK), .Q(n8056), .QN(n20965)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6568), .CK(CLK), .Q(n8057), .QN(n20966)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6567), .CK(CLK), .Q(n8058), .QN(n20967)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6566), .CK(CLK), .Q(n8059), .QN(n20968)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6565), .CK(CLK), .Q(n8060), .QN(n20969)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6564), .CK(CLK), .Q(n8061), .QN(n20970)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6563), .CK(CLK), .Q(n8062), .QN(n20971)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6562), .CK(CLK), .Q(n8063), .QN(n20972)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6561), .CK(CLK), .Q(n8064), .QN(n20973)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6560), .CK(CLK), .Q(n8065), .QN(n20974)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6559), .CK(CLK), .Q(n8066), .QN(n20975)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6558), .CK(CLK), .Q(n8067), .QN(n20976)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6557), .CK(CLK), .Q(n8068), .QN(n20977)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6556), .CK(CLK), .Q(n8069), .QN(n20978)
         );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5311), .CK(CLK), .Q(n24027), .QN(n20157) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5310), .CK(CLK), .Q(n24026), .QN(n20158) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5309), .CK(CLK), .Q(n24025), .QN(n20159) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5308), .CK(CLK), .Q(n24024), .QN(n20160) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5307), .CK(CLK), .Q(n24023), .QN(n20161) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5306), .CK(CLK), .Q(n24022), .QN(n20162) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5305), .CK(CLK), .Q(n24021), .QN(n20163) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5304), .CK(CLK), .Q(n24020), .QN(n20164) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5303), .CK(CLK), .Q(n24019), .QN(n20165) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5302), .CK(CLK), .Q(n24018), .QN(n20166) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5301), .CK(CLK), .Q(n24017), .QN(n20167) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5300), .CK(CLK), .Q(n24016), .QN(n20168) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5299), .CK(CLK), .Q(n24015), .QN(n20169) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5298), .CK(CLK), .Q(n24014), .QN(n20170) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5297), .CK(CLK), .Q(n24013), .QN(n20171) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5296), .CK(CLK), .Q(n24012), .QN(n20172) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5295), .CK(CLK), .Q(n24011), .QN(n20173) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5294), .CK(CLK), .Q(n24010), .QN(n20174) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5293), .CK(CLK), .Q(n24009), .QN(n20175) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5292), .CK(CLK), .Q(n24008), .QN(n20176) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5291), .CK(CLK), .Q(n24007), .QN(n20177) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5290), .CK(CLK), .Q(n24006), .QN(n20178) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5289), .CK(CLK), .Q(n24005), .QN(n20179) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5288), .CK(CLK), .Q(n24004), .QN(n20180) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5287), .CK(CLK), .Q(n24003), .QN(n20181) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5286), .CK(CLK), .Q(n24002), .QN(n20182) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5285), .CK(CLK), .Q(n24001), .QN(n20183) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5284), .CK(CLK), .Q(n24000), .QN(n20184) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5283), .CK(CLK), .Q(n23999), .QN(n20185) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5282), .CK(CLK), .Q(n23998), .QN(n20186) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5281), .CK(CLK), .Q(n23997), .QN(n19708) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5280), .CK(CLK), .Q(n23996), .QN(n19709) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5279), .CK(CLK), .Q(n23995), .QN(n19710) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5278), .CK(CLK), .Q(n23994), .QN(n19711) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5277), .CK(CLK), .Q(n23993), .QN(n19712) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5276), .CK(CLK), .Q(n23992), .QN(n19713) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6299), .CK(CLK), .Q(n8326), .QN(n21051)
         );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6298), .CK(CLK), .Q(n8327), .QN(n21052)
         );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6297), .CK(CLK), .Q(n8328), .QN(n21053)
         );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6296), .CK(CLK), .Q(n8329), .QN(n21054)
         );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6295), .CK(CLK), .Q(n8330), .QN(n21055)
         );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6294), .CK(CLK), .Q(n8331), .QN(n21056)
         );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6293), .CK(CLK), .Q(n8332), .QN(n21057)
         );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6292), .CK(CLK), .Q(n8333), .QN(n21058)
         );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6291), .CK(CLK), .Q(n8334), .QN(n21059)
         );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6290), .CK(CLK), .Q(n8335), .QN(n21060)
         );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6289), .CK(CLK), .Q(n8336), .QN(n21061)
         );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6288), .CK(CLK), .Q(n8337), .QN(n21062)
         );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6287), .CK(CLK), .Q(n8338), .QN(n21063)
         );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6286), .CK(CLK), .Q(n8339), .QN(n21064)
         );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6285), .CK(CLK), .Q(n8340), .QN(n21065)
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6284), .CK(CLK), .Q(n8341), .QN(n21066)
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6283), .CK(CLK), .Q(n8342), .QN(n21067)
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6282), .CK(CLK), .Q(n8343), .QN(n21068)
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6281), .CK(CLK), .Q(n8344), .QN(n21069)
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6280), .CK(CLK), .Q(n8345), .QN(n21070)
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6279), .CK(CLK), .Q(n8346), .QN(n21071)
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6278), .CK(CLK), .Q(n8347), .QN(n21072)
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6277), .CK(CLK), .Q(n8348), .QN(n21073)
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6276), .CK(CLK), .Q(n8349), .QN(n21074)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6555), .CK(CLK), .Q(n8070), .QN(n21075)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6554), .CK(CLK), .Q(n8071), .QN(n21076)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6553), .CK(CLK), .Q(n8072), .QN(n21077)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6552), .CK(CLK), .Q(n8073), .QN(n21078)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6551), .CK(CLK), .Q(n8074), .QN(n21079)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6550), .CK(CLK), .Q(n8075), .QN(n21080)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6549), .CK(CLK), .Q(n8076), .QN(n21081)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6548), .CK(CLK), .Q(n8077), .QN(n21082)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6547), .CK(CLK), .Q(n8078), .QN(n21083)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6546), .CK(CLK), .Q(n8079), .QN(n21084)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6545), .CK(CLK), .Q(n8080), .QN(n21085)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6544), .CK(CLK), .Q(n8081), .QN(n21086)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6543), .CK(CLK), .Q(n8082), .QN(n21087)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6542), .CK(CLK), .Q(n8083), .QN(n21088)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6541), .CK(CLK), .Q(n8084), .QN(n21089)
         );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6540), .CK(CLK), .Q(n8085), .QN(n21090)
         );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6539), .CK(CLK), .Q(n8086), .QN(n21091)
         );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6538), .CK(CLK), .Q(n8087), .QN(n21092)
         );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6537), .CK(CLK), .Q(n8088), .QN(n21093)
         );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6536), .CK(CLK), .Q(n8089), .QN(n21094)
         );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6535), .CK(CLK), .Q(n8090), .QN(n21095)
         );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6534), .CK(CLK), .Q(n8091), .QN(n21096)
         );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6533), .CK(CLK), .Q(n8092), .QN(n21097)
         );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6532), .CK(CLK), .Q(n8093), .QN(n21098)
         );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5183), .CK(CLK), .Q(n8674), .QN(n20547)
         );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5182), .CK(CLK), .Q(n8675), .QN(n20548)
         );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5181), .CK(CLK), .Q(n8676), .QN(n20549)
         );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5180), .CK(CLK), .Q(n8677), .QN(n20550)
         );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5179), .CK(CLK), .Q(n8678), .QN(n20551)
         );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5178), .CK(CLK), .Q(n8679), .QN(n20552)
         );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5177), .CK(CLK), .Q(n8680), .QN(n20553)
         );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5176), .CK(CLK), .Q(n8681), .QN(n20554)
         );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5175), .CK(CLK), .Q(n8682), .QN(n20555)
         );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5174), .CK(CLK), .Q(n8683), .QN(n20556)
         );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5173), .CK(CLK), .Q(n8684), .QN(n20557)
         );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5172), .CK(CLK), .Q(n8685), .QN(n20558)
         );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5171), .CK(CLK), .Q(n8686), .QN(n20559)
         );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5170), .CK(CLK), .Q(n8687), .QN(n20560)
         );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5169), .CK(CLK), .Q(n8688), .QN(n20561)
         );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5168), .CK(CLK), .Q(n8689), .QN(n20562)
         );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5167), .CK(CLK), .Q(n8690), .QN(n20563)
         );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5166), .CK(CLK), .Q(n8691), .QN(n20564)
         );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5165), .CK(CLK), .Q(n8692), .QN(n20565)
         );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5164), .CK(CLK), .Q(n8693), .QN(n20566)
         );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5163), .CK(CLK), .Q(n8694), .QN(n20567)
         );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5162), .CK(CLK), .Q(n8695), .QN(n20568)
         );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5161), .CK(CLK), .Q(n8696), .QN(n20569)
         );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5160), .CK(CLK), .Q(n8697), .QN(n20570)
         );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5159), .CK(CLK), .Q(n8698), .QN(n20571)
         );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5158), .CK(CLK), .Q(n8699), .QN(n20572)
         );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5157), .CK(CLK), .Q(n8700), .QN(n20573)
         );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5156), .CK(CLK), .Q(n8701), .QN(n20574)
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5155), .CK(CLK), .Q(n8702), .QN(n20575)
         );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5154), .CK(CLK), .Q(n8703), .QN(n20576)
         );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5153), .CK(CLK), .Q(n8704), .QN(n20577)
         );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5152), .CK(CLK), .Q(n8705), .QN(n20578)
         );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5151), .CK(CLK), .Q(n8706), .QN(n20579)
         );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5150), .CK(CLK), .Q(n8707), .QN(n20580)
         );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5149), .CK(CLK), .Q(n8708), .QN(n20581)
         );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5148), .CK(CLK), .Q(n8709), .QN(n20582)
         );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5439), .CK(CLK), .Q(n8354), .QN(n20583)
         );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5438), .CK(CLK), .Q(n8355), .QN(n20584)
         );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5437), .CK(CLK), .Q(n8356), .QN(n20585)
         );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5436), .CK(CLK), .Q(n8357), .QN(n20586)
         );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5435), .CK(CLK), .Q(n8358), .QN(n20587)
         );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5434), .CK(CLK), .Q(n8359), .QN(n20588)
         );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5433), .CK(CLK), .Q(n8360), .QN(n20589)
         );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5432), .CK(CLK), .Q(n8361), .QN(n20590)
         );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5431), .CK(CLK), .Q(n8362), .QN(n20591)
         );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5430), .CK(CLK), .Q(n8363), .QN(n20592)
         );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5429), .CK(CLK), .Q(n8364), .QN(n20593)
         );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5428), .CK(CLK), .Q(n8365), .QN(n20594)
         );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5427), .CK(CLK), .Q(n8366), .QN(n20595)
         );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5426), .CK(CLK), .Q(n8367), .QN(n20596)
         );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5425), .CK(CLK), .Q(n8368), .QN(n20597)
         );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5424), .CK(CLK), .Q(n8369), .QN(n20598)
         );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5423), .CK(CLK), .Q(n8370), .QN(n20599)
         );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5422), .CK(CLK), .Q(n8371), .QN(n20600)
         );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5421), .CK(CLK), .Q(n8372), .QN(n20601)
         );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5420), .CK(CLK), .Q(n8373), .QN(n20602)
         );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5419), .CK(CLK), .Q(n8374), .QN(n20603)
         );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5418), .CK(CLK), .Q(n8375), .QN(n20604)
         );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5417), .CK(CLK), .Q(n8376), .QN(n20605)
         );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5416), .CK(CLK), .Q(n8377), .QN(n20606)
         );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5415), .CK(CLK), .Q(n8378), .QN(n20607)
         );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5414), .CK(CLK), .Q(n8379), .QN(n20608)
         );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5413), .CK(CLK), .Q(n8380), .QN(n20609)
         );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5412), .CK(CLK), .Q(n8381), .QN(n20610)
         );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5411), .CK(CLK), .Q(n8382), .QN(n20611)
         );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5410), .CK(CLK), .Q(n8383), .QN(n20612)
         );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5409), .CK(CLK), .Q(n8384), .QN(n20613)
         );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5408), .CK(CLK), .Q(n8385), .QN(n20614)
         );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5407), .CK(CLK), .Q(n8386), .QN(n20615)
         );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5406), .CK(CLK), .Q(n8387), .QN(n20616)
         );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5405), .CK(CLK), .Q(n8388), .QN(n20617)
         );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5404), .CK(CLK), .Q(n8389), .QN(n20618)
         );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5275), .CK(CLK), .Q(n23991), .QN(n19714) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5274), .CK(CLK), .Q(n23990), .QN(n19715) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5273), .CK(CLK), .Q(n23989), .QN(n19716) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5272), .CK(CLK), .Q(n23988), .QN(n19717) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5271), .CK(CLK), .Q(n23987), .QN(n19718) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5270), .CK(CLK), .Q(n23986), .QN(n19719) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5269), .CK(CLK), .Q(n23985), .QN(n19720) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5268), .CK(CLK), .Q(n23984), .QN(n19721) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5267), .CK(CLK), .Q(n23983), .QN(n19722) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5266), .CK(CLK), .Q(n23982), .QN(n19723) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5265), .CK(CLK), .Q(n23981), .QN(n19724) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5264), .CK(CLK), .Q(n23980), .QN(n19725) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5263), .CK(CLK), .Q(n23979), .QN(n19726) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5262), .CK(CLK), .Q(n23978), .QN(n19727) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5261), .CK(CLK), .Q(n23977), .QN(n19728)
         );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5260), .CK(CLK), .Q(n23976), .QN(n19729)
         );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5259), .CK(CLK), .Q(n23975), .QN(n19730)
         );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5258), .CK(CLK), .Q(n23974), .QN(n19731)
         );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5257), .CK(CLK), .Q(n23973), .QN(n19732)
         );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5256), .CK(CLK), .Q(n23972), .QN(n19733)
         );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5255), .CK(CLK), .Q(n23971), .QN(n19734)
         );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5254), .CK(CLK), .Q(n23970), .QN(n19735)
         );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5253), .CK(CLK), .Q(n23969), .QN(n19736)
         );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5252), .CK(CLK), .Q(n23968), .QN(n19737)
         );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5147), .CK(CLK), .Q(n8710), .QN(n20727)
         );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5146), .CK(CLK), .Q(n8711), .QN(n20728)
         );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5145), .CK(CLK), .Q(n8712), .QN(n20729)
         );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5144), .CK(CLK), .Q(n8713), .QN(n20730)
         );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5143), .CK(CLK), .Q(n8714), .QN(n20731)
         );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5142), .CK(CLK), .Q(n8715), .QN(n20732)
         );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5141), .CK(CLK), .Q(n8716), .QN(n20733)
         );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5140), .CK(CLK), .Q(n8717), .QN(n20734)
         );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5139), .CK(CLK), .Q(n8718), .QN(n20735)
         );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5138), .CK(CLK), .Q(n8719), .QN(n20736)
         );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5137), .CK(CLK), .Q(n8720), .QN(n20737)
         );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5136), .CK(CLK), .Q(n8721), .QN(n20738)
         );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5135), .CK(CLK), .Q(n8722), .QN(n20739)
         );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5134), .CK(CLK), .Q(n8723), .QN(n20740)
         );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5133), .CK(CLK), .Q(n8724), .QN(n20741)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5132), .CK(CLK), .Q(n8725), .QN(n20742)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5131), .CK(CLK), .Q(n8726), .QN(n20743)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5130), .CK(CLK), .Q(n8727), .QN(n20744)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5129), .CK(CLK), .Q(n8728), .QN(n20745)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5128), .CK(CLK), .Q(n8729), .QN(n20746)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5127), .CK(CLK), .Q(n8730), .QN(n20747)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5126), .CK(CLK), .Q(n8731), .QN(n20748)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5125), .CK(CLK), .Q(n8732), .QN(n20749)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5124), .CK(CLK), .Q(n8733), .QN(n20750)
         );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5403), .CK(CLK), .Q(n8390), .QN(n20751)
         );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5402), .CK(CLK), .Q(n8391), .QN(n20752)
         );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5401), .CK(CLK), .Q(n8392), .QN(n20753)
         );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5400), .CK(CLK), .Q(n8393), .QN(n20754)
         );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5399), .CK(CLK), .Q(n8394), .QN(n20755)
         );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5398), .CK(CLK), .Q(n8395), .QN(n20756)
         );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5397), .CK(CLK), .Q(n8396), .QN(n20757)
         );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5396), .CK(CLK), .Q(n8397), .QN(n20758)
         );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5395), .CK(CLK), .Q(n8398), .QN(n20759)
         );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5394), .CK(CLK), .Q(n8399), .QN(n20760)
         );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5393), .CK(CLK), .Q(n8400), .QN(n20761)
         );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5392), .CK(CLK), .Q(n8401), .QN(n20762)
         );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5391), .CK(CLK), .Q(n8402), .QN(n20763)
         );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5390), .CK(CLK), .Q(n8403), .QN(n20764)
         );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5389), .CK(CLK), .Q(n8404), .QN(n20765)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5388), .CK(CLK), .Q(n8405), .QN(n20766)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5387), .CK(CLK), .Q(n8406), .QN(n20767)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5386), .CK(CLK), .Q(n8407), .QN(n20768)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5385), .CK(CLK), .Q(n8408), .QN(n20769)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5384), .CK(CLK), .Q(n8409), .QN(n20770)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5383), .CK(CLK), .Q(n8410), .QN(n20771)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5382), .CK(CLK), .Q(n8411), .QN(n20772)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5381), .CK(CLK), .Q(n8412), .QN(n20773)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5380), .CK(CLK), .Q(n8413), .QN(n20774)
         );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n7042), .CK(CLK), .Q(n7647), .QN(n21148)
         );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n7043), .CK(CLK), .Q(n7646), .QN(n21149)
         );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7041), .CK(CLK), .Q(n7648), .QN(n21150)
         );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7040), .CK(CLK), .Q(n7649), .QN(n21151)
         );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7039), .CK(CLK), .Q(n7650), .QN(n21152)
         );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7038), .CK(CLK), .Q(n7651), .QN(n21153)
         );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7037), .CK(CLK), .Q(n7652), .QN(n21154)
         );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7036), .CK(CLK), .Q(n7653), .QN(n21155)
         );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7035), .CK(CLK), .Q(n7654), .QN(n21156)
         );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7034), .CK(CLK), .Q(n7655), .QN(n21157)
         );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7033), .CK(CLK), .Q(n7656), .QN(n21158)
         );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7032), .CK(CLK), .Q(n7657), .QN(n21159)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7008), .CK(CLK), .Q(n7681), .QN(n21160)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7007), .CK(CLK), .Q(n7682), .QN(n21161)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7006), .CK(CLK), .Q(n7683), .QN(n21162)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7005), .CK(CLK), .Q(n7684), .QN(n21163)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7004), .CK(CLK), .Q(n7685), .QN(n21164)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7003), .CK(CLK), .Q(n7686), .QN(n21165)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7002), .CK(CLK), .Q(n7687), .QN(n21166)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7001), .CK(CLK), .Q(n7688), .QN(n21167)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7000), .CK(CLK), .Q(n7689), .QN(n21168)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n6999), .CK(CLK), .Q(n7690), .QN(n21169)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n6998), .CK(CLK), .Q(n7691), .QN(n21170)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n6997), .CK(CLK), .Q(n7692), .QN(n21171)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n6996), .CK(CLK), .Q(n7693), .QN(n21172)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n6995), .CK(CLK), .Q(n7694), .QN(n21173)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n6994), .CK(CLK), .Q(n7695), .QN(n21174)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n6993), .CK(CLK), .Q(n7696), .QN(n21175)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n6992), .CK(CLK), .Q(n7697), .QN(n21176)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n6991), .CK(CLK), .Q(n7698), .QN(n21177)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n6990), .CK(CLK), .Q(n7699), .QN(n21178)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n6989), .CK(CLK), .Q(n7700), .QN(n21179)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n6988), .CK(CLK), .Q(n7701), .QN(n21180)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n6987), .CK(CLK), .Q(n7702), .QN(n21181)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n6986), .CK(CLK), .Q(n7703), .QN(n21182)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n6985), .CK(CLK), .Q(n7704), .QN(n21183)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n6984), .CK(CLK), .Q(n7705), .QN(n21184)
         );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n6983), .CK(CLK), .Q(n7706), .QN(n21185)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n6982), .CK(CLK), .Q(n7707), .QN(n21186)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n6980), .CK(CLK), .Q(n7709), .QN(n21187)
         );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5379), .CK(CLK), .Q(n7966), .QN(n20527)
         );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5378), .CK(CLK), .Q(n7967), .QN(n20528)
         );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5377), .CK(CLK), .Q(n7968), .QN(n20529)
         );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5376), .CK(CLK), .Q(n7969), .QN(n20530)
         );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5375), .CK(CLK), .Q(n7970), .QN(n20847)
         );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5374), .CK(CLK), .Q(n7971), .QN(n20848)
         );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5373), .CK(CLK), .Q(n7972), .QN(n20849)
         );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5372), .CK(CLK), .Q(n7973), .QN(n20850)
         );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5371), .CK(CLK), .Q(n7974), .QN(n20851)
         );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5370), .CK(CLK), .Q(n7975), .QN(n20852)
         );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5369), .CK(CLK), .Q(n7976), .QN(n20853)
         );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5368), .CK(CLK), .Q(n7977), .QN(n20854)
         );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5367), .CK(CLK), .Q(n7978), .QN(n20855)
         );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5366), .CK(CLK), .Q(n7979), .QN(n20856)
         );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5365), .CK(CLK), .Q(n7980), .QN(n20857)
         );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5364), .CK(CLK), .Q(n7981), .QN(n20858)
         );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5363), .CK(CLK), .Q(n7982), .QN(n20859)
         );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5362), .CK(CLK), .Q(n7983), .QN(n20860)
         );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5361), .CK(CLK), .Q(n7984), .QN(n20861)
         );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5360), .CK(CLK), .Q(n7985), .QN(n20862)
         );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5359), .CK(CLK), .Q(n7986), .QN(n20863)
         );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5358), .CK(CLK), .Q(n7987), .QN(n20864)
         );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5357), .CK(CLK), .Q(n7988), .QN(n20865)
         );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5356), .CK(CLK), .Q(n7989), .QN(n20866)
         );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5355), .CK(CLK), .Q(n7990), .QN(n20867)
         );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5354), .CK(CLK), .Q(n7991), .QN(n20868)
         );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5353), .CK(CLK), .Q(n7992), .QN(n20869)
         );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5352), .CK(CLK), .Q(n7993), .QN(n20870)
         );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5351), .CK(CLK), .Q(n7994), .QN(n20871)
         );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5350), .CK(CLK), .Q(n7995), .QN(n20872)
         );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5349), .CK(CLK), .Q(n7996), .QN(n20873)
         );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5348), .CK(CLK), .Q(n7997), .QN(n20874)
         );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5347), .CK(CLK), .Q(n7998), .QN(n20875)
         );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5346), .CK(CLK), .Q(n7999), .QN(n20876)
         );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5345), .CK(CLK), .Q(n8000), .QN(n20877)
         );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5344), .CK(CLK), .Q(n8001), .QN(n20878)
         );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5343), .CK(CLK), .Q(n8002), .QN(n20879)
         );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5342), .CK(CLK), .Q(n8003), .QN(n20880)
         );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5341), .CK(CLK), .Q(n8004), .QN(n20881)
         );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5340), .CK(CLK), .Q(n8005), .QN(n20882)
         );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5339), .CK(CLK), .Q(n8006), .QN(n20883)
         );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5338), .CK(CLK), .Q(n8007), .QN(n20884)
         );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5337), .CK(CLK), .Q(n8008), .QN(n20885)
         );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5336), .CK(CLK), .Q(n8009), .QN(n20886)
         );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5335), .CK(CLK), .Q(n8010), .QN(n20887)
         );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5334), .CK(CLK), .Q(n8011), .QN(n20888)
         );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5333), .CK(CLK), .Q(n8012), .QN(n20889)
         );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5332), .CK(CLK), .Q(n8013), .QN(n20890)
         );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5331), .CK(CLK), .Q(n8014), .QN(n20891)
         );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5330), .CK(CLK), .Q(n8015), .QN(n20892)
         );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5329), .CK(CLK), .Q(n8016), .QN(n20893)
         );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5328), .CK(CLK), .Q(n8017), .QN(n20894)
         );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5327), .CK(CLK), .Q(n8018), .QN(n20895)
         );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5326), .CK(CLK), .Q(n8019), .QN(n20896)
         );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5325), .CK(CLK), .Q(n8020), .QN(n20897)
         );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5324), .CK(CLK), .Q(n8021), .QN(n20898)
         );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5323), .CK(CLK), .Q(n8022), .QN(n20899)
         );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5322), .CK(CLK), .Q(n8023), .QN(n20900)
         );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5321), .CK(CLK), .Q(n8024), .QN(n20901)
         );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5320), .CK(CLK), .Q(n8025), .QN(n20902)
         );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5319), .CK(CLK), .Q(n8026), .QN(n20903)
         );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5318), .CK(CLK), .Q(n8027), .QN(n20904)
         );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5317), .CK(CLK), .Q(n8028), .QN(n20905)
         );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5316), .CK(CLK), .Q(n8029), .QN(n20906)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n4995), .CK(CLK), .Q(OUT2[63]) );
  DFF_X1 \OUT2_reg[62]  ( .D(n4994), .CK(CLK), .Q(OUT2[62]) );
  DFF_X1 \OUT2_reg[61]  ( .D(n4993), .CK(CLK), .Q(OUT2[61]) );
  DFF_X1 \OUT2_reg[60]  ( .D(n4992), .CK(CLK), .Q(OUT2[60]) );
  DFF_X1 \OUT2_reg[59]  ( .D(n4991), .CK(CLK), .Q(OUT2[59]) );
  DFF_X1 \OUT2_reg[58]  ( .D(n4990), .CK(CLK), .Q(OUT2[58]) );
  DFF_X1 \OUT2_reg[57]  ( .D(n4989), .CK(CLK), .Q(OUT2[57]) );
  DFF_X1 \OUT2_reg[56]  ( .D(n4988), .CK(CLK), .Q(OUT2[56]) );
  DFF_X1 \OUT2_reg[55]  ( .D(n4987), .CK(CLK), .Q(OUT2[55]) );
  DFF_X1 \OUT2_reg[54]  ( .D(n4986), .CK(CLK), .Q(OUT2[54]) );
  DFF_X1 \OUT2_reg[53]  ( .D(n4985), .CK(CLK), .Q(OUT2[53]) );
  DFF_X1 \OUT2_reg[52]  ( .D(n4984), .CK(CLK), .Q(OUT2[52]) );
  DFF_X1 \OUT2_reg[51]  ( .D(n4983), .CK(CLK), .Q(OUT2[51]) );
  DFF_X1 \OUT2_reg[50]  ( .D(n4982), .CK(CLK), .Q(OUT2[50]) );
  DFF_X1 \OUT2_reg[49]  ( .D(n4981), .CK(CLK), .Q(OUT2[49]) );
  DFF_X1 \OUT2_reg[48]  ( .D(n4980), .CK(CLK), .Q(OUT2[48]) );
  DFF_X1 \OUT2_reg[47]  ( .D(n4979), .CK(CLK), .Q(OUT2[47]) );
  DFF_X1 \OUT2_reg[46]  ( .D(n4978), .CK(CLK), .Q(OUT2[46]) );
  DFF_X1 \OUT2_reg[45]  ( .D(n4977), .CK(CLK), .Q(OUT2[45]) );
  DFF_X1 \OUT2_reg[44]  ( .D(n4976), .CK(CLK), .Q(OUT2[44]) );
  DFF_X1 \OUT2_reg[43]  ( .D(n4975), .CK(CLK), .Q(OUT2[43]) );
  DFF_X1 \OUT2_reg[42]  ( .D(n4974), .CK(CLK), .Q(OUT2[42]) );
  DFF_X1 \OUT2_reg[41]  ( .D(n4973), .CK(CLK), .Q(OUT2[41]) );
  DFF_X1 \OUT2_reg[40]  ( .D(n4972), .CK(CLK), .Q(OUT2[40]) );
  NOR2_X1 U18625 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n22542) );
  INV_X1 U18626 ( .A(n24832), .ZN(n24818) );
  INV_X1 U18627 ( .A(n24832), .ZN(n24817) );
  INV_X1 U18628 ( .A(n25549), .ZN(n25535) );
  INV_X1 U18629 ( .A(n25549), .ZN(n25536) );
  INV_X1 U18630 ( .A(n24833), .ZN(n24819) );
  INV_X1 U18631 ( .A(n25343), .ZN(n25329) );
  INV_X1 U18632 ( .A(n25343), .ZN(n25328) );
  INV_X1 U18633 ( .A(n25274), .ZN(n25260) );
  INV_X1 U18634 ( .A(n25274), .ZN(n25261) );
  INV_X1 U18635 ( .A(n25189), .ZN(n25175) );
  INV_X1 U18636 ( .A(n25189), .ZN(n25176) );
  INV_X1 U18637 ( .A(n25104), .ZN(n25090) );
  INV_X1 U18638 ( .A(n25104), .ZN(n25091) );
  INV_X1 U18639 ( .A(n25053), .ZN(n25039) );
  INV_X1 U18640 ( .A(n25053), .ZN(n25040) );
  INV_X1 U18641 ( .A(n25036), .ZN(n25022) );
  INV_X1 U18642 ( .A(n25036), .ZN(n25023) );
  INV_X1 U18643 ( .A(n24866), .ZN(n24852) );
  INV_X1 U18644 ( .A(n24866), .ZN(n24853) );
  INV_X1 U18645 ( .A(n24934), .ZN(n24920) );
  INV_X1 U18646 ( .A(n24934), .ZN(n24921) );
  INV_X1 U18647 ( .A(n24968), .ZN(n24954) );
  INV_X1 U18648 ( .A(n24968), .ZN(n24955) );
  INV_X1 U18649 ( .A(n24985), .ZN(n24971) );
  INV_X1 U18650 ( .A(n24985), .ZN(n24972) );
  INV_X1 U18651 ( .A(n25121), .ZN(n25107) );
  INV_X1 U18652 ( .A(n25121), .ZN(n25108) );
  INV_X1 U18653 ( .A(n25138), .ZN(n25124) );
  INV_X1 U18654 ( .A(n25138), .ZN(n25125) );
  INV_X1 U18655 ( .A(n25172), .ZN(n25158) );
  INV_X1 U18656 ( .A(n25172), .ZN(n25159) );
  INV_X1 U18657 ( .A(n25002), .ZN(n24988) );
  INV_X1 U18658 ( .A(n25002), .ZN(n24989) );
  INV_X1 U18659 ( .A(n25240), .ZN(n25226) );
  INV_X1 U18660 ( .A(n25240), .ZN(n25227) );
  INV_X1 U18661 ( .A(n25223), .ZN(n25209) );
  INV_X1 U18662 ( .A(n25223), .ZN(n25210) );
  INV_X1 U18663 ( .A(n25155), .ZN(n25141) );
  INV_X1 U18664 ( .A(n25155), .ZN(n25142) );
  INV_X1 U18665 ( .A(n24900), .ZN(n24886) );
  INV_X1 U18666 ( .A(n24900), .ZN(n24887) );
  INV_X1 U18667 ( .A(n25257), .ZN(n25243) );
  INV_X1 U18668 ( .A(n25257), .ZN(n25244) );
  INV_X1 U18669 ( .A(n25087), .ZN(n25073) );
  INV_X1 U18670 ( .A(n25087), .ZN(n25074) );
  INV_X1 U18671 ( .A(n25019), .ZN(n25005) );
  INV_X1 U18672 ( .A(n25019), .ZN(n25006) );
  INV_X1 U18673 ( .A(n24917), .ZN(n24903) );
  INV_X1 U18674 ( .A(n24917), .ZN(n24904) );
  INV_X1 U18675 ( .A(n24849), .ZN(n24835) );
  INV_X1 U18676 ( .A(n24849), .ZN(n24836) );
  INV_X1 U18677 ( .A(n25070), .ZN(n25056) );
  INV_X1 U18678 ( .A(n25070), .ZN(n25057) );
  INV_X1 U18679 ( .A(n25325), .ZN(n25311) );
  INV_X1 U18680 ( .A(n25325), .ZN(n25312) );
  INV_X1 U18681 ( .A(n25206), .ZN(n25192) );
  INV_X1 U18682 ( .A(n25206), .ZN(n25193) );
  INV_X1 U18683 ( .A(n25308), .ZN(n25294) );
  INV_X1 U18684 ( .A(n25308), .ZN(n25295) );
  INV_X1 U18685 ( .A(n24883), .ZN(n24869) );
  INV_X1 U18686 ( .A(n24883), .ZN(n24870) );
  INV_X1 U18687 ( .A(n24951), .ZN(n24937) );
  INV_X1 U18688 ( .A(n24951), .ZN(n24938) );
  INV_X1 U18689 ( .A(n25291), .ZN(n25277) );
  INV_X1 U18690 ( .A(n25291), .ZN(n25278) );
  BUF_X1 U18691 ( .A(n24814), .Z(n24832) );
  BUF_X1 U18692 ( .A(n25550), .Z(n25549) );
  BUF_X1 U18693 ( .A(n24813), .Z(n24831) );
  BUF_X1 U18694 ( .A(n24813), .Z(n24830) );
  BUF_X1 U18695 ( .A(n24813), .Z(n24829) );
  BUF_X1 U18696 ( .A(n24812), .Z(n24828) );
  BUF_X1 U18697 ( .A(n24812), .Z(n24827) );
  BUF_X1 U18698 ( .A(n24812), .Z(n24826) );
  BUF_X1 U18699 ( .A(n24811), .Z(n24825) );
  BUF_X1 U18700 ( .A(n24811), .Z(n24824) );
  BUF_X1 U18701 ( .A(n24811), .Z(n24823) );
  BUF_X1 U18702 ( .A(n24810), .Z(n24822) );
  BUF_X1 U18703 ( .A(n24810), .Z(n24821) );
  BUF_X1 U18704 ( .A(n24810), .Z(n24820) );
  BUF_X1 U18705 ( .A(n25550), .Z(n25537) );
  BUF_X1 U18706 ( .A(n25550), .Z(n25538) );
  BUF_X1 U18707 ( .A(n25550), .Z(n25539) );
  BUF_X1 U18708 ( .A(n25550), .Z(n25540) );
  BUF_X1 U18709 ( .A(n25550), .Z(n25541) );
  BUF_X1 U18710 ( .A(n25550), .Z(n25542) );
  BUF_X1 U18711 ( .A(n25550), .Z(n25543) );
  BUF_X1 U18712 ( .A(n25537), .Z(n25544) );
  BUF_X1 U18713 ( .A(n25538), .Z(n25545) );
  BUF_X1 U18714 ( .A(n25539), .Z(n25546) );
  BUF_X1 U18715 ( .A(n25540), .Z(n25547) );
  BUF_X1 U18716 ( .A(n25541), .Z(n25548) );
  BUF_X1 U18717 ( .A(n24814), .Z(n24833) );
  BUF_X1 U18718 ( .A(n22602), .Z(n24442) );
  BUF_X1 U18719 ( .A(n22602), .Z(n24438) );
  BUF_X1 U18720 ( .A(n22602), .Z(n24439) );
  BUF_X1 U18721 ( .A(n22602), .Z(n24440) );
  BUF_X1 U18722 ( .A(n22602), .Z(n24441) );
  BUF_X1 U18723 ( .A(n22571), .Z(n24586) );
  BUF_X1 U18724 ( .A(n22571), .Z(n24582) );
  BUF_X1 U18725 ( .A(n22571), .Z(n24583) );
  BUF_X1 U18726 ( .A(n22571), .Z(n24584) );
  BUF_X1 U18727 ( .A(n22571), .Z(n24585) );
  BUF_X1 U18728 ( .A(n22577), .Z(n24556) );
  BUF_X1 U18729 ( .A(n22577), .Z(n24552) );
  BUF_X1 U18730 ( .A(n22577), .Z(n24553) );
  BUF_X1 U18731 ( .A(n22577), .Z(n24554) );
  BUF_X1 U18732 ( .A(n22577), .Z(n24555) );
  BUF_X1 U18733 ( .A(n22594), .Z(n24490) );
  BUF_X1 U18734 ( .A(n22594), .Z(n24486) );
  BUF_X1 U18735 ( .A(n22594), .Z(n24487) );
  BUF_X1 U18736 ( .A(n22594), .Z(n24488) );
  BUF_X1 U18737 ( .A(n22594), .Z(n24489) );
  BUF_X1 U18738 ( .A(n22574), .Z(n24568) );
  BUF_X1 U18739 ( .A(n22574), .Z(n24564) );
  BUF_X1 U18740 ( .A(n22574), .Z(n24565) );
  BUF_X1 U18741 ( .A(n22574), .Z(n24566) );
  BUF_X1 U18742 ( .A(n22574), .Z(n24567) );
  BUF_X1 U18743 ( .A(n25003), .Z(n25002) );
  BUF_X1 U18744 ( .A(n25241), .Z(n25240) );
  BUF_X1 U18745 ( .A(n25224), .Z(n25223) );
  BUF_X1 U18746 ( .A(n25156), .Z(n25155) );
  BUF_X1 U18747 ( .A(n24901), .Z(n24900) );
  BUF_X1 U18748 ( .A(n25258), .Z(n25257) );
  BUF_X1 U18749 ( .A(n25088), .Z(n25087) );
  BUF_X1 U18750 ( .A(n25020), .Z(n25019) );
  BUF_X1 U18751 ( .A(n24918), .Z(n24917) );
  BUF_X1 U18752 ( .A(n24850), .Z(n24849) );
  BUF_X1 U18753 ( .A(n25071), .Z(n25070) );
  BUF_X1 U18754 ( .A(n25326), .Z(n25325) );
  BUF_X1 U18755 ( .A(n25207), .Z(n25206) );
  BUF_X1 U18756 ( .A(n25309), .Z(n25308) );
  BUF_X1 U18757 ( .A(n25344), .Z(n25342) );
  BUF_X1 U18758 ( .A(n25275), .Z(n25274) );
  BUF_X1 U18759 ( .A(n25190), .Z(n25189) );
  BUF_X1 U18760 ( .A(n25105), .Z(n25104) );
  BUF_X1 U18761 ( .A(n25054), .Z(n25053) );
  BUF_X1 U18762 ( .A(n25037), .Z(n25036) );
  BUF_X1 U18763 ( .A(n24867), .Z(n24866) );
  BUF_X1 U18764 ( .A(n24884), .Z(n24883) );
  BUF_X1 U18765 ( .A(n24935), .Z(n24934) );
  BUF_X1 U18766 ( .A(n24952), .Z(n24951) );
  BUF_X1 U18767 ( .A(n24969), .Z(n24968) );
  BUF_X1 U18768 ( .A(n24986), .Z(n24985) );
  BUF_X1 U18769 ( .A(n25122), .Z(n25121) );
  BUF_X1 U18770 ( .A(n25139), .Z(n25138) );
  BUF_X1 U18771 ( .A(n25173), .Z(n25172) );
  BUF_X1 U18772 ( .A(n25292), .Z(n25291) );
  BUF_X1 U18773 ( .A(n25344), .Z(n25331) );
  BUF_X1 U18774 ( .A(n25344), .Z(n25332) );
  BUF_X1 U18775 ( .A(n25344), .Z(n25333) );
  BUF_X1 U18776 ( .A(n25344), .Z(n25334) );
  BUF_X1 U18777 ( .A(n25331), .Z(n25341) );
  BUF_X1 U18778 ( .A(n25344), .Z(n25330) );
  BUF_X1 U18779 ( .A(n25003), .Z(n24990) );
  BUF_X1 U18780 ( .A(n25003), .Z(n24991) );
  BUF_X1 U18781 ( .A(n25003), .Z(n24992) );
  BUF_X1 U18782 ( .A(n25003), .Z(n24993) );
  BUF_X1 U18783 ( .A(n25241), .Z(n25228) );
  BUF_X1 U18784 ( .A(n25241), .Z(n25229) );
  BUF_X1 U18785 ( .A(n25241), .Z(n25230) );
  BUF_X1 U18786 ( .A(n25241), .Z(n25231) );
  BUF_X1 U18787 ( .A(n25224), .Z(n25211) );
  BUF_X1 U18788 ( .A(n25224), .Z(n25212) );
  BUF_X1 U18789 ( .A(n25224), .Z(n25213) );
  BUF_X1 U18790 ( .A(n25224), .Z(n25214) );
  BUF_X1 U18791 ( .A(n25156), .Z(n25143) );
  BUF_X1 U18792 ( .A(n25156), .Z(n25144) );
  BUF_X1 U18793 ( .A(n25156), .Z(n25145) );
  BUF_X1 U18794 ( .A(n25156), .Z(n25146) );
  BUF_X1 U18795 ( .A(n25003), .Z(n24994) );
  BUF_X1 U18796 ( .A(n25003), .Z(n24995) );
  BUF_X1 U18797 ( .A(n25003), .Z(n24996) );
  BUF_X1 U18798 ( .A(n24990), .Z(n24997) );
  BUF_X1 U18799 ( .A(n24991), .Z(n24998) );
  BUF_X1 U18800 ( .A(n24992), .Z(n24999) );
  BUF_X1 U18801 ( .A(n24993), .Z(n25000) );
  BUF_X1 U18802 ( .A(n24994), .Z(n25001) );
  BUF_X1 U18803 ( .A(n25241), .Z(n25232) );
  BUF_X1 U18804 ( .A(n25241), .Z(n25233) );
  BUF_X1 U18805 ( .A(n25241), .Z(n25234) );
  BUF_X1 U18806 ( .A(n25228), .Z(n25235) );
  BUF_X1 U18807 ( .A(n25229), .Z(n25236) );
  BUF_X1 U18808 ( .A(n25230), .Z(n25237) );
  BUF_X1 U18809 ( .A(n25231), .Z(n25238) );
  BUF_X1 U18810 ( .A(n25232), .Z(n25239) );
  BUF_X1 U18811 ( .A(n25224), .Z(n25215) );
  BUF_X1 U18812 ( .A(n25224), .Z(n25216) );
  BUF_X1 U18813 ( .A(n25224), .Z(n25217) );
  BUF_X1 U18814 ( .A(n25211), .Z(n25218) );
  BUF_X1 U18815 ( .A(n25212), .Z(n25219) );
  BUF_X1 U18816 ( .A(n25213), .Z(n25220) );
  BUF_X1 U18817 ( .A(n25214), .Z(n25221) );
  BUF_X1 U18818 ( .A(n25215), .Z(n25222) );
  BUF_X1 U18819 ( .A(n25156), .Z(n25147) );
  BUF_X1 U18820 ( .A(n25156), .Z(n25148) );
  BUF_X1 U18821 ( .A(n25156), .Z(n25149) );
  BUF_X1 U18822 ( .A(n25143), .Z(n25150) );
  BUF_X1 U18823 ( .A(n25144), .Z(n25151) );
  BUF_X1 U18824 ( .A(n25145), .Z(n25152) );
  BUF_X1 U18825 ( .A(n25146), .Z(n25153) );
  BUF_X1 U18826 ( .A(n25147), .Z(n25154) );
  BUF_X1 U18827 ( .A(n24901), .Z(n24888) );
  BUF_X1 U18828 ( .A(n24901), .Z(n24889) );
  BUF_X1 U18829 ( .A(n24901), .Z(n24890) );
  BUF_X1 U18830 ( .A(n24901), .Z(n24891) );
  BUF_X1 U18831 ( .A(n24901), .Z(n24892) );
  BUF_X1 U18832 ( .A(n24901), .Z(n24893) );
  BUF_X1 U18833 ( .A(n24901), .Z(n24894) );
  BUF_X1 U18834 ( .A(n24888), .Z(n24895) );
  BUF_X1 U18835 ( .A(n24889), .Z(n24896) );
  BUF_X1 U18836 ( .A(n24890), .Z(n24897) );
  BUF_X1 U18837 ( .A(n24891), .Z(n24898) );
  BUF_X1 U18838 ( .A(n24892), .Z(n24899) );
  BUF_X1 U18839 ( .A(n25258), .Z(n25245) );
  BUF_X1 U18840 ( .A(n25258), .Z(n25246) );
  BUF_X1 U18841 ( .A(n25258), .Z(n25247) );
  BUF_X1 U18842 ( .A(n25258), .Z(n25248) );
  BUF_X1 U18843 ( .A(n25088), .Z(n25075) );
  BUF_X1 U18844 ( .A(n25088), .Z(n25076) );
  BUF_X1 U18845 ( .A(n25088), .Z(n25077) );
  BUF_X1 U18846 ( .A(n25088), .Z(n25078) );
  BUF_X1 U18847 ( .A(n25020), .Z(n25007) );
  BUF_X1 U18848 ( .A(n25020), .Z(n25008) );
  BUF_X1 U18849 ( .A(n25020), .Z(n25009) );
  BUF_X1 U18850 ( .A(n25020), .Z(n25010) );
  BUF_X1 U18851 ( .A(n24918), .Z(n24905) );
  BUF_X1 U18852 ( .A(n24918), .Z(n24906) );
  BUF_X1 U18853 ( .A(n24918), .Z(n24907) );
  BUF_X1 U18854 ( .A(n24918), .Z(n24908) );
  BUF_X1 U18855 ( .A(n24850), .Z(n24837) );
  BUF_X1 U18856 ( .A(n24850), .Z(n24838) );
  BUF_X1 U18857 ( .A(n24850), .Z(n24839) );
  BUF_X1 U18858 ( .A(n24850), .Z(n24840) );
  BUF_X1 U18859 ( .A(n25258), .Z(n25249) );
  BUF_X1 U18860 ( .A(n25258), .Z(n25250) );
  BUF_X1 U18861 ( .A(n25258), .Z(n25251) );
  BUF_X1 U18862 ( .A(n25245), .Z(n25252) );
  BUF_X1 U18863 ( .A(n25246), .Z(n25253) );
  BUF_X1 U18864 ( .A(n25247), .Z(n25254) );
  BUF_X1 U18865 ( .A(n25248), .Z(n25255) );
  BUF_X1 U18866 ( .A(n25249), .Z(n25256) );
  BUF_X1 U18867 ( .A(n25088), .Z(n25079) );
  BUF_X1 U18868 ( .A(n25088), .Z(n25080) );
  BUF_X1 U18869 ( .A(n25088), .Z(n25081) );
  BUF_X1 U18870 ( .A(n25075), .Z(n25082) );
  BUF_X1 U18871 ( .A(n25076), .Z(n25083) );
  BUF_X1 U18872 ( .A(n25077), .Z(n25084) );
  BUF_X1 U18873 ( .A(n25078), .Z(n25085) );
  BUF_X1 U18874 ( .A(n25079), .Z(n25086) );
  BUF_X1 U18875 ( .A(n25020), .Z(n25011) );
  BUF_X1 U18876 ( .A(n25020), .Z(n25012) );
  BUF_X1 U18877 ( .A(n25020), .Z(n25013) );
  BUF_X1 U18878 ( .A(n25007), .Z(n25014) );
  BUF_X1 U18879 ( .A(n25008), .Z(n25015) );
  BUF_X1 U18880 ( .A(n25009), .Z(n25016) );
  BUF_X1 U18881 ( .A(n25010), .Z(n25017) );
  BUF_X1 U18882 ( .A(n25011), .Z(n25018) );
  BUF_X1 U18883 ( .A(n24918), .Z(n24909) );
  BUF_X1 U18884 ( .A(n24918), .Z(n24910) );
  BUF_X1 U18885 ( .A(n24918), .Z(n24911) );
  BUF_X1 U18886 ( .A(n24905), .Z(n24912) );
  BUF_X1 U18887 ( .A(n24906), .Z(n24913) );
  BUF_X1 U18888 ( .A(n24907), .Z(n24914) );
  BUF_X1 U18889 ( .A(n24908), .Z(n24915) );
  BUF_X1 U18890 ( .A(n24909), .Z(n24916) );
  BUF_X1 U18891 ( .A(n24850), .Z(n24841) );
  BUF_X1 U18892 ( .A(n24850), .Z(n24842) );
  BUF_X1 U18893 ( .A(n24850), .Z(n24843) );
  BUF_X1 U18894 ( .A(n24837), .Z(n24844) );
  BUF_X1 U18895 ( .A(n24838), .Z(n24845) );
  BUF_X1 U18896 ( .A(n24839), .Z(n24846) );
  BUF_X1 U18897 ( .A(n24840), .Z(n24847) );
  BUF_X1 U18898 ( .A(n24841), .Z(n24848) );
  BUF_X1 U18899 ( .A(n25071), .Z(n25058) );
  BUF_X1 U18900 ( .A(n25071), .Z(n25059) );
  BUF_X1 U18901 ( .A(n25071), .Z(n25060) );
  BUF_X1 U18902 ( .A(n25071), .Z(n25061) );
  BUF_X1 U18903 ( .A(n25071), .Z(n25062) );
  BUF_X1 U18904 ( .A(n25071), .Z(n25063) );
  BUF_X1 U18905 ( .A(n25071), .Z(n25064) );
  BUF_X1 U18906 ( .A(n25058), .Z(n25065) );
  BUF_X1 U18907 ( .A(n25059), .Z(n25066) );
  BUF_X1 U18908 ( .A(n25060), .Z(n25067) );
  BUF_X1 U18909 ( .A(n25061), .Z(n25068) );
  BUF_X1 U18910 ( .A(n25062), .Z(n25069) );
  BUF_X1 U18911 ( .A(n25326), .Z(n25313) );
  BUF_X1 U18912 ( .A(n25326), .Z(n25314) );
  BUF_X1 U18913 ( .A(n25326), .Z(n25315) );
  BUF_X1 U18914 ( .A(n25326), .Z(n25316) );
  BUF_X1 U18915 ( .A(n25207), .Z(n25194) );
  BUF_X1 U18916 ( .A(n25207), .Z(n25195) );
  BUF_X1 U18917 ( .A(n25207), .Z(n25196) );
  BUF_X1 U18918 ( .A(n25207), .Z(n25197) );
  BUF_X1 U18919 ( .A(n25309), .Z(n25296) );
  BUF_X1 U18920 ( .A(n25309), .Z(n25297) );
  BUF_X1 U18921 ( .A(n25309), .Z(n25298) );
  BUF_X1 U18922 ( .A(n25309), .Z(n25299) );
  BUF_X1 U18923 ( .A(n25326), .Z(n25317) );
  BUF_X1 U18924 ( .A(n25326), .Z(n25318) );
  BUF_X1 U18925 ( .A(n25326), .Z(n25319) );
  BUF_X1 U18926 ( .A(n25313), .Z(n25320) );
  BUF_X1 U18927 ( .A(n25314), .Z(n25321) );
  BUF_X1 U18928 ( .A(n25315), .Z(n25322) );
  BUF_X1 U18929 ( .A(n25316), .Z(n25323) );
  BUF_X1 U18930 ( .A(n25317), .Z(n25324) );
  BUF_X1 U18931 ( .A(n25207), .Z(n25198) );
  BUF_X1 U18932 ( .A(n25207), .Z(n25199) );
  BUF_X1 U18933 ( .A(n25207), .Z(n25200) );
  BUF_X1 U18934 ( .A(n25194), .Z(n25201) );
  BUF_X1 U18935 ( .A(n25195), .Z(n25202) );
  BUF_X1 U18936 ( .A(n25196), .Z(n25203) );
  BUF_X1 U18937 ( .A(n25197), .Z(n25204) );
  BUF_X1 U18938 ( .A(n25198), .Z(n25205) );
  BUF_X1 U18939 ( .A(n25309), .Z(n25300) );
  BUF_X1 U18940 ( .A(n25309), .Z(n25301) );
  BUF_X1 U18941 ( .A(n25309), .Z(n25302) );
  BUF_X1 U18942 ( .A(n25296), .Z(n25303) );
  BUF_X1 U18943 ( .A(n25297), .Z(n25304) );
  BUF_X1 U18944 ( .A(n25298), .Z(n25305) );
  BUF_X1 U18945 ( .A(n25299), .Z(n25306) );
  BUF_X1 U18946 ( .A(n25300), .Z(n25307) );
  BUF_X1 U18947 ( .A(n24884), .Z(n24877) );
  BUF_X1 U18948 ( .A(n24877), .Z(n24878) );
  BUF_X1 U18949 ( .A(n24871), .Z(n24879) );
  BUF_X1 U18950 ( .A(n24872), .Z(n24880) );
  BUF_X1 U18951 ( .A(n24873), .Z(n24881) );
  BUF_X1 U18952 ( .A(n24874), .Z(n24882) );
  BUF_X1 U18953 ( .A(n25344), .Z(n25335) );
  BUF_X1 U18954 ( .A(n25344), .Z(n25336) );
  BUF_X1 U18955 ( .A(n25332), .Z(n25337) );
  BUF_X1 U18956 ( .A(n25333), .Z(n25338) );
  BUF_X1 U18957 ( .A(n25334), .Z(n25339) );
  BUF_X1 U18958 ( .A(n25330), .Z(n25340) );
  BUF_X1 U18959 ( .A(n25275), .Z(n25262) );
  BUF_X1 U18960 ( .A(n25275), .Z(n25263) );
  BUF_X1 U18961 ( .A(n25275), .Z(n25264) );
  BUF_X1 U18962 ( .A(n25275), .Z(n25265) );
  BUF_X1 U18963 ( .A(n25190), .Z(n25177) );
  BUF_X1 U18964 ( .A(n25190), .Z(n25178) );
  BUF_X1 U18965 ( .A(n25190), .Z(n25179) );
  BUF_X1 U18966 ( .A(n25190), .Z(n25180) );
  BUF_X1 U18967 ( .A(n25105), .Z(n25092) );
  BUF_X1 U18968 ( .A(n25105), .Z(n25093) );
  BUF_X1 U18969 ( .A(n25105), .Z(n25094) );
  BUF_X1 U18970 ( .A(n25105), .Z(n25095) );
  BUF_X1 U18971 ( .A(n25054), .Z(n25041) );
  BUF_X1 U18972 ( .A(n25054), .Z(n25042) );
  BUF_X1 U18973 ( .A(n25054), .Z(n25043) );
  BUF_X1 U18974 ( .A(n25054), .Z(n25044) );
  BUF_X1 U18975 ( .A(n25037), .Z(n25024) );
  BUF_X1 U18976 ( .A(n25037), .Z(n25025) );
  BUF_X1 U18977 ( .A(n25037), .Z(n25026) );
  BUF_X1 U18978 ( .A(n25037), .Z(n25027) );
  BUF_X1 U18979 ( .A(n25275), .Z(n25266) );
  BUF_X1 U18980 ( .A(n25275), .Z(n25267) );
  BUF_X1 U18981 ( .A(n25275), .Z(n25268) );
  BUF_X1 U18982 ( .A(n25262), .Z(n25269) );
  BUF_X1 U18983 ( .A(n25263), .Z(n25270) );
  BUF_X1 U18984 ( .A(n25264), .Z(n25271) );
  BUF_X1 U18985 ( .A(n25265), .Z(n25272) );
  BUF_X1 U18986 ( .A(n25266), .Z(n25273) );
  BUF_X1 U18987 ( .A(n25190), .Z(n25181) );
  BUF_X1 U18988 ( .A(n25190), .Z(n25182) );
  BUF_X1 U18989 ( .A(n25190), .Z(n25183) );
  BUF_X1 U18990 ( .A(n25177), .Z(n25184) );
  BUF_X1 U18991 ( .A(n25178), .Z(n25185) );
  BUF_X1 U18992 ( .A(n25179), .Z(n25186) );
  BUF_X1 U18993 ( .A(n25180), .Z(n25187) );
  BUF_X1 U18994 ( .A(n25181), .Z(n25188) );
  BUF_X1 U18995 ( .A(n25105), .Z(n25096) );
  BUF_X1 U18996 ( .A(n25105), .Z(n25097) );
  BUF_X1 U18997 ( .A(n25105), .Z(n25098) );
  BUF_X1 U18998 ( .A(n25092), .Z(n25099) );
  BUF_X1 U18999 ( .A(n25093), .Z(n25100) );
  BUF_X1 U19000 ( .A(n25094), .Z(n25101) );
  BUF_X1 U19001 ( .A(n25095), .Z(n25102) );
  BUF_X1 U19002 ( .A(n25096), .Z(n25103) );
  BUF_X1 U19003 ( .A(n25054), .Z(n25045) );
  BUF_X1 U19004 ( .A(n25054), .Z(n25046) );
  BUF_X1 U19005 ( .A(n25054), .Z(n25047) );
  BUF_X1 U19006 ( .A(n25041), .Z(n25048) );
  BUF_X1 U19007 ( .A(n25042), .Z(n25049) );
  BUF_X1 U19008 ( .A(n25043), .Z(n25050) );
  BUF_X1 U19009 ( .A(n25044), .Z(n25051) );
  BUF_X1 U19010 ( .A(n25045), .Z(n25052) );
  BUF_X1 U19011 ( .A(n25037), .Z(n25028) );
  BUF_X1 U19012 ( .A(n25037), .Z(n25029) );
  BUF_X1 U19013 ( .A(n25037), .Z(n25030) );
  BUF_X1 U19014 ( .A(n25024), .Z(n25031) );
  BUF_X1 U19015 ( .A(n25025), .Z(n25032) );
  BUF_X1 U19016 ( .A(n25026), .Z(n25033) );
  BUF_X1 U19017 ( .A(n25027), .Z(n25034) );
  BUF_X1 U19018 ( .A(n25028), .Z(n25035) );
  BUF_X1 U19019 ( .A(n24867), .Z(n24854) );
  BUF_X1 U19020 ( .A(n24867), .Z(n24855) );
  BUF_X1 U19021 ( .A(n24867), .Z(n24856) );
  BUF_X1 U19022 ( .A(n24867), .Z(n24857) );
  BUF_X1 U19023 ( .A(n24867), .Z(n24858) );
  BUF_X1 U19024 ( .A(n24867), .Z(n24859) );
  BUF_X1 U19025 ( .A(n24867), .Z(n24860) );
  BUF_X1 U19026 ( .A(n24854), .Z(n24861) );
  BUF_X1 U19027 ( .A(n24855), .Z(n24862) );
  BUF_X1 U19028 ( .A(n24856), .Z(n24863) );
  BUF_X1 U19029 ( .A(n24857), .Z(n24864) );
  BUF_X1 U19030 ( .A(n24858), .Z(n24865) );
  BUF_X1 U19031 ( .A(n24884), .Z(n24871) );
  BUF_X1 U19032 ( .A(n24884), .Z(n24872) );
  BUF_X1 U19033 ( .A(n24884), .Z(n24873) );
  BUF_X1 U19034 ( .A(n24884), .Z(n24874) );
  BUF_X1 U19035 ( .A(n24884), .Z(n24875) );
  BUF_X1 U19036 ( .A(n24884), .Z(n24876) );
  BUF_X1 U19037 ( .A(n24935), .Z(n24922) );
  BUF_X1 U19038 ( .A(n24935), .Z(n24923) );
  BUF_X1 U19039 ( .A(n24935), .Z(n24924) );
  BUF_X1 U19040 ( .A(n24935), .Z(n24925) );
  BUF_X1 U19041 ( .A(n24935), .Z(n24926) );
  BUF_X1 U19042 ( .A(n24935), .Z(n24927) );
  BUF_X1 U19043 ( .A(n24935), .Z(n24928) );
  BUF_X1 U19044 ( .A(n24922), .Z(n24929) );
  BUF_X1 U19045 ( .A(n24923), .Z(n24930) );
  BUF_X1 U19046 ( .A(n24924), .Z(n24931) );
  BUF_X1 U19047 ( .A(n24925), .Z(n24932) );
  BUF_X1 U19048 ( .A(n24926), .Z(n24933) );
  BUF_X1 U19049 ( .A(n24952), .Z(n24939) );
  BUF_X1 U19050 ( .A(n24952), .Z(n24940) );
  BUF_X1 U19051 ( .A(n24952), .Z(n24941) );
  BUF_X1 U19052 ( .A(n24952), .Z(n24942) );
  BUF_X1 U19053 ( .A(n24952), .Z(n24943) );
  BUF_X1 U19054 ( .A(n24952), .Z(n24944) );
  BUF_X1 U19055 ( .A(n24952), .Z(n24945) );
  BUF_X1 U19056 ( .A(n24939), .Z(n24946) );
  BUF_X1 U19057 ( .A(n24940), .Z(n24947) );
  BUF_X1 U19058 ( .A(n24941), .Z(n24948) );
  BUF_X1 U19059 ( .A(n24942), .Z(n24949) );
  BUF_X1 U19060 ( .A(n24943), .Z(n24950) );
  BUF_X1 U19061 ( .A(n24969), .Z(n24956) );
  BUF_X1 U19062 ( .A(n24969), .Z(n24957) );
  BUF_X1 U19063 ( .A(n24969), .Z(n24958) );
  BUF_X1 U19064 ( .A(n24969), .Z(n24959) );
  BUF_X1 U19065 ( .A(n24969), .Z(n24960) );
  BUF_X1 U19066 ( .A(n24969), .Z(n24961) );
  BUF_X1 U19067 ( .A(n24969), .Z(n24962) );
  BUF_X1 U19068 ( .A(n24956), .Z(n24963) );
  BUF_X1 U19069 ( .A(n24957), .Z(n24964) );
  BUF_X1 U19070 ( .A(n24958), .Z(n24965) );
  BUF_X1 U19071 ( .A(n24959), .Z(n24966) );
  BUF_X1 U19072 ( .A(n24960), .Z(n24967) );
  BUF_X1 U19073 ( .A(n24986), .Z(n24973) );
  BUF_X1 U19074 ( .A(n24986), .Z(n24974) );
  BUF_X1 U19075 ( .A(n24986), .Z(n24975) );
  BUF_X1 U19076 ( .A(n24986), .Z(n24976) );
  BUF_X1 U19077 ( .A(n24986), .Z(n24977) );
  BUF_X1 U19078 ( .A(n24986), .Z(n24978) );
  BUF_X1 U19079 ( .A(n24986), .Z(n24979) );
  BUF_X1 U19080 ( .A(n24973), .Z(n24980) );
  BUF_X1 U19081 ( .A(n24974), .Z(n24981) );
  BUF_X1 U19082 ( .A(n24975), .Z(n24982) );
  BUF_X1 U19083 ( .A(n24976), .Z(n24983) );
  BUF_X1 U19084 ( .A(n24977), .Z(n24984) );
  BUF_X1 U19085 ( .A(n25122), .Z(n25109) );
  BUF_X1 U19086 ( .A(n25122), .Z(n25110) );
  BUF_X1 U19087 ( .A(n25122), .Z(n25111) );
  BUF_X1 U19088 ( .A(n25122), .Z(n25112) );
  BUF_X1 U19089 ( .A(n25122), .Z(n25113) );
  BUF_X1 U19090 ( .A(n25122), .Z(n25114) );
  BUF_X1 U19091 ( .A(n25122), .Z(n25115) );
  BUF_X1 U19092 ( .A(n25109), .Z(n25116) );
  BUF_X1 U19093 ( .A(n25110), .Z(n25117) );
  BUF_X1 U19094 ( .A(n25111), .Z(n25118) );
  BUF_X1 U19095 ( .A(n25112), .Z(n25119) );
  BUF_X1 U19096 ( .A(n25113), .Z(n25120) );
  BUF_X1 U19097 ( .A(n25139), .Z(n25126) );
  BUF_X1 U19098 ( .A(n25139), .Z(n25127) );
  BUF_X1 U19099 ( .A(n25139), .Z(n25128) );
  BUF_X1 U19100 ( .A(n25139), .Z(n25129) );
  BUF_X1 U19101 ( .A(n25139), .Z(n25130) );
  BUF_X1 U19102 ( .A(n25139), .Z(n25131) );
  BUF_X1 U19103 ( .A(n25139), .Z(n25132) );
  BUF_X1 U19104 ( .A(n25126), .Z(n25133) );
  BUF_X1 U19105 ( .A(n25127), .Z(n25134) );
  BUF_X1 U19106 ( .A(n25128), .Z(n25135) );
  BUF_X1 U19107 ( .A(n25129), .Z(n25136) );
  BUF_X1 U19108 ( .A(n25130), .Z(n25137) );
  BUF_X1 U19109 ( .A(n25173), .Z(n25160) );
  BUF_X1 U19110 ( .A(n25173), .Z(n25161) );
  BUF_X1 U19111 ( .A(n25173), .Z(n25162) );
  BUF_X1 U19112 ( .A(n25173), .Z(n25163) );
  BUF_X1 U19113 ( .A(n25173), .Z(n25164) );
  BUF_X1 U19114 ( .A(n25173), .Z(n25165) );
  BUF_X1 U19115 ( .A(n25173), .Z(n25166) );
  BUF_X1 U19116 ( .A(n25160), .Z(n25167) );
  BUF_X1 U19117 ( .A(n25161), .Z(n25168) );
  BUF_X1 U19118 ( .A(n25162), .Z(n25169) );
  BUF_X1 U19119 ( .A(n25163), .Z(n25170) );
  BUF_X1 U19120 ( .A(n25164), .Z(n25171) );
  BUF_X1 U19121 ( .A(n25292), .Z(n25279) );
  BUF_X1 U19122 ( .A(n25292), .Z(n25280) );
  BUF_X1 U19123 ( .A(n25292), .Z(n25281) );
  BUF_X1 U19124 ( .A(n25292), .Z(n25282) );
  BUF_X1 U19125 ( .A(n25292), .Z(n25283) );
  BUF_X1 U19126 ( .A(n25292), .Z(n25284) );
  BUF_X1 U19127 ( .A(n25292), .Z(n25285) );
  BUF_X1 U19128 ( .A(n25279), .Z(n25286) );
  BUF_X1 U19129 ( .A(n25280), .Z(n25287) );
  BUF_X1 U19130 ( .A(n25281), .Z(n25288) );
  BUF_X1 U19131 ( .A(n25282), .Z(n25289) );
  BUF_X1 U19132 ( .A(n25283), .Z(n25290) );
  BUF_X1 U19133 ( .A(n25335), .Z(n25343) );
  BUF_X1 U19134 ( .A(n24815), .Z(n24813) );
  BUF_X1 U19135 ( .A(n24815), .Z(n24812) );
  BUF_X1 U19136 ( .A(n24816), .Z(n24811) );
  BUF_X1 U19137 ( .A(n24816), .Z(n24810) );
  BUF_X1 U19138 ( .A(n24815), .Z(n24814) );
  INV_X1 U19139 ( .A(n25534), .ZN(n25550) );
  BUF_X1 U19140 ( .A(n22598), .Z(n24466) );
  BUF_X1 U19141 ( .A(n22598), .Z(n24462) );
  BUF_X1 U19142 ( .A(n22598), .Z(n24463) );
  BUF_X1 U19143 ( .A(n22598), .Z(n24464) );
  BUF_X1 U19144 ( .A(n22598), .Z(n24465) );
  BUF_X1 U19145 ( .A(n21307), .Z(n24786) );
  BUF_X1 U19146 ( .A(n21312), .Z(n24762) );
  BUF_X1 U19147 ( .A(n21317), .Z(n24738) );
  BUF_X1 U19148 ( .A(n21322), .Z(n24714) );
  BUF_X1 U19149 ( .A(n21331), .Z(n24690) );
  BUF_X1 U19150 ( .A(n21336), .Z(n24666) );
  BUF_X1 U19151 ( .A(n21341), .Z(n24642) );
  BUF_X1 U19152 ( .A(n21346), .Z(n24618) );
  BUF_X1 U19153 ( .A(n21307), .Z(n24787) );
  BUF_X1 U19154 ( .A(n21312), .Z(n24763) );
  BUF_X1 U19155 ( .A(n21317), .Z(n24739) );
  BUF_X1 U19156 ( .A(n21322), .Z(n24715) );
  BUF_X1 U19157 ( .A(n21331), .Z(n24691) );
  BUF_X1 U19158 ( .A(n21336), .Z(n24667) );
  BUF_X1 U19159 ( .A(n21341), .Z(n24643) );
  BUF_X1 U19160 ( .A(n21346), .Z(n24619) );
  BUF_X1 U19161 ( .A(n21307), .Z(n24788) );
  BUF_X1 U19162 ( .A(n21312), .Z(n24764) );
  BUF_X1 U19163 ( .A(n21317), .Z(n24740) );
  BUF_X1 U19164 ( .A(n21322), .Z(n24716) );
  BUF_X1 U19165 ( .A(n21331), .Z(n24692) );
  BUF_X1 U19166 ( .A(n21336), .Z(n24668) );
  BUF_X1 U19167 ( .A(n21341), .Z(n24644) );
  BUF_X1 U19168 ( .A(n21346), .Z(n24620) );
  BUF_X1 U19169 ( .A(n21307), .Z(n24789) );
  BUF_X1 U19170 ( .A(n21312), .Z(n24765) );
  BUF_X1 U19171 ( .A(n21317), .Z(n24741) );
  BUF_X1 U19172 ( .A(n21322), .Z(n24717) );
  BUF_X1 U19173 ( .A(n21331), .Z(n24693) );
  BUF_X1 U19174 ( .A(n21336), .Z(n24669) );
  BUF_X1 U19175 ( .A(n21341), .Z(n24645) );
  BUF_X1 U19176 ( .A(n21346), .Z(n24621) );
  BUF_X1 U19177 ( .A(n21307), .Z(n24790) );
  BUF_X1 U19178 ( .A(n21312), .Z(n24766) );
  BUF_X1 U19179 ( .A(n21317), .Z(n24742) );
  BUF_X1 U19180 ( .A(n21322), .Z(n24718) );
  BUF_X1 U19181 ( .A(n21331), .Z(n24694) );
  BUF_X1 U19182 ( .A(n21336), .Z(n24670) );
  BUF_X1 U19183 ( .A(n21341), .Z(n24646) );
  BUF_X1 U19184 ( .A(n21346), .Z(n24622) );
  BUF_X1 U19185 ( .A(n22607), .Z(n24418) );
  BUF_X1 U19186 ( .A(n22607), .Z(n24414) );
  BUF_X1 U19187 ( .A(n22607), .Z(n24415) );
  BUF_X1 U19188 ( .A(n22607), .Z(n24416) );
  BUF_X1 U19189 ( .A(n22607), .Z(n24417) );
  BUF_X1 U19190 ( .A(n21302), .Z(n24792) );
  BUF_X1 U19191 ( .A(n21302), .Z(n24793) );
  BUF_X1 U19192 ( .A(n21302), .Z(n24794) );
  BUF_X1 U19193 ( .A(n21302), .Z(n24795) );
  BUF_X1 U19194 ( .A(n21302), .Z(n24796) );
  BUF_X1 U19195 ( .A(n22586), .Z(n24514) );
  BUF_X1 U19196 ( .A(n22586), .Z(n24510) );
  BUF_X1 U19197 ( .A(n22586), .Z(n24511) );
  BUF_X1 U19198 ( .A(n22586), .Z(n24512) );
  BUF_X1 U19199 ( .A(n22586), .Z(n24513) );
  BUF_X1 U19200 ( .A(n22576), .Z(n24562) );
  BUF_X1 U19201 ( .A(n22581), .Z(n24538) );
  BUF_X1 U19202 ( .A(n22576), .Z(n24558) );
  BUF_X1 U19203 ( .A(n22581), .Z(n24534) );
  BUF_X1 U19204 ( .A(n22576), .Z(n24559) );
  BUF_X1 U19205 ( .A(n22581), .Z(n24535) );
  BUF_X1 U19206 ( .A(n22576), .Z(n24560) );
  BUF_X1 U19207 ( .A(n22581), .Z(n24536) );
  BUF_X1 U19208 ( .A(n22576), .Z(n24561) );
  BUF_X1 U19209 ( .A(n22581), .Z(n24537) );
  BUF_X1 U19210 ( .A(n21308), .Z(n24780) );
  BUF_X1 U19211 ( .A(n21313), .Z(n24756) );
  BUF_X1 U19212 ( .A(n21318), .Z(n24732) );
  BUF_X1 U19213 ( .A(n21323), .Z(n24708) );
  BUF_X1 U19214 ( .A(n21332), .Z(n24684) );
  BUF_X1 U19215 ( .A(n21337), .Z(n24660) );
  BUF_X1 U19216 ( .A(n21342), .Z(n24636) );
  BUF_X1 U19217 ( .A(n21347), .Z(n24612) );
  BUF_X1 U19218 ( .A(n21308), .Z(n24781) );
  BUF_X1 U19219 ( .A(n21313), .Z(n24757) );
  BUF_X1 U19220 ( .A(n21318), .Z(n24733) );
  BUF_X1 U19221 ( .A(n21323), .Z(n24709) );
  BUF_X1 U19222 ( .A(n21332), .Z(n24685) );
  BUF_X1 U19223 ( .A(n21337), .Z(n24661) );
  BUF_X1 U19224 ( .A(n21342), .Z(n24637) );
  BUF_X1 U19225 ( .A(n21347), .Z(n24613) );
  BUF_X1 U19226 ( .A(n21308), .Z(n24782) );
  BUF_X1 U19227 ( .A(n21313), .Z(n24758) );
  BUF_X1 U19228 ( .A(n21318), .Z(n24734) );
  BUF_X1 U19229 ( .A(n21323), .Z(n24710) );
  BUF_X1 U19230 ( .A(n21332), .Z(n24686) );
  BUF_X1 U19231 ( .A(n21337), .Z(n24662) );
  BUF_X1 U19232 ( .A(n21342), .Z(n24638) );
  BUF_X1 U19233 ( .A(n21347), .Z(n24614) );
  BUF_X1 U19234 ( .A(n21308), .Z(n24783) );
  BUF_X1 U19235 ( .A(n21313), .Z(n24759) );
  BUF_X1 U19236 ( .A(n21318), .Z(n24735) );
  BUF_X1 U19237 ( .A(n21323), .Z(n24711) );
  BUF_X1 U19238 ( .A(n21332), .Z(n24687) );
  BUF_X1 U19239 ( .A(n21337), .Z(n24663) );
  BUF_X1 U19240 ( .A(n21342), .Z(n24639) );
  BUF_X1 U19241 ( .A(n21347), .Z(n24615) );
  BUF_X1 U19242 ( .A(n21308), .Z(n24784) );
  BUF_X1 U19243 ( .A(n21313), .Z(n24760) );
  BUF_X1 U19244 ( .A(n21318), .Z(n24736) );
  BUF_X1 U19245 ( .A(n21323), .Z(n24712) );
  BUF_X1 U19246 ( .A(n21332), .Z(n24688) );
  BUF_X1 U19247 ( .A(n21337), .Z(n24664) );
  BUF_X1 U19248 ( .A(n21342), .Z(n24640) );
  BUF_X1 U19249 ( .A(n21347), .Z(n24616) );
  BUF_X1 U19250 ( .A(n22603), .Z(n24436) );
  BUF_X1 U19251 ( .A(n22603), .Z(n24432) );
  BUF_X1 U19252 ( .A(n22603), .Z(n24433) );
  BUF_X1 U19253 ( .A(n22603), .Z(n24434) );
  BUF_X1 U19254 ( .A(n22603), .Z(n24435) );
  BUF_X1 U19255 ( .A(n22568), .Z(n24598) );
  BUF_X1 U19256 ( .A(n22583), .Z(n24526) );
  BUF_X1 U19257 ( .A(n22573), .Z(n24574) );
  BUF_X1 U19258 ( .A(n22578), .Z(n24550) );
  BUF_X1 U19259 ( .A(n22568), .Z(n24595) );
  BUF_X1 U19260 ( .A(n22583), .Z(n24523) );
  BUF_X1 U19261 ( .A(n22573), .Z(n24571) );
  BUF_X1 U19262 ( .A(n22578), .Z(n24547) );
  BUF_X1 U19263 ( .A(n22568), .Z(n24596) );
  BUF_X1 U19264 ( .A(n22583), .Z(n24524) );
  BUF_X1 U19265 ( .A(n22573), .Z(n24572) );
  BUF_X1 U19266 ( .A(n22578), .Z(n24548) );
  BUF_X1 U19267 ( .A(n22568), .Z(n24597) );
  BUF_X1 U19268 ( .A(n22583), .Z(n24525) );
  BUF_X1 U19269 ( .A(n22573), .Z(n24573) );
  BUF_X1 U19270 ( .A(n22578), .Z(n24549) );
  BUF_X1 U19271 ( .A(n22601), .Z(n24448) );
  BUF_X1 U19272 ( .A(n22601), .Z(n24444) );
  BUF_X1 U19273 ( .A(n22601), .Z(n24445) );
  BUF_X1 U19274 ( .A(n22601), .Z(n24446) );
  BUF_X1 U19275 ( .A(n22601), .Z(n24447) );
  BUF_X1 U19276 ( .A(n22587), .Z(n24508) );
  BUF_X1 U19277 ( .A(n22587), .Z(n24504) );
  BUF_X1 U19278 ( .A(n22587), .Z(n24505) );
  BUF_X1 U19279 ( .A(n22587), .Z(n24506) );
  BUF_X1 U19280 ( .A(n22587), .Z(n24507) );
  BUF_X1 U19281 ( .A(n22599), .Z(n24460) );
  BUF_X1 U19282 ( .A(n22599), .Z(n24456) );
  BUF_X1 U19283 ( .A(n22599), .Z(n24457) );
  BUF_X1 U19284 ( .A(n22599), .Z(n24458) );
  BUF_X1 U19285 ( .A(n22599), .Z(n24459) );
  BUF_X1 U19286 ( .A(n22600), .Z(n24454) );
  BUF_X1 U19287 ( .A(n22600), .Z(n24450) );
  BUF_X1 U19288 ( .A(n22600), .Z(n24451) );
  BUF_X1 U19289 ( .A(n22600), .Z(n24452) );
  BUF_X1 U19290 ( .A(n22600), .Z(n24453) );
  BUF_X1 U19291 ( .A(n22572), .Z(n24580) );
  BUF_X1 U19292 ( .A(n22582), .Z(n24532) );
  BUF_X1 U19293 ( .A(n22572), .Z(n24576) );
  BUF_X1 U19294 ( .A(n22582), .Z(n24528) );
  BUF_X1 U19295 ( .A(n22572), .Z(n24577) );
  BUF_X1 U19296 ( .A(n22582), .Z(n24529) );
  BUF_X1 U19297 ( .A(n22572), .Z(n24578) );
  BUF_X1 U19298 ( .A(n22582), .Z(n24530) );
  BUF_X1 U19299 ( .A(n22572), .Z(n24579) );
  BUF_X1 U19300 ( .A(n22582), .Z(n24531) );
  BUF_X1 U19301 ( .A(n22588), .Z(n24502) );
  BUF_X1 U19302 ( .A(n22588), .Z(n24498) );
  BUF_X1 U19303 ( .A(n22588), .Z(n24499) );
  BUF_X1 U19304 ( .A(n22588), .Z(n24500) );
  BUF_X1 U19305 ( .A(n22588), .Z(n24501) );
  BUF_X1 U19306 ( .A(n25555), .Z(n25562) );
  BUF_X1 U19307 ( .A(n25556), .Z(n25563) );
  BUF_X1 U19308 ( .A(n25555), .Z(n25561) );
  BUF_X1 U19309 ( .A(n25555), .Z(n25560) );
  BUF_X1 U19310 ( .A(n25554), .Z(n25559) );
  BUF_X1 U19311 ( .A(n25554), .Z(n25558) );
  BUF_X1 U19312 ( .A(n25554), .Z(n25557) );
  BUF_X1 U19313 ( .A(n21310), .Z(n24774) );
  BUF_X1 U19314 ( .A(n21315), .Z(n24750) );
  BUF_X1 U19315 ( .A(n21320), .Z(n24726) );
  BUF_X1 U19316 ( .A(n21325), .Z(n24702) );
  BUF_X1 U19317 ( .A(n21334), .Z(n24678) );
  BUF_X1 U19318 ( .A(n21339), .Z(n24654) );
  BUF_X1 U19319 ( .A(n21344), .Z(n24630) );
  BUF_X1 U19320 ( .A(n21349), .Z(n24606) );
  BUF_X1 U19321 ( .A(n21310), .Z(n24775) );
  BUF_X1 U19322 ( .A(n21315), .Z(n24751) );
  BUF_X1 U19323 ( .A(n21320), .Z(n24727) );
  BUF_X1 U19324 ( .A(n21325), .Z(n24703) );
  BUF_X1 U19325 ( .A(n21334), .Z(n24679) );
  BUF_X1 U19326 ( .A(n21339), .Z(n24655) );
  BUF_X1 U19327 ( .A(n21344), .Z(n24631) );
  BUF_X1 U19328 ( .A(n21349), .Z(n24607) );
  BUF_X1 U19329 ( .A(n21310), .Z(n24776) );
  BUF_X1 U19330 ( .A(n21315), .Z(n24752) );
  BUF_X1 U19331 ( .A(n21320), .Z(n24728) );
  BUF_X1 U19332 ( .A(n21325), .Z(n24704) );
  BUF_X1 U19333 ( .A(n21334), .Z(n24680) );
  BUF_X1 U19334 ( .A(n21339), .Z(n24656) );
  BUF_X1 U19335 ( .A(n21344), .Z(n24632) );
  BUF_X1 U19336 ( .A(n21349), .Z(n24608) );
  BUF_X1 U19337 ( .A(n21310), .Z(n24777) );
  BUF_X1 U19338 ( .A(n21315), .Z(n24753) );
  BUF_X1 U19339 ( .A(n21320), .Z(n24729) );
  BUF_X1 U19340 ( .A(n21325), .Z(n24705) );
  BUF_X1 U19341 ( .A(n21334), .Z(n24681) );
  BUF_X1 U19342 ( .A(n21339), .Z(n24657) );
  BUF_X1 U19343 ( .A(n21344), .Z(n24633) );
  BUF_X1 U19344 ( .A(n21349), .Z(n24609) );
  BUF_X1 U19345 ( .A(n21310), .Z(n24778) );
  BUF_X1 U19346 ( .A(n21315), .Z(n24754) );
  BUF_X1 U19347 ( .A(n21320), .Z(n24730) );
  BUF_X1 U19348 ( .A(n21325), .Z(n24706) );
  BUF_X1 U19349 ( .A(n21334), .Z(n24682) );
  BUF_X1 U19350 ( .A(n21339), .Z(n24658) );
  BUF_X1 U19351 ( .A(n21344), .Z(n24634) );
  BUF_X1 U19352 ( .A(n21349), .Z(n24610) );
  BUF_X1 U19353 ( .A(n22593), .Z(n24496) );
  BUF_X1 U19354 ( .A(n22595), .Z(n24484) );
  BUF_X1 U19355 ( .A(n22597), .Z(n24472) );
  BUF_X1 U19356 ( .A(n22610), .Z(n24406) );
  BUF_X1 U19357 ( .A(n22605), .Z(n24430) );
  BUF_X1 U19358 ( .A(n22593), .Z(n24492) );
  BUF_X1 U19359 ( .A(n22595), .Z(n24480) );
  BUF_X1 U19360 ( .A(n22597), .Z(n24468) );
  BUF_X1 U19361 ( .A(n22610), .Z(n24402) );
  BUF_X1 U19362 ( .A(n22605), .Z(n24426) );
  BUF_X1 U19363 ( .A(n22593), .Z(n24493) );
  BUF_X1 U19364 ( .A(n22595), .Z(n24481) );
  BUF_X1 U19365 ( .A(n22597), .Z(n24469) );
  BUF_X1 U19366 ( .A(n22610), .Z(n24403) );
  BUF_X1 U19367 ( .A(n22605), .Z(n24427) );
  BUF_X1 U19368 ( .A(n22593), .Z(n24494) );
  BUF_X1 U19369 ( .A(n22595), .Z(n24482) );
  BUF_X1 U19370 ( .A(n22597), .Z(n24470) );
  BUF_X1 U19371 ( .A(n22610), .Z(n24404) );
  BUF_X1 U19372 ( .A(n22605), .Z(n24428) );
  BUF_X1 U19373 ( .A(n22593), .Z(n24495) );
  BUF_X1 U19374 ( .A(n22595), .Z(n24483) );
  BUF_X1 U19375 ( .A(n22597), .Z(n24471) );
  BUF_X1 U19376 ( .A(n22610), .Z(n24405) );
  BUF_X1 U19377 ( .A(n22605), .Z(n24429) );
  BUF_X1 U19378 ( .A(n21311), .Z(n24768) );
  BUF_X1 U19379 ( .A(n21316), .Z(n24744) );
  BUF_X1 U19380 ( .A(n21321), .Z(n24720) );
  BUF_X1 U19381 ( .A(n21326), .Z(n24696) );
  BUF_X1 U19382 ( .A(n21335), .Z(n24672) );
  BUF_X1 U19383 ( .A(n21340), .Z(n24648) );
  BUF_X1 U19384 ( .A(n21345), .Z(n24624) );
  BUF_X1 U19385 ( .A(n21350), .Z(n24600) );
  BUF_X1 U19386 ( .A(n21311), .Z(n24769) );
  BUF_X1 U19387 ( .A(n21316), .Z(n24745) );
  BUF_X1 U19388 ( .A(n21321), .Z(n24721) );
  BUF_X1 U19389 ( .A(n21326), .Z(n24697) );
  BUF_X1 U19390 ( .A(n21335), .Z(n24673) );
  BUF_X1 U19391 ( .A(n21340), .Z(n24649) );
  BUF_X1 U19392 ( .A(n21345), .Z(n24625) );
  BUF_X1 U19393 ( .A(n21350), .Z(n24601) );
  BUF_X1 U19394 ( .A(n21311), .Z(n24770) );
  BUF_X1 U19395 ( .A(n21316), .Z(n24746) );
  BUF_X1 U19396 ( .A(n21321), .Z(n24722) );
  BUF_X1 U19397 ( .A(n21326), .Z(n24698) );
  BUF_X1 U19398 ( .A(n21335), .Z(n24674) );
  BUF_X1 U19399 ( .A(n21340), .Z(n24650) );
  BUF_X1 U19400 ( .A(n21345), .Z(n24626) );
  BUF_X1 U19401 ( .A(n21350), .Z(n24602) );
  BUF_X1 U19402 ( .A(n21311), .Z(n24771) );
  BUF_X1 U19403 ( .A(n21316), .Z(n24747) );
  BUF_X1 U19404 ( .A(n21321), .Z(n24723) );
  BUF_X1 U19405 ( .A(n21326), .Z(n24699) );
  BUF_X1 U19406 ( .A(n21335), .Z(n24675) );
  BUF_X1 U19407 ( .A(n21340), .Z(n24651) );
  BUF_X1 U19408 ( .A(n21345), .Z(n24627) );
  BUF_X1 U19409 ( .A(n21350), .Z(n24603) );
  BUF_X1 U19410 ( .A(n21311), .Z(n24772) );
  BUF_X1 U19411 ( .A(n21316), .Z(n24748) );
  BUF_X1 U19412 ( .A(n21321), .Z(n24724) );
  BUF_X1 U19413 ( .A(n21326), .Z(n24700) );
  BUF_X1 U19414 ( .A(n21335), .Z(n24676) );
  BUF_X1 U19415 ( .A(n21340), .Z(n24652) );
  BUF_X1 U19416 ( .A(n21345), .Z(n24628) );
  BUF_X1 U19417 ( .A(n21350), .Z(n24604) );
  BUF_X1 U19418 ( .A(n22596), .Z(n24478) );
  BUF_X1 U19419 ( .A(n22611), .Z(n24400) );
  BUF_X1 U19420 ( .A(n22606), .Z(n24424) );
  BUF_X1 U19421 ( .A(n22596), .Z(n24474) );
  BUF_X1 U19422 ( .A(n22611), .Z(n24396) );
  BUF_X1 U19423 ( .A(n22606), .Z(n24420) );
  BUF_X1 U19424 ( .A(n22596), .Z(n24475) );
  BUF_X1 U19425 ( .A(n22611), .Z(n24397) );
  BUF_X1 U19426 ( .A(n22606), .Z(n24421) );
  BUF_X1 U19427 ( .A(n22596), .Z(n24476) );
  BUF_X1 U19428 ( .A(n22611), .Z(n24398) );
  BUF_X1 U19429 ( .A(n22606), .Z(n24422) );
  BUF_X1 U19430 ( .A(n22596), .Z(n24477) );
  BUF_X1 U19431 ( .A(n22611), .Z(n24399) );
  BUF_X1 U19432 ( .A(n22606), .Z(n24423) );
  NAND2_X1 U19433 ( .A1(n23754), .A2(n23755), .ZN(n22594) );
  NAND2_X1 U19434 ( .A1(n23739), .A2(n23744), .ZN(n22574) );
  BUF_X1 U19435 ( .A(n22569), .Z(n24592) );
  BUF_X1 U19436 ( .A(n22584), .Z(n24520) );
  BUF_X1 U19437 ( .A(n22579), .Z(n24544) );
  BUF_X1 U19438 ( .A(n22569), .Z(n24588) );
  BUF_X1 U19439 ( .A(n22584), .Z(n24516) );
  BUF_X1 U19440 ( .A(n22579), .Z(n24540) );
  BUF_X1 U19441 ( .A(n22569), .Z(n24589) );
  BUF_X1 U19442 ( .A(n22584), .Z(n24517) );
  BUF_X1 U19443 ( .A(n22579), .Z(n24541) );
  BUF_X1 U19444 ( .A(n22569), .Z(n24590) );
  BUF_X1 U19445 ( .A(n22584), .Z(n24518) );
  BUF_X1 U19446 ( .A(n22579), .Z(n24542) );
  BUF_X1 U19447 ( .A(n22569), .Z(n24591) );
  BUF_X1 U19448 ( .A(n22584), .Z(n24519) );
  BUF_X1 U19449 ( .A(n22579), .Z(n24543) );
  BUF_X1 U19450 ( .A(n22568), .Z(n24594) );
  BUF_X1 U19451 ( .A(n22583), .Z(n24522) );
  BUF_X1 U19452 ( .A(n22573), .Z(n24570) );
  BUF_X1 U19453 ( .A(n22578), .Z(n24546) );
  BUF_X1 U19454 ( .A(n25556), .Z(n25564) );
  AND2_X1 U19455 ( .A1(n23739), .A2(n23740), .ZN(n22571) );
  AND2_X1 U19456 ( .A1(n23739), .A2(n23737), .ZN(n22577) );
  AND2_X1 U19457 ( .A1(n23739), .A2(n23747), .ZN(n22602) );
  BUF_X1 U19458 ( .A(n21189), .Z(n25534) );
  OAI21_X1 U19459 ( .B1(n21253), .B2(n21254), .A(n25562), .ZN(n21189) );
  BUF_X1 U19460 ( .A(n21296), .Z(n24815) );
  BUF_X1 U19461 ( .A(n21296), .Z(n24816) );
  INV_X1 U19462 ( .A(n24987), .ZN(n25003) );
  INV_X1 U19463 ( .A(n25208), .ZN(n25224) );
  INV_X1 U19464 ( .A(n25140), .ZN(n25156) );
  INV_X1 U19465 ( .A(n24885), .ZN(n24901) );
  INV_X1 U19466 ( .A(n25072), .ZN(n25088) );
  INV_X1 U19467 ( .A(n25004), .ZN(n25020) );
  INV_X1 U19468 ( .A(n24902), .ZN(n24918) );
  INV_X1 U19469 ( .A(n24834), .ZN(n24850) );
  INV_X1 U19470 ( .A(n25055), .ZN(n25071) );
  INV_X1 U19471 ( .A(n25191), .ZN(n25207) );
  INV_X1 U19472 ( .A(n25174), .ZN(n25190) );
  INV_X1 U19473 ( .A(n25089), .ZN(n25105) );
  INV_X1 U19474 ( .A(n25038), .ZN(n25054) );
  INV_X1 U19475 ( .A(n25021), .ZN(n25037) );
  INV_X1 U19476 ( .A(n24851), .ZN(n24867) );
  INV_X1 U19477 ( .A(n24868), .ZN(n24884) );
  INV_X1 U19478 ( .A(n24919), .ZN(n24935) );
  INV_X1 U19479 ( .A(n24936), .ZN(n24952) );
  INV_X1 U19480 ( .A(n24953), .ZN(n24969) );
  INV_X1 U19481 ( .A(n24970), .ZN(n24986) );
  INV_X1 U19482 ( .A(n25106), .ZN(n25122) );
  INV_X1 U19483 ( .A(n25123), .ZN(n25139) );
  INV_X1 U19484 ( .A(n25157), .ZN(n25173) );
  INV_X1 U19485 ( .A(n25225), .ZN(n25241) );
  INV_X1 U19486 ( .A(n25242), .ZN(n25258) );
  INV_X1 U19487 ( .A(n25310), .ZN(n25326) );
  INV_X1 U19488 ( .A(n25293), .ZN(n25309) );
  INV_X1 U19489 ( .A(n25327), .ZN(n25344) );
  INV_X1 U19490 ( .A(n25259), .ZN(n25275) );
  INV_X1 U19491 ( .A(n25276), .ZN(n25292) );
  OAI22_X1 U19492 ( .A1(n21151), .A2(n24497), .B1(n20525), .B2(n24491), .ZN(
        n22663) );
  OAI22_X1 U19493 ( .A1(n21150), .A2(n24497), .B1(n20524), .B2(n24491), .ZN(
        n22645) );
  OAI22_X1 U19494 ( .A1(n21148), .A2(n24497), .B1(n20523), .B2(n24491), .ZN(
        n22627) );
  OAI22_X1 U19495 ( .A1(n21149), .A2(n24497), .B1(n20522), .B2(n24491), .ZN(
        n22592) );
  OAI22_X1 U19496 ( .A1(n19271), .A2(n24485), .B1(n20261), .B2(n24479), .ZN(
        n22662) );
  OAI22_X1 U19497 ( .A1(n19270), .A2(n24485), .B1(n20260), .B2(n24479), .ZN(
        n22644) );
  OAI22_X1 U19498 ( .A1(n19269), .A2(n24485), .B1(n20259), .B2(n24479), .ZN(
        n22626) );
  OAI22_X1 U19499 ( .A1(n19268), .A2(n24485), .B1(n20258), .B2(n24479), .ZN(
        n22591) );
  OAI22_X1 U19500 ( .A1(n20542), .A2(n24473), .B1(n19207), .B2(n24467), .ZN(
        n22661) );
  OAI22_X1 U19501 ( .A1(n20541), .A2(n24473), .B1(n19206), .B2(n24467), .ZN(
        n22643) );
  OAI22_X1 U19502 ( .A1(n20540), .A2(n24473), .B1(n19205), .B2(n24467), .ZN(
        n22625) );
  OAI22_X1 U19503 ( .A1(n20539), .A2(n24473), .B1(n19204), .B2(n24467), .ZN(
        n22590) );
  OAI22_X1 U19504 ( .A1(n21159), .A2(n24496), .B1(n20698), .B2(n24490), .ZN(
        n22807) );
  OAI22_X1 U19505 ( .A1(n21158), .A2(n24496), .B1(n20697), .B2(n24490), .ZN(
        n22789) );
  OAI22_X1 U19506 ( .A1(n21157), .A2(n24496), .B1(n20696), .B2(n24490), .ZN(
        n22771) );
  OAI22_X1 U19507 ( .A1(n21156), .A2(n24496), .B1(n20695), .B2(n24490), .ZN(
        n22753) );
  OAI22_X1 U19508 ( .A1(n21155), .A2(n24496), .B1(n20694), .B2(n24490), .ZN(
        n22735) );
  OAI22_X1 U19509 ( .A1(n21154), .A2(n24496), .B1(n20693), .B2(n24490), .ZN(
        n22717) );
  OAI22_X1 U19510 ( .A1(n21153), .A2(n24496), .B1(n20692), .B2(n24490), .ZN(
        n22699) );
  OAI22_X1 U19511 ( .A1(n21152), .A2(n24496), .B1(n20691), .B2(n24490), .ZN(
        n22681) );
  OAI22_X1 U19512 ( .A1(n21187), .A2(n24492), .B1(n20846), .B2(n24486), .ZN(
        n23753) );
  OAI22_X1 U19513 ( .A1(n21147), .A2(n24492), .B1(n20845), .B2(n24486), .ZN(
        n23725) );
  OAI22_X1 U19514 ( .A1(n21186), .A2(n24492), .B1(n20844), .B2(n24486), .ZN(
        n23707) );
  OAI22_X1 U19515 ( .A1(n21185), .A2(n24492), .B1(n20843), .B2(n24486), .ZN(
        n23689) );
  OAI22_X1 U19516 ( .A1(n21184), .A2(n24492), .B1(n20842), .B2(n24486), .ZN(
        n23671) );
  OAI22_X1 U19517 ( .A1(n21183), .A2(n24492), .B1(n20841), .B2(n24486), .ZN(
        n23653) );
  OAI22_X1 U19518 ( .A1(n21182), .A2(n24492), .B1(n20840), .B2(n24486), .ZN(
        n23635) );
  OAI22_X1 U19519 ( .A1(n21181), .A2(n24492), .B1(n20839), .B2(n24486), .ZN(
        n23617) );
  OAI22_X1 U19520 ( .A1(n21180), .A2(n24492), .B1(n20838), .B2(n24486), .ZN(
        n23599) );
  OAI22_X1 U19521 ( .A1(n21179), .A2(n24492), .B1(n20837), .B2(n24486), .ZN(
        n23581) );
  OAI22_X1 U19522 ( .A1(n21178), .A2(n24492), .B1(n20836), .B2(n24486), .ZN(
        n23563) );
  OAI22_X1 U19523 ( .A1(n21177), .A2(n24492), .B1(n20835), .B2(n24486), .ZN(
        n23545) );
  OAI22_X1 U19524 ( .A1(n21176), .A2(n24493), .B1(n20834), .B2(n24487), .ZN(
        n23527) );
  OAI22_X1 U19525 ( .A1(n21175), .A2(n24493), .B1(n20833), .B2(n24487), .ZN(
        n23509) );
  OAI22_X1 U19526 ( .A1(n21174), .A2(n24493), .B1(n20832), .B2(n24487), .ZN(
        n23491) );
  OAI22_X1 U19527 ( .A1(n21173), .A2(n24493), .B1(n20831), .B2(n24487), .ZN(
        n23473) );
  OAI22_X1 U19528 ( .A1(n21172), .A2(n24493), .B1(n20830), .B2(n24487), .ZN(
        n23455) );
  OAI22_X1 U19529 ( .A1(n21171), .A2(n24493), .B1(n20829), .B2(n24487), .ZN(
        n23437) );
  OAI22_X1 U19530 ( .A1(n21170), .A2(n24493), .B1(n20828), .B2(n24487), .ZN(
        n23419) );
  OAI22_X1 U19531 ( .A1(n21169), .A2(n24493), .B1(n20827), .B2(n24487), .ZN(
        n23401) );
  OAI22_X1 U19532 ( .A1(n21168), .A2(n24493), .B1(n20826), .B2(n24487), .ZN(
        n23383) );
  OAI22_X1 U19533 ( .A1(n21167), .A2(n24493), .B1(n20825), .B2(n24487), .ZN(
        n23365) );
  OAI22_X1 U19534 ( .A1(n21166), .A2(n24493), .B1(n20824), .B2(n24487), .ZN(
        n23347) );
  OAI22_X1 U19535 ( .A1(n21165), .A2(n24493), .B1(n20823), .B2(n24487), .ZN(
        n23329) );
  OAI22_X1 U19536 ( .A1(n21164), .A2(n24494), .B1(n20726), .B2(n24488), .ZN(
        n23311) );
  OAI22_X1 U19537 ( .A1(n21163), .A2(n24494), .B1(n20725), .B2(n24488), .ZN(
        n23293) );
  OAI22_X1 U19538 ( .A1(n21162), .A2(n24494), .B1(n20724), .B2(n24488), .ZN(
        n23275) );
  OAI22_X1 U19539 ( .A1(n21161), .A2(n24494), .B1(n20723), .B2(n24488), .ZN(
        n23257) );
  OAI22_X1 U19540 ( .A1(n21160), .A2(n24494), .B1(n20722), .B2(n24488), .ZN(
        n23239) );
  OAI22_X1 U19541 ( .A1(n20998), .A2(n24471), .B1(n19227), .B2(n24465), .ZN(
        n23021) );
  OAI22_X1 U19542 ( .A1(n20997), .A2(n24471), .B1(n19226), .B2(n24465), .ZN(
        n23003) );
  OAI22_X1 U19543 ( .A1(n20996), .A2(n24471), .B1(n19225), .B2(n24465), .ZN(
        n22985) );
  OAI22_X1 U19544 ( .A1(n20995), .A2(n24471), .B1(n19224), .B2(n24465), .ZN(
        n22967) );
  OAI22_X1 U19545 ( .A1(n20994), .A2(n24471), .B1(n19223), .B2(n24465), .ZN(
        n22949) );
  OAI22_X1 U19546 ( .A1(n20993), .A2(n24471), .B1(n19222), .B2(n24465), .ZN(
        n22931) );
  OAI22_X1 U19547 ( .A1(n20992), .A2(n24471), .B1(n19221), .B2(n24465), .ZN(
        n22913) );
  OAI22_X1 U19548 ( .A1(n20991), .A2(n24471), .B1(n19220), .B2(n24465), .ZN(
        n22895) );
  OAI22_X1 U19549 ( .A1(n20990), .A2(n24472), .B1(n19219), .B2(n24466), .ZN(
        n22877) );
  OAI22_X1 U19550 ( .A1(n20989), .A2(n24472), .B1(n19218), .B2(n24466), .ZN(
        n22859) );
  OAI22_X1 U19551 ( .A1(n20988), .A2(n24472), .B1(n19217), .B2(n24466), .ZN(
        n22841) );
  OAI22_X1 U19552 ( .A1(n20987), .A2(n24472), .B1(n19216), .B2(n24466), .ZN(
        n22823) );
  OAI22_X1 U19553 ( .A1(n20986), .A2(n24472), .B1(n19215), .B2(n24466), .ZN(
        n22805) );
  OAI22_X1 U19554 ( .A1(n20985), .A2(n24472), .B1(n19214), .B2(n24466), .ZN(
        n22787) );
  OAI22_X1 U19555 ( .A1(n20984), .A2(n24472), .B1(n19213), .B2(n24466), .ZN(
        n22769) );
  OAI22_X1 U19556 ( .A1(n20983), .A2(n24472), .B1(n19212), .B2(n24466), .ZN(
        n22751) );
  OAI22_X1 U19557 ( .A1(n20982), .A2(n24472), .B1(n19211), .B2(n24466), .ZN(
        n22733) );
  OAI22_X1 U19558 ( .A1(n20981), .A2(n24472), .B1(n19210), .B2(n24466), .ZN(
        n22715) );
  OAI22_X1 U19559 ( .A1(n20980), .A2(n24472), .B1(n19209), .B2(n24466), .ZN(
        n22697) );
  OAI22_X1 U19560 ( .A1(n20979), .A2(n24472), .B1(n19208), .B2(n24466), .ZN(
        n22679) );
  OAI22_X1 U19561 ( .A1(n21122), .A2(n24468), .B1(n19267), .B2(n24462), .ZN(
        n23751) );
  OAI22_X1 U19562 ( .A1(n21121), .A2(n24468), .B1(n19266), .B2(n24462), .ZN(
        n23723) );
  OAI22_X1 U19563 ( .A1(n21120), .A2(n24468), .B1(n19265), .B2(n24462), .ZN(
        n23705) );
  OAI22_X1 U19564 ( .A1(n21119), .A2(n24468), .B1(n19264), .B2(n24462), .ZN(
        n23687) );
  OAI22_X1 U19565 ( .A1(n21118), .A2(n24468), .B1(n19263), .B2(n24462), .ZN(
        n23669) );
  OAI22_X1 U19566 ( .A1(n21117), .A2(n24468), .B1(n19262), .B2(n24462), .ZN(
        n23651) );
  OAI22_X1 U19567 ( .A1(n21116), .A2(n24468), .B1(n19261), .B2(n24462), .ZN(
        n23633) );
  OAI22_X1 U19568 ( .A1(n21115), .A2(n24468), .B1(n19260), .B2(n24462), .ZN(
        n23615) );
  OAI22_X1 U19569 ( .A1(n21114), .A2(n24468), .B1(n19259), .B2(n24462), .ZN(
        n23597) );
  OAI22_X1 U19570 ( .A1(n21113), .A2(n24468), .B1(n19258), .B2(n24462), .ZN(
        n23579) );
  OAI22_X1 U19571 ( .A1(n21112), .A2(n24468), .B1(n19257), .B2(n24462), .ZN(
        n23561) );
  OAI22_X1 U19572 ( .A1(n21111), .A2(n24468), .B1(n19256), .B2(n24462), .ZN(
        n23543) );
  OAI22_X1 U19573 ( .A1(n21110), .A2(n24469), .B1(n19255), .B2(n24463), .ZN(
        n23525) );
  OAI22_X1 U19574 ( .A1(n21109), .A2(n24469), .B1(n19254), .B2(n24463), .ZN(
        n23507) );
  OAI22_X1 U19575 ( .A1(n21108), .A2(n24469), .B1(n19253), .B2(n24463), .ZN(
        n23489) );
  OAI22_X1 U19576 ( .A1(n21107), .A2(n24469), .B1(n19252), .B2(n24463), .ZN(
        n23471) );
  OAI22_X1 U19577 ( .A1(n21106), .A2(n24469), .B1(n19251), .B2(n24463), .ZN(
        n23453) );
  OAI22_X1 U19578 ( .A1(n21105), .A2(n24469), .B1(n19250), .B2(n24463), .ZN(
        n23435) );
  OAI22_X1 U19579 ( .A1(n21104), .A2(n24469), .B1(n19249), .B2(n24463), .ZN(
        n23417) );
  OAI22_X1 U19580 ( .A1(n21103), .A2(n24469), .B1(n19248), .B2(n24463), .ZN(
        n23399) );
  OAI22_X1 U19581 ( .A1(n21102), .A2(n24469), .B1(n19247), .B2(n24463), .ZN(
        n23381) );
  OAI22_X1 U19582 ( .A1(n21101), .A2(n24469), .B1(n19246), .B2(n24463), .ZN(
        n23363) );
  OAI22_X1 U19583 ( .A1(n21100), .A2(n24469), .B1(n19245), .B2(n24463), .ZN(
        n23345) );
  OAI22_X1 U19584 ( .A1(n21099), .A2(n24469), .B1(n19244), .B2(n24463), .ZN(
        n23327) );
  OAI22_X1 U19585 ( .A1(n21014), .A2(n24470), .B1(n19243), .B2(n24464), .ZN(
        n23309) );
  OAI22_X1 U19586 ( .A1(n21013), .A2(n24470), .B1(n19242), .B2(n24464), .ZN(
        n23291) );
  OAI22_X1 U19587 ( .A1(n21012), .A2(n24470), .B1(n19241), .B2(n24464), .ZN(
        n23273) );
  OAI22_X1 U19588 ( .A1(n21011), .A2(n24470), .B1(n19240), .B2(n24464), .ZN(
        n23255) );
  OAI22_X1 U19589 ( .A1(n21010), .A2(n24470), .B1(n19239), .B2(n24464), .ZN(
        n23237) );
  OAI22_X1 U19590 ( .A1(n21009), .A2(n24470), .B1(n19238), .B2(n24464), .ZN(
        n23219) );
  OAI22_X1 U19591 ( .A1(n21008), .A2(n24470), .B1(n19237), .B2(n24464), .ZN(
        n23201) );
  OAI22_X1 U19592 ( .A1(n21007), .A2(n24470), .B1(n19236), .B2(n24464), .ZN(
        n23183) );
  OAI22_X1 U19593 ( .A1(n21006), .A2(n24470), .B1(n19235), .B2(n24464), .ZN(
        n23165) );
  OAI22_X1 U19594 ( .A1(n21005), .A2(n24470), .B1(n19234), .B2(n24464), .ZN(
        n23147) );
  OAI22_X1 U19595 ( .A1(n21004), .A2(n24470), .B1(n19233), .B2(n24464), .ZN(
        n23129) );
  OAI22_X1 U19596 ( .A1(n21003), .A2(n24470), .B1(n19232), .B2(n24464), .ZN(
        n23111) );
  OAI22_X1 U19597 ( .A1(n21002), .A2(n24471), .B1(n19231), .B2(n24465), .ZN(
        n23093) );
  OAI22_X1 U19598 ( .A1(n21001), .A2(n24471), .B1(n19230), .B2(n24465), .ZN(
        n23075) );
  OAI22_X1 U19599 ( .A1(n21000), .A2(n24471), .B1(n19229), .B2(n24465), .ZN(
        n23057) );
  OAI22_X1 U19600 ( .A1(n20999), .A2(n24471), .B1(n19228), .B2(n24465), .ZN(
        n23039) );
  OAI22_X1 U19601 ( .A1(n19291), .A2(n24483), .B1(n20357), .B2(n24477), .ZN(
        n23022) );
  OAI22_X1 U19602 ( .A1(n19290), .A2(n24483), .B1(n20356), .B2(n24477), .ZN(
        n23004) );
  OAI22_X1 U19603 ( .A1(n19289), .A2(n24483), .B1(n20355), .B2(n24477), .ZN(
        n22986) );
  OAI22_X1 U19604 ( .A1(n19288), .A2(n24483), .B1(n20354), .B2(n24477), .ZN(
        n22968) );
  OAI22_X1 U19605 ( .A1(n19287), .A2(n24483), .B1(n20353), .B2(n24477), .ZN(
        n22950) );
  OAI22_X1 U19606 ( .A1(n19286), .A2(n24483), .B1(n20352), .B2(n24477), .ZN(
        n22932) );
  OAI22_X1 U19607 ( .A1(n19285), .A2(n24483), .B1(n20351), .B2(n24477), .ZN(
        n22914) );
  OAI22_X1 U19608 ( .A1(n19284), .A2(n24483), .B1(n20350), .B2(n24477), .ZN(
        n22896) );
  OAI22_X1 U19609 ( .A1(n19283), .A2(n24484), .B1(n20349), .B2(n24478), .ZN(
        n22878) );
  OAI22_X1 U19610 ( .A1(n19282), .A2(n24484), .B1(n20348), .B2(n24478), .ZN(
        n22860) );
  OAI22_X1 U19611 ( .A1(n19281), .A2(n24484), .B1(n20347), .B2(n24478), .ZN(
        n22842) );
  OAI22_X1 U19612 ( .A1(n19280), .A2(n24484), .B1(n20346), .B2(n24478), .ZN(
        n22824) );
  OAI22_X1 U19613 ( .A1(n19279), .A2(n24484), .B1(n20345), .B2(n24478), .ZN(
        n22806) );
  OAI22_X1 U19614 ( .A1(n19278), .A2(n24484), .B1(n20344), .B2(n24478), .ZN(
        n22788) );
  OAI22_X1 U19615 ( .A1(n19277), .A2(n24484), .B1(n20343), .B2(n24478), .ZN(
        n22770) );
  OAI22_X1 U19616 ( .A1(n19276), .A2(n24484), .B1(n20342), .B2(n24478), .ZN(
        n22752) );
  OAI22_X1 U19617 ( .A1(n19275), .A2(n24484), .B1(n20341), .B2(n24478), .ZN(
        n22734) );
  OAI22_X1 U19618 ( .A1(n19274), .A2(n24484), .B1(n20340), .B2(n24478), .ZN(
        n22716) );
  OAI22_X1 U19619 ( .A1(n19273), .A2(n24484), .B1(n20339), .B2(n24478), .ZN(
        n22698) );
  OAI22_X1 U19620 ( .A1(n19272), .A2(n24484), .B1(n20338), .B2(n24478), .ZN(
        n22680) );
  OAI22_X1 U19621 ( .A1(n19331), .A2(n24480), .B1(n20445), .B2(n24474), .ZN(
        n23752) );
  OAI22_X1 U19622 ( .A1(n19330), .A2(n24480), .B1(n20444), .B2(n24474), .ZN(
        n23724) );
  OAI22_X1 U19623 ( .A1(n19329), .A2(n24480), .B1(n20443), .B2(n24474), .ZN(
        n23706) );
  OAI22_X1 U19624 ( .A1(n19328), .A2(n24480), .B1(n20442), .B2(n24474), .ZN(
        n23688) );
  OAI22_X1 U19625 ( .A1(n19327), .A2(n24480), .B1(n20441), .B2(n24474), .ZN(
        n23670) );
  OAI22_X1 U19626 ( .A1(n19326), .A2(n24480), .B1(n20440), .B2(n24474), .ZN(
        n23652) );
  OAI22_X1 U19627 ( .A1(n19325), .A2(n24480), .B1(n20439), .B2(n24474), .ZN(
        n23634) );
  OAI22_X1 U19628 ( .A1(n19324), .A2(n24480), .B1(n20438), .B2(n24474), .ZN(
        n23616) );
  OAI22_X1 U19629 ( .A1(n19323), .A2(n24480), .B1(n20437), .B2(n24474), .ZN(
        n23598) );
  OAI22_X1 U19630 ( .A1(n19322), .A2(n24480), .B1(n20436), .B2(n24474), .ZN(
        n23580) );
  OAI22_X1 U19631 ( .A1(n19321), .A2(n24480), .B1(n20435), .B2(n24474), .ZN(
        n23562) );
  OAI22_X1 U19632 ( .A1(n19320), .A2(n24480), .B1(n20434), .B2(n24474), .ZN(
        n23544) );
  OAI22_X1 U19633 ( .A1(n19319), .A2(n24481), .B1(n20433), .B2(n24475), .ZN(
        n23526) );
  OAI22_X1 U19634 ( .A1(n19318), .A2(n24481), .B1(n20432), .B2(n24475), .ZN(
        n23508) );
  OAI22_X1 U19635 ( .A1(n19317), .A2(n24481), .B1(n20431), .B2(n24475), .ZN(
        n23490) );
  OAI22_X1 U19636 ( .A1(n19316), .A2(n24481), .B1(n20430), .B2(n24475), .ZN(
        n23472) );
  OAI22_X1 U19637 ( .A1(n19315), .A2(n24481), .B1(n20429), .B2(n24475), .ZN(
        n23454) );
  OAI22_X1 U19638 ( .A1(n19314), .A2(n24481), .B1(n20428), .B2(n24475), .ZN(
        n23436) );
  OAI22_X1 U19639 ( .A1(n19313), .A2(n24481), .B1(n20427), .B2(n24475), .ZN(
        n23418) );
  OAI22_X1 U19640 ( .A1(n19312), .A2(n24481), .B1(n20426), .B2(n24475), .ZN(
        n23400) );
  OAI22_X1 U19641 ( .A1(n19311), .A2(n24481), .B1(n20425), .B2(n24475), .ZN(
        n23382) );
  OAI22_X1 U19642 ( .A1(n19310), .A2(n24481), .B1(n20424), .B2(n24475), .ZN(
        n23364) );
  OAI22_X1 U19643 ( .A1(n19309), .A2(n24481), .B1(n20423), .B2(n24475), .ZN(
        n23346) );
  OAI22_X1 U19644 ( .A1(n19308), .A2(n24481), .B1(n20422), .B2(n24475), .ZN(
        n23328) );
  OAI22_X1 U19645 ( .A1(n19307), .A2(n24482), .B1(n20373), .B2(n24476), .ZN(
        n23310) );
  OAI22_X1 U19646 ( .A1(n19306), .A2(n24482), .B1(n20372), .B2(n24476), .ZN(
        n23292) );
  OAI22_X1 U19647 ( .A1(n19305), .A2(n24482), .B1(n20371), .B2(n24476), .ZN(
        n23274) );
  OAI22_X1 U19648 ( .A1(n19304), .A2(n24482), .B1(n20370), .B2(n24476), .ZN(
        n23256) );
  OAI22_X1 U19649 ( .A1(n19303), .A2(n24482), .B1(n20369), .B2(n24476), .ZN(
        n23238) );
  OAI22_X1 U19650 ( .A1(n19302), .A2(n24482), .B1(n20368), .B2(n24476), .ZN(
        n23220) );
  OAI22_X1 U19651 ( .A1(n19301), .A2(n24482), .B1(n20367), .B2(n24476), .ZN(
        n23202) );
  OAI22_X1 U19652 ( .A1(n19300), .A2(n24482), .B1(n20366), .B2(n24476), .ZN(
        n23184) );
  OAI22_X1 U19653 ( .A1(n19299), .A2(n24482), .B1(n20365), .B2(n24476), .ZN(
        n23166) );
  OAI22_X1 U19654 ( .A1(n19298), .A2(n24482), .B1(n20364), .B2(n24476), .ZN(
        n23148) );
  OAI22_X1 U19655 ( .A1(n19297), .A2(n24482), .B1(n20363), .B2(n24476), .ZN(
        n23130) );
  OAI22_X1 U19656 ( .A1(n19296), .A2(n24482), .B1(n20362), .B2(n24476), .ZN(
        n23112) );
  OAI22_X1 U19657 ( .A1(n19295), .A2(n24483), .B1(n20361), .B2(n24477), .ZN(
        n23094) );
  OAI22_X1 U19658 ( .A1(n19294), .A2(n24483), .B1(n20360), .B2(n24477), .ZN(
        n23076) );
  OAI22_X1 U19659 ( .A1(n19293), .A2(n24483), .B1(n20359), .B2(n24477), .ZN(
        n23058) );
  OAI22_X1 U19660 ( .A1(n19292), .A2(n24483), .B1(n20358), .B2(n24477), .ZN(
        n23040) );
  OAI22_X1 U19661 ( .A1(n25330), .A2(n25345), .B1(n25328), .B2(n21187), .ZN(
        n6980) );
  OAI22_X1 U19662 ( .A1(n25330), .A2(n25351), .B1(n25329), .B2(n21186), .ZN(
        n6982) );
  OAI22_X1 U19663 ( .A1(n25330), .A2(n25354), .B1(n25329), .B2(n21185), .ZN(
        n6983) );
  OAI22_X1 U19664 ( .A1(n25330), .A2(n25357), .B1(n25329), .B2(n21184), .ZN(
        n6984) );
  OAI22_X1 U19665 ( .A1(n25331), .A2(n25360), .B1(n25329), .B2(n21183), .ZN(
        n6985) );
  OAI22_X1 U19666 ( .A1(n25331), .A2(n25363), .B1(n25329), .B2(n21182), .ZN(
        n6986) );
  OAI22_X1 U19667 ( .A1(n25331), .A2(n25366), .B1(n25329), .B2(n21181), .ZN(
        n6987) );
  OAI22_X1 U19668 ( .A1(n25331), .A2(n25369), .B1(n25329), .B2(n21180), .ZN(
        n6988) );
  OAI22_X1 U19669 ( .A1(n25331), .A2(n25372), .B1(n25329), .B2(n21179), .ZN(
        n6989) );
  OAI22_X1 U19670 ( .A1(n25332), .A2(n25375), .B1(n25329), .B2(n21178), .ZN(
        n6990) );
  OAI22_X1 U19671 ( .A1(n25332), .A2(n25378), .B1(n25329), .B2(n21177), .ZN(
        n6991) );
  OAI22_X1 U19672 ( .A1(n25332), .A2(n25381), .B1(n25329), .B2(n21176), .ZN(
        n6992) );
  OAI22_X1 U19673 ( .A1(n25332), .A2(n25384), .B1(n25329), .B2(n21175), .ZN(
        n6993) );
  OAI22_X1 U19674 ( .A1(n25332), .A2(n25387), .B1(n25329), .B2(n21174), .ZN(
        n6994) );
  OAI22_X1 U19675 ( .A1(n25333), .A2(n25390), .B1(n25328), .B2(n21173), .ZN(
        n6995) );
  OAI22_X1 U19676 ( .A1(n25333), .A2(n25393), .B1(n25328), .B2(n21172), .ZN(
        n6996) );
  OAI22_X1 U19677 ( .A1(n25333), .A2(n25396), .B1(n25328), .B2(n21171), .ZN(
        n6997) );
  OAI22_X1 U19678 ( .A1(n25333), .A2(n25399), .B1(n25328), .B2(n21170), .ZN(
        n6998) );
  OAI22_X1 U19679 ( .A1(n25333), .A2(n25402), .B1(n25328), .B2(n21169), .ZN(
        n6999) );
  OAI22_X1 U19680 ( .A1(n25334), .A2(n25405), .B1(n25328), .B2(n21168), .ZN(
        n7000) );
  OAI22_X1 U19681 ( .A1(n25334), .A2(n25408), .B1(n25328), .B2(n21167), .ZN(
        n7001) );
  OAI22_X1 U19682 ( .A1(n25334), .A2(n25411), .B1(n25328), .B2(n21166), .ZN(
        n7002) );
  OAI22_X1 U19683 ( .A1(n25334), .A2(n25414), .B1(n25328), .B2(n21165), .ZN(
        n7003) );
  OAI22_X1 U19684 ( .A1(n25334), .A2(n25417), .B1(n25328), .B2(n21164), .ZN(
        n7004) );
  OAI22_X1 U19685 ( .A1(n25335), .A2(n25420), .B1(n25328), .B2(n21163), .ZN(
        n7005) );
  OAI22_X1 U19686 ( .A1(n25335), .A2(n25423), .B1(n25328), .B2(n21162), .ZN(
        n7006) );
  OAI22_X1 U19687 ( .A1(n25335), .A2(n25426), .B1(n25328), .B2(n21161), .ZN(
        n7007) );
  OAI22_X1 U19688 ( .A1(n25335), .A2(n25429), .B1(n25327), .B2(n21160), .ZN(
        n7008) );
  OAI22_X1 U19689 ( .A1(n25340), .A2(n25501), .B1(n25329), .B2(n21159), .ZN(
        n7032) );
  OAI22_X1 U19690 ( .A1(n25340), .A2(n25504), .B1(n25328), .B2(n21158), .ZN(
        n7033) );
  OAI22_X1 U19691 ( .A1(n25340), .A2(n25507), .B1(n25327), .B2(n21157), .ZN(
        n7034) );
  OAI22_X1 U19692 ( .A1(n25341), .A2(n25510), .B1(n25329), .B2(n21156), .ZN(
        n7035) );
  OAI22_X1 U19693 ( .A1(n25341), .A2(n25513), .B1(n25328), .B2(n21155), .ZN(
        n7036) );
  OAI22_X1 U19694 ( .A1(n25341), .A2(n25516), .B1(n25327), .B2(n21154), .ZN(
        n7037) );
  OAI22_X1 U19695 ( .A1(n25341), .A2(n25519), .B1(n25329), .B2(n21153), .ZN(
        n7038) );
  OAI22_X1 U19696 ( .A1(n25341), .A2(n25522), .B1(n25328), .B2(n21152), .ZN(
        n7039) );
  OAI22_X1 U19697 ( .A1(n25342), .A2(n25525), .B1(n25327), .B2(n21151), .ZN(
        n7040) );
  OAI22_X1 U19698 ( .A1(n25342), .A2(n25528), .B1(n25329), .B2(n21150), .ZN(
        n7041) );
  OAI22_X1 U19699 ( .A1(n25342), .A2(n25551), .B1(n25328), .B2(n21149), .ZN(
        n7043) );
  OAI22_X1 U19700 ( .A1(n25342), .A2(n25531), .B1(n25327), .B2(n21148), .ZN(
        n7042) );
  OAI22_X1 U19701 ( .A1(n24990), .A2(n25346), .B1(n24988), .B2(n21146), .ZN(
        n5700) );
  OAI22_X1 U19702 ( .A1(n24990), .A2(n25349), .B1(n24988), .B2(n21145), .ZN(
        n5701) );
  OAI22_X1 U19703 ( .A1(n24990), .A2(n25352), .B1(n24988), .B2(n21144), .ZN(
        n5702) );
  OAI22_X1 U19704 ( .A1(n24990), .A2(n25355), .B1(n24988), .B2(n21143), .ZN(
        n5703) );
  OAI22_X1 U19705 ( .A1(n24990), .A2(n25358), .B1(n24988), .B2(n21142), .ZN(
        n5704) );
  OAI22_X1 U19706 ( .A1(n24991), .A2(n25361), .B1(n24988), .B2(n21141), .ZN(
        n5705) );
  OAI22_X1 U19707 ( .A1(n24991), .A2(n25364), .B1(n24988), .B2(n21140), .ZN(
        n5706) );
  OAI22_X1 U19708 ( .A1(n24991), .A2(n25367), .B1(n24988), .B2(n21139), .ZN(
        n5707) );
  OAI22_X1 U19709 ( .A1(n24991), .A2(n25370), .B1(n24988), .B2(n21138), .ZN(
        n5708) );
  OAI22_X1 U19710 ( .A1(n24991), .A2(n25373), .B1(n24988), .B2(n21137), .ZN(
        n5709) );
  OAI22_X1 U19711 ( .A1(n24992), .A2(n25376), .B1(n24988), .B2(n21136), .ZN(
        n5710) );
  OAI22_X1 U19712 ( .A1(n24992), .A2(n25379), .B1(n24988), .B2(n21135), .ZN(
        n5711) );
  OAI22_X1 U19713 ( .A1(n24992), .A2(n25382), .B1(n24989), .B2(n21134), .ZN(
        n5712) );
  OAI22_X1 U19714 ( .A1(n24992), .A2(n25385), .B1(n24989), .B2(n21133), .ZN(
        n5713) );
  OAI22_X1 U19715 ( .A1(n24992), .A2(n25388), .B1(n24989), .B2(n21132), .ZN(
        n5714) );
  OAI22_X1 U19716 ( .A1(n24993), .A2(n25391), .B1(n24989), .B2(n21131), .ZN(
        n5715) );
  OAI22_X1 U19717 ( .A1(n24993), .A2(n25394), .B1(n24989), .B2(n21130), .ZN(
        n5716) );
  OAI22_X1 U19718 ( .A1(n24993), .A2(n25397), .B1(n24989), .B2(n21129), .ZN(
        n5717) );
  OAI22_X1 U19719 ( .A1(n24993), .A2(n25400), .B1(n24989), .B2(n21128), .ZN(
        n5718) );
  OAI22_X1 U19720 ( .A1(n24993), .A2(n25403), .B1(n24989), .B2(n21127), .ZN(
        n5719) );
  OAI22_X1 U19721 ( .A1(n24994), .A2(n25406), .B1(n24989), .B2(n21126), .ZN(
        n5720) );
  OAI22_X1 U19722 ( .A1(n24994), .A2(n25409), .B1(n24989), .B2(n21125), .ZN(
        n5721) );
  OAI22_X1 U19723 ( .A1(n24994), .A2(n25412), .B1(n24989), .B2(n21124), .ZN(
        n5722) );
  OAI22_X1 U19724 ( .A1(n24994), .A2(n25415), .B1(n24989), .B2(n21123), .ZN(
        n5723) );
  OAI22_X1 U19725 ( .A1(n25228), .A2(n25345), .B1(n25226), .B2(n21122), .ZN(
        n6596) );
  OAI22_X1 U19726 ( .A1(n25228), .A2(n25348), .B1(n25226), .B2(n21121), .ZN(
        n6597) );
  OAI22_X1 U19727 ( .A1(n25228), .A2(n25351), .B1(n25226), .B2(n21120), .ZN(
        n6598) );
  OAI22_X1 U19728 ( .A1(n25228), .A2(n25354), .B1(n25226), .B2(n21119), .ZN(
        n6599) );
  OAI22_X1 U19729 ( .A1(n25228), .A2(n25357), .B1(n25226), .B2(n21118), .ZN(
        n6600) );
  OAI22_X1 U19730 ( .A1(n25229), .A2(n25360), .B1(n25226), .B2(n21117), .ZN(
        n6601) );
  OAI22_X1 U19731 ( .A1(n25229), .A2(n25363), .B1(n25226), .B2(n21116), .ZN(
        n6602) );
  OAI22_X1 U19732 ( .A1(n25229), .A2(n25366), .B1(n25226), .B2(n21115), .ZN(
        n6603) );
  OAI22_X1 U19733 ( .A1(n25229), .A2(n25369), .B1(n25226), .B2(n21114), .ZN(
        n6604) );
  OAI22_X1 U19734 ( .A1(n25229), .A2(n25372), .B1(n25226), .B2(n21113), .ZN(
        n6605) );
  OAI22_X1 U19735 ( .A1(n25230), .A2(n25375), .B1(n25226), .B2(n21112), .ZN(
        n6606) );
  OAI22_X1 U19736 ( .A1(n25230), .A2(n25378), .B1(n25226), .B2(n21111), .ZN(
        n6607) );
  OAI22_X1 U19737 ( .A1(n25230), .A2(n25381), .B1(n25227), .B2(n21110), .ZN(
        n6608) );
  OAI22_X1 U19738 ( .A1(n25230), .A2(n25384), .B1(n25227), .B2(n21109), .ZN(
        n6609) );
  OAI22_X1 U19739 ( .A1(n25230), .A2(n25387), .B1(n25227), .B2(n21108), .ZN(
        n6610) );
  OAI22_X1 U19740 ( .A1(n25231), .A2(n25390), .B1(n25227), .B2(n21107), .ZN(
        n6611) );
  OAI22_X1 U19741 ( .A1(n25231), .A2(n25393), .B1(n25227), .B2(n21106), .ZN(
        n6612) );
  OAI22_X1 U19742 ( .A1(n25231), .A2(n25396), .B1(n25227), .B2(n21105), .ZN(
        n6613) );
  OAI22_X1 U19743 ( .A1(n25231), .A2(n25399), .B1(n25227), .B2(n21104), .ZN(
        n6614) );
  OAI22_X1 U19744 ( .A1(n25231), .A2(n25402), .B1(n25227), .B2(n21103), .ZN(
        n6615) );
  OAI22_X1 U19745 ( .A1(n25232), .A2(n25405), .B1(n25227), .B2(n21102), .ZN(
        n6616) );
  OAI22_X1 U19746 ( .A1(n25232), .A2(n25408), .B1(n25227), .B2(n21101), .ZN(
        n6617) );
  OAI22_X1 U19747 ( .A1(n25232), .A2(n25411), .B1(n25227), .B2(n21100), .ZN(
        n6618) );
  OAI22_X1 U19748 ( .A1(n25232), .A2(n25414), .B1(n25227), .B2(n21099), .ZN(
        n6619) );
  OAI22_X1 U19749 ( .A1(n25211), .A2(n25345), .B1(n25209), .B2(n21098), .ZN(
        n6532) );
  OAI22_X1 U19750 ( .A1(n25211), .A2(n25348), .B1(n25209), .B2(n21097), .ZN(
        n6533) );
  OAI22_X1 U19751 ( .A1(n25211), .A2(n25351), .B1(n25209), .B2(n21096), .ZN(
        n6534) );
  OAI22_X1 U19752 ( .A1(n25211), .A2(n25354), .B1(n25209), .B2(n21095), .ZN(
        n6535) );
  OAI22_X1 U19753 ( .A1(n25211), .A2(n25357), .B1(n25209), .B2(n21094), .ZN(
        n6536) );
  OAI22_X1 U19754 ( .A1(n25212), .A2(n25360), .B1(n25209), .B2(n21093), .ZN(
        n6537) );
  OAI22_X1 U19755 ( .A1(n25212), .A2(n25363), .B1(n25209), .B2(n21092), .ZN(
        n6538) );
  OAI22_X1 U19756 ( .A1(n25212), .A2(n25366), .B1(n25209), .B2(n21091), .ZN(
        n6539) );
  OAI22_X1 U19757 ( .A1(n25212), .A2(n25369), .B1(n25209), .B2(n21090), .ZN(
        n6540) );
  OAI22_X1 U19758 ( .A1(n25212), .A2(n25372), .B1(n25209), .B2(n21089), .ZN(
        n6541) );
  OAI22_X1 U19759 ( .A1(n25213), .A2(n25375), .B1(n25209), .B2(n21088), .ZN(
        n6542) );
  OAI22_X1 U19760 ( .A1(n25213), .A2(n25378), .B1(n25209), .B2(n21087), .ZN(
        n6543) );
  OAI22_X1 U19761 ( .A1(n25213), .A2(n25381), .B1(n25210), .B2(n21086), .ZN(
        n6544) );
  OAI22_X1 U19762 ( .A1(n25213), .A2(n25384), .B1(n25210), .B2(n21085), .ZN(
        n6545) );
  OAI22_X1 U19763 ( .A1(n25213), .A2(n25387), .B1(n25210), .B2(n21084), .ZN(
        n6546) );
  OAI22_X1 U19764 ( .A1(n25214), .A2(n25390), .B1(n25210), .B2(n21083), .ZN(
        n6547) );
  OAI22_X1 U19765 ( .A1(n25214), .A2(n25393), .B1(n25210), .B2(n21082), .ZN(
        n6548) );
  OAI22_X1 U19766 ( .A1(n25214), .A2(n25396), .B1(n25210), .B2(n21081), .ZN(
        n6549) );
  OAI22_X1 U19767 ( .A1(n25214), .A2(n25399), .B1(n25210), .B2(n21080), .ZN(
        n6550) );
  OAI22_X1 U19768 ( .A1(n25214), .A2(n25402), .B1(n25210), .B2(n21079), .ZN(
        n6551) );
  OAI22_X1 U19769 ( .A1(n25215), .A2(n25405), .B1(n25210), .B2(n21078), .ZN(
        n6552) );
  OAI22_X1 U19770 ( .A1(n25215), .A2(n25408), .B1(n25210), .B2(n21077), .ZN(
        n6553) );
  OAI22_X1 U19771 ( .A1(n25215), .A2(n25411), .B1(n25210), .B2(n21076), .ZN(
        n6554) );
  OAI22_X1 U19772 ( .A1(n25215), .A2(n25414), .B1(n25210), .B2(n21075), .ZN(
        n6555) );
  OAI22_X1 U19773 ( .A1(n25143), .A2(n25346), .B1(n25141), .B2(n21074), .ZN(
        n6276) );
  OAI22_X1 U19774 ( .A1(n25143), .A2(n25349), .B1(n25141), .B2(n21073), .ZN(
        n6277) );
  OAI22_X1 U19775 ( .A1(n25143), .A2(n25352), .B1(n25141), .B2(n21072), .ZN(
        n6278) );
  OAI22_X1 U19776 ( .A1(n25143), .A2(n25355), .B1(n25141), .B2(n21071), .ZN(
        n6279) );
  OAI22_X1 U19777 ( .A1(n25143), .A2(n25358), .B1(n25141), .B2(n21070), .ZN(
        n6280) );
  OAI22_X1 U19778 ( .A1(n25144), .A2(n25361), .B1(n25141), .B2(n21069), .ZN(
        n6281) );
  OAI22_X1 U19779 ( .A1(n25144), .A2(n25364), .B1(n25141), .B2(n21068), .ZN(
        n6282) );
  OAI22_X1 U19780 ( .A1(n25144), .A2(n25367), .B1(n25141), .B2(n21067), .ZN(
        n6283) );
  OAI22_X1 U19781 ( .A1(n25144), .A2(n25370), .B1(n25141), .B2(n21066), .ZN(
        n6284) );
  OAI22_X1 U19782 ( .A1(n25144), .A2(n25373), .B1(n25141), .B2(n21065), .ZN(
        n6285) );
  OAI22_X1 U19783 ( .A1(n25145), .A2(n25376), .B1(n25141), .B2(n21064), .ZN(
        n6286) );
  OAI22_X1 U19784 ( .A1(n25145), .A2(n25379), .B1(n25141), .B2(n21063), .ZN(
        n6287) );
  OAI22_X1 U19785 ( .A1(n25145), .A2(n25382), .B1(n25142), .B2(n21062), .ZN(
        n6288) );
  OAI22_X1 U19786 ( .A1(n25145), .A2(n25385), .B1(n25142), .B2(n21061), .ZN(
        n6289) );
  OAI22_X1 U19787 ( .A1(n25145), .A2(n25388), .B1(n25142), .B2(n21060), .ZN(
        n6290) );
  OAI22_X1 U19788 ( .A1(n25146), .A2(n25391), .B1(n25142), .B2(n21059), .ZN(
        n6291) );
  OAI22_X1 U19789 ( .A1(n25146), .A2(n25394), .B1(n25142), .B2(n21058), .ZN(
        n6292) );
  OAI22_X1 U19790 ( .A1(n25146), .A2(n25397), .B1(n25142), .B2(n21057), .ZN(
        n6293) );
  OAI22_X1 U19791 ( .A1(n25146), .A2(n25400), .B1(n25142), .B2(n21056), .ZN(
        n6294) );
  OAI22_X1 U19792 ( .A1(n25146), .A2(n25403), .B1(n25142), .B2(n21055), .ZN(
        n6295) );
  OAI22_X1 U19793 ( .A1(n25147), .A2(n25406), .B1(n25142), .B2(n21054), .ZN(
        n6296) );
  OAI22_X1 U19794 ( .A1(n25147), .A2(n25409), .B1(n25142), .B2(n21053), .ZN(
        n6297) );
  OAI22_X1 U19795 ( .A1(n25147), .A2(n25412), .B1(n25142), .B2(n21052), .ZN(
        n6298) );
  OAI22_X1 U19796 ( .A1(n25147), .A2(n25415), .B1(n25142), .B2(n21051), .ZN(
        n6299) );
  OAI22_X1 U19797 ( .A1(n25245), .A2(n25345), .B1(n25243), .B2(n20846), .ZN(
        n6660) );
  OAI22_X1 U19798 ( .A1(n25245), .A2(n25348), .B1(n25243), .B2(n20845), .ZN(
        n6661) );
  OAI22_X1 U19799 ( .A1(n25245), .A2(n25351), .B1(n25243), .B2(n20844), .ZN(
        n6662) );
  OAI22_X1 U19800 ( .A1(n25245), .A2(n25354), .B1(n25243), .B2(n20843), .ZN(
        n6663) );
  OAI22_X1 U19801 ( .A1(n25245), .A2(n25357), .B1(n25243), .B2(n20842), .ZN(
        n6664) );
  OAI22_X1 U19802 ( .A1(n25246), .A2(n25360), .B1(n25243), .B2(n20841), .ZN(
        n6665) );
  OAI22_X1 U19803 ( .A1(n25246), .A2(n25363), .B1(n25243), .B2(n20840), .ZN(
        n6666) );
  OAI22_X1 U19804 ( .A1(n25246), .A2(n25366), .B1(n25243), .B2(n20839), .ZN(
        n6667) );
  OAI22_X1 U19805 ( .A1(n25246), .A2(n25369), .B1(n25243), .B2(n20838), .ZN(
        n6668) );
  OAI22_X1 U19806 ( .A1(n25246), .A2(n25372), .B1(n25243), .B2(n20837), .ZN(
        n6669) );
  OAI22_X1 U19807 ( .A1(n25247), .A2(n25375), .B1(n25243), .B2(n20836), .ZN(
        n6670) );
  OAI22_X1 U19808 ( .A1(n25247), .A2(n25378), .B1(n25243), .B2(n20835), .ZN(
        n6671) );
  OAI22_X1 U19809 ( .A1(n25247), .A2(n25381), .B1(n25244), .B2(n20834), .ZN(
        n6672) );
  OAI22_X1 U19810 ( .A1(n25247), .A2(n25384), .B1(n25244), .B2(n20833), .ZN(
        n6673) );
  OAI22_X1 U19811 ( .A1(n25247), .A2(n25387), .B1(n25244), .B2(n20832), .ZN(
        n6674) );
  OAI22_X1 U19812 ( .A1(n25248), .A2(n25390), .B1(n25244), .B2(n20831), .ZN(
        n6675) );
  OAI22_X1 U19813 ( .A1(n25248), .A2(n25393), .B1(n25244), .B2(n20830), .ZN(
        n6676) );
  OAI22_X1 U19814 ( .A1(n25248), .A2(n25396), .B1(n25244), .B2(n20829), .ZN(
        n6677) );
  OAI22_X1 U19815 ( .A1(n25248), .A2(n25399), .B1(n25244), .B2(n20828), .ZN(
        n6678) );
  OAI22_X1 U19816 ( .A1(n25248), .A2(n25402), .B1(n25244), .B2(n20827), .ZN(
        n6679) );
  OAI22_X1 U19817 ( .A1(n25249), .A2(n25405), .B1(n25244), .B2(n20826), .ZN(
        n6680) );
  OAI22_X1 U19818 ( .A1(n25249), .A2(n25408), .B1(n25244), .B2(n20825), .ZN(
        n6681) );
  OAI22_X1 U19819 ( .A1(n25249), .A2(n25411), .B1(n25244), .B2(n20824), .ZN(
        n6682) );
  OAI22_X1 U19820 ( .A1(n25249), .A2(n25414), .B1(n25244), .B2(n20823), .ZN(
        n6683) );
  OAI22_X1 U19821 ( .A1(n25075), .A2(n25346), .B1(n25073), .B2(n20822), .ZN(
        n6020) );
  OAI22_X1 U19822 ( .A1(n25075), .A2(n25349), .B1(n25073), .B2(n20821), .ZN(
        n6021) );
  OAI22_X1 U19823 ( .A1(n25075), .A2(n25352), .B1(n25073), .B2(n20820), .ZN(
        n6022) );
  OAI22_X1 U19824 ( .A1(n25075), .A2(n25355), .B1(n25073), .B2(n20819), .ZN(
        n6023) );
  OAI22_X1 U19825 ( .A1(n25075), .A2(n25358), .B1(n25073), .B2(n20818), .ZN(
        n6024) );
  OAI22_X1 U19826 ( .A1(n25076), .A2(n25361), .B1(n25073), .B2(n20817), .ZN(
        n6025) );
  OAI22_X1 U19827 ( .A1(n25076), .A2(n25364), .B1(n25073), .B2(n20816), .ZN(
        n6026) );
  OAI22_X1 U19828 ( .A1(n25076), .A2(n25367), .B1(n25073), .B2(n20815), .ZN(
        n6027) );
  OAI22_X1 U19829 ( .A1(n25076), .A2(n25370), .B1(n25073), .B2(n20814), .ZN(
        n6028) );
  OAI22_X1 U19830 ( .A1(n25076), .A2(n25373), .B1(n25073), .B2(n20813), .ZN(
        n6029) );
  OAI22_X1 U19831 ( .A1(n25077), .A2(n25376), .B1(n25073), .B2(n20812), .ZN(
        n6030) );
  OAI22_X1 U19832 ( .A1(n25077), .A2(n25379), .B1(n25073), .B2(n20811), .ZN(
        n6031) );
  OAI22_X1 U19833 ( .A1(n25077), .A2(n25382), .B1(n25074), .B2(n20810), .ZN(
        n6032) );
  OAI22_X1 U19834 ( .A1(n25077), .A2(n25385), .B1(n25074), .B2(n20809), .ZN(
        n6033) );
  OAI22_X1 U19835 ( .A1(n25077), .A2(n25388), .B1(n25074), .B2(n20808), .ZN(
        n6034) );
  OAI22_X1 U19836 ( .A1(n25078), .A2(n25391), .B1(n25074), .B2(n20807), .ZN(
        n6035) );
  OAI22_X1 U19837 ( .A1(n25078), .A2(n25394), .B1(n25074), .B2(n20806), .ZN(
        n6036) );
  OAI22_X1 U19838 ( .A1(n25078), .A2(n25397), .B1(n25074), .B2(n20805), .ZN(
        n6037) );
  OAI22_X1 U19839 ( .A1(n25078), .A2(n25400), .B1(n25074), .B2(n20804), .ZN(
        n6038) );
  OAI22_X1 U19840 ( .A1(n25078), .A2(n25403), .B1(n25074), .B2(n20803), .ZN(
        n6039) );
  OAI22_X1 U19841 ( .A1(n25079), .A2(n25406), .B1(n25074), .B2(n20802), .ZN(
        n6040) );
  OAI22_X1 U19842 ( .A1(n25079), .A2(n25409), .B1(n25074), .B2(n20801), .ZN(
        n6041) );
  OAI22_X1 U19843 ( .A1(n25079), .A2(n25412), .B1(n25074), .B2(n20800), .ZN(
        n6042) );
  OAI22_X1 U19844 ( .A1(n25079), .A2(n25415), .B1(n25074), .B2(n20799), .ZN(
        n6043) );
  OAI22_X1 U19845 ( .A1(n25007), .A2(n25346), .B1(n25005), .B2(n20798), .ZN(
        n5764) );
  OAI22_X1 U19846 ( .A1(n25007), .A2(n25349), .B1(n25005), .B2(n20797), .ZN(
        n5765) );
  OAI22_X1 U19847 ( .A1(n25007), .A2(n25352), .B1(n25005), .B2(n20796), .ZN(
        n5766) );
  OAI22_X1 U19848 ( .A1(n25007), .A2(n25355), .B1(n25005), .B2(n20795), .ZN(
        n5767) );
  OAI22_X1 U19849 ( .A1(n25007), .A2(n25358), .B1(n25005), .B2(n20794), .ZN(
        n5768) );
  OAI22_X1 U19850 ( .A1(n25008), .A2(n25361), .B1(n25005), .B2(n20793), .ZN(
        n5769) );
  OAI22_X1 U19851 ( .A1(n25008), .A2(n25364), .B1(n25005), .B2(n20792), .ZN(
        n5770) );
  OAI22_X1 U19852 ( .A1(n25008), .A2(n25367), .B1(n25005), .B2(n20791), .ZN(
        n5771) );
  OAI22_X1 U19853 ( .A1(n25008), .A2(n25370), .B1(n25005), .B2(n20790), .ZN(
        n5772) );
  OAI22_X1 U19854 ( .A1(n25008), .A2(n25373), .B1(n25005), .B2(n20789), .ZN(
        n5773) );
  OAI22_X1 U19855 ( .A1(n25009), .A2(n25376), .B1(n25005), .B2(n20788), .ZN(
        n5774) );
  OAI22_X1 U19856 ( .A1(n25009), .A2(n25379), .B1(n25005), .B2(n20787), .ZN(
        n5775) );
  OAI22_X1 U19857 ( .A1(n25009), .A2(n25382), .B1(n25006), .B2(n20786), .ZN(
        n5776) );
  OAI22_X1 U19858 ( .A1(n25009), .A2(n25385), .B1(n25006), .B2(n20785), .ZN(
        n5777) );
  OAI22_X1 U19859 ( .A1(n25009), .A2(n25388), .B1(n25006), .B2(n20784), .ZN(
        n5778) );
  OAI22_X1 U19860 ( .A1(n25010), .A2(n25391), .B1(n25006), .B2(n20783), .ZN(
        n5779) );
  OAI22_X1 U19861 ( .A1(n25010), .A2(n25394), .B1(n25006), .B2(n20782), .ZN(
        n5780) );
  OAI22_X1 U19862 ( .A1(n25010), .A2(n25397), .B1(n25006), .B2(n20781), .ZN(
        n5781) );
  OAI22_X1 U19863 ( .A1(n25010), .A2(n25400), .B1(n25006), .B2(n20780), .ZN(
        n5782) );
  OAI22_X1 U19864 ( .A1(n25010), .A2(n25403), .B1(n25006), .B2(n20779), .ZN(
        n5783) );
  OAI22_X1 U19865 ( .A1(n25011), .A2(n25406), .B1(n25006), .B2(n20778), .ZN(
        n5784) );
  OAI22_X1 U19866 ( .A1(n25011), .A2(n25409), .B1(n25006), .B2(n20777), .ZN(
        n5785) );
  OAI22_X1 U19867 ( .A1(n25011), .A2(n25412), .B1(n25006), .B2(n20776), .ZN(
        n5786) );
  OAI22_X1 U19868 ( .A1(n25011), .A2(n25415), .B1(n25006), .B2(n20775), .ZN(
        n5787) );
  OAI22_X1 U19869 ( .A1(n24905), .A2(n25347), .B1(n24903), .B2(n20774), .ZN(
        n5380) );
  OAI22_X1 U19870 ( .A1(n24905), .A2(n25350), .B1(n24903), .B2(n20773), .ZN(
        n5381) );
  OAI22_X1 U19871 ( .A1(n24905), .A2(n25353), .B1(n24903), .B2(n20772), .ZN(
        n5382) );
  OAI22_X1 U19872 ( .A1(n24905), .A2(n25356), .B1(n24903), .B2(n20771), .ZN(
        n5383) );
  OAI22_X1 U19873 ( .A1(n24905), .A2(n25359), .B1(n24903), .B2(n20770), .ZN(
        n5384) );
  OAI22_X1 U19874 ( .A1(n24906), .A2(n25362), .B1(n24903), .B2(n20769), .ZN(
        n5385) );
  OAI22_X1 U19875 ( .A1(n24906), .A2(n25365), .B1(n24903), .B2(n20768), .ZN(
        n5386) );
  OAI22_X1 U19876 ( .A1(n24906), .A2(n25368), .B1(n24903), .B2(n20767), .ZN(
        n5387) );
  OAI22_X1 U19877 ( .A1(n24906), .A2(n25371), .B1(n24903), .B2(n20766), .ZN(
        n5388) );
  OAI22_X1 U19878 ( .A1(n24906), .A2(n25374), .B1(n24903), .B2(n20765), .ZN(
        n5389) );
  OAI22_X1 U19879 ( .A1(n24907), .A2(n25377), .B1(n24903), .B2(n20764), .ZN(
        n5390) );
  OAI22_X1 U19880 ( .A1(n24907), .A2(n25380), .B1(n24903), .B2(n20763), .ZN(
        n5391) );
  OAI22_X1 U19881 ( .A1(n24907), .A2(n25383), .B1(n24904), .B2(n20762), .ZN(
        n5392) );
  OAI22_X1 U19882 ( .A1(n24907), .A2(n25386), .B1(n24904), .B2(n20761), .ZN(
        n5393) );
  OAI22_X1 U19883 ( .A1(n24907), .A2(n25389), .B1(n24904), .B2(n20760), .ZN(
        n5394) );
  OAI22_X1 U19884 ( .A1(n24908), .A2(n25392), .B1(n24904), .B2(n20759), .ZN(
        n5395) );
  OAI22_X1 U19885 ( .A1(n24908), .A2(n25395), .B1(n24904), .B2(n20758), .ZN(
        n5396) );
  OAI22_X1 U19886 ( .A1(n24908), .A2(n25398), .B1(n24904), .B2(n20757), .ZN(
        n5397) );
  OAI22_X1 U19887 ( .A1(n24908), .A2(n25401), .B1(n24904), .B2(n20756), .ZN(
        n5398) );
  OAI22_X1 U19888 ( .A1(n24908), .A2(n25404), .B1(n24904), .B2(n20755), .ZN(
        n5399) );
  OAI22_X1 U19889 ( .A1(n24909), .A2(n25407), .B1(n24904), .B2(n20754), .ZN(
        n5400) );
  OAI22_X1 U19890 ( .A1(n24909), .A2(n25410), .B1(n24904), .B2(n20753), .ZN(
        n5401) );
  OAI22_X1 U19891 ( .A1(n24909), .A2(n25413), .B1(n24904), .B2(n20752), .ZN(
        n5402) );
  OAI22_X1 U19892 ( .A1(n24909), .A2(n25416), .B1(n24904), .B2(n20751), .ZN(
        n5403) );
  OAI22_X1 U19893 ( .A1(n24837), .A2(n25347), .B1(n24835), .B2(n20750), .ZN(
        n5124) );
  OAI22_X1 U19894 ( .A1(n24837), .A2(n25350), .B1(n24835), .B2(n20749), .ZN(
        n5125) );
  OAI22_X1 U19895 ( .A1(n24837), .A2(n25353), .B1(n24835), .B2(n20748), .ZN(
        n5126) );
  OAI22_X1 U19896 ( .A1(n24837), .A2(n25356), .B1(n24835), .B2(n20747), .ZN(
        n5127) );
  OAI22_X1 U19897 ( .A1(n24837), .A2(n25359), .B1(n24835), .B2(n20746), .ZN(
        n5128) );
  OAI22_X1 U19898 ( .A1(n24838), .A2(n25362), .B1(n24835), .B2(n20745), .ZN(
        n5129) );
  OAI22_X1 U19899 ( .A1(n24838), .A2(n25365), .B1(n24835), .B2(n20744), .ZN(
        n5130) );
  OAI22_X1 U19900 ( .A1(n24838), .A2(n25368), .B1(n24835), .B2(n20743), .ZN(
        n5131) );
  OAI22_X1 U19901 ( .A1(n24838), .A2(n25371), .B1(n24835), .B2(n20742), .ZN(
        n5132) );
  OAI22_X1 U19902 ( .A1(n24838), .A2(n25374), .B1(n24835), .B2(n20741), .ZN(
        n5133) );
  OAI22_X1 U19903 ( .A1(n24839), .A2(n25377), .B1(n24835), .B2(n20740), .ZN(
        n5134) );
  OAI22_X1 U19904 ( .A1(n24839), .A2(n25380), .B1(n24835), .B2(n20739), .ZN(
        n5135) );
  OAI22_X1 U19905 ( .A1(n24839), .A2(n25383), .B1(n24836), .B2(n20738), .ZN(
        n5136) );
  OAI22_X1 U19906 ( .A1(n24839), .A2(n25386), .B1(n24836), .B2(n20737), .ZN(
        n5137) );
  OAI22_X1 U19907 ( .A1(n24839), .A2(n25389), .B1(n24836), .B2(n20736), .ZN(
        n5138) );
  OAI22_X1 U19908 ( .A1(n24840), .A2(n25392), .B1(n24836), .B2(n20735), .ZN(
        n5139) );
  OAI22_X1 U19909 ( .A1(n24840), .A2(n25395), .B1(n24836), .B2(n20734), .ZN(
        n5140) );
  OAI22_X1 U19910 ( .A1(n24840), .A2(n25398), .B1(n24836), .B2(n20733), .ZN(
        n5141) );
  OAI22_X1 U19911 ( .A1(n24840), .A2(n25401), .B1(n24836), .B2(n20732), .ZN(
        n5142) );
  OAI22_X1 U19912 ( .A1(n24840), .A2(n25404), .B1(n24836), .B2(n20731), .ZN(
        n5143) );
  OAI22_X1 U19913 ( .A1(n24841), .A2(n25407), .B1(n24836), .B2(n20730), .ZN(
        n5144) );
  OAI22_X1 U19914 ( .A1(n24841), .A2(n25410), .B1(n24836), .B2(n20729), .ZN(
        n5145) );
  OAI22_X1 U19915 ( .A1(n24841), .A2(n25413), .B1(n24836), .B2(n20728), .ZN(
        n5146) );
  OAI22_X1 U19916 ( .A1(n24841), .A2(n25416), .B1(n24836), .B2(n20727), .ZN(
        n5147) );
  OAI22_X1 U19917 ( .A1(n25058), .A2(n25346), .B1(n25056), .B2(n20505), .ZN(
        n5956) );
  OAI22_X1 U19918 ( .A1(n25058), .A2(n25349), .B1(n25056), .B2(n20504), .ZN(
        n5957) );
  OAI22_X1 U19919 ( .A1(n25058), .A2(n25352), .B1(n25056), .B2(n20503), .ZN(
        n5958) );
  OAI22_X1 U19920 ( .A1(n25058), .A2(n25355), .B1(n25056), .B2(n20502), .ZN(
        n5959) );
  OAI22_X1 U19921 ( .A1(n25058), .A2(n25358), .B1(n25056), .B2(n20501), .ZN(
        n5960) );
  OAI22_X1 U19922 ( .A1(n25059), .A2(n25361), .B1(n25056), .B2(n20500), .ZN(
        n5961) );
  OAI22_X1 U19923 ( .A1(n25059), .A2(n25364), .B1(n25056), .B2(n20499), .ZN(
        n5962) );
  OAI22_X1 U19924 ( .A1(n25059), .A2(n25367), .B1(n25056), .B2(n20498), .ZN(
        n5963) );
  OAI22_X1 U19925 ( .A1(n25059), .A2(n25370), .B1(n25056), .B2(n20497), .ZN(
        n5964) );
  OAI22_X1 U19926 ( .A1(n25059), .A2(n25373), .B1(n25056), .B2(n20496), .ZN(
        n5965) );
  OAI22_X1 U19927 ( .A1(n25060), .A2(n25376), .B1(n25056), .B2(n20495), .ZN(
        n5966) );
  OAI22_X1 U19928 ( .A1(n25060), .A2(n25379), .B1(n25056), .B2(n20494), .ZN(
        n5967) );
  OAI22_X1 U19929 ( .A1(n25060), .A2(n25382), .B1(n25057), .B2(n20493), .ZN(
        n5968) );
  OAI22_X1 U19930 ( .A1(n25060), .A2(n25385), .B1(n25057), .B2(n20492), .ZN(
        n5969) );
  OAI22_X1 U19931 ( .A1(n25060), .A2(n25388), .B1(n25057), .B2(n20491), .ZN(
        n5970) );
  OAI22_X1 U19932 ( .A1(n25061), .A2(n25391), .B1(n25057), .B2(n20490), .ZN(
        n5971) );
  OAI22_X1 U19933 ( .A1(n25061), .A2(n25394), .B1(n25057), .B2(n20489), .ZN(
        n5972) );
  OAI22_X1 U19934 ( .A1(n25061), .A2(n25397), .B1(n25057), .B2(n20488), .ZN(
        n5973) );
  OAI22_X1 U19935 ( .A1(n25061), .A2(n25400), .B1(n25057), .B2(n20487), .ZN(
        n5974) );
  OAI22_X1 U19936 ( .A1(n25061), .A2(n25403), .B1(n25057), .B2(n20486), .ZN(
        n5975) );
  OAI22_X1 U19937 ( .A1(n25062), .A2(n25406), .B1(n25057), .B2(n20485), .ZN(
        n5976) );
  OAI22_X1 U19938 ( .A1(n25062), .A2(n25409), .B1(n25057), .B2(n20484), .ZN(
        n5977) );
  OAI22_X1 U19939 ( .A1(n25062), .A2(n25412), .B1(n25057), .B2(n20483), .ZN(
        n5978) );
  OAI22_X1 U19940 ( .A1(n25062), .A2(n25415), .B1(n25057), .B2(n20482), .ZN(
        n5979) );
  OAI22_X1 U19941 ( .A1(n25313), .A2(n25345), .B1(n25311), .B2(n20445), .ZN(
        n6916) );
  OAI22_X1 U19942 ( .A1(n25313), .A2(n25348), .B1(n25311), .B2(n20444), .ZN(
        n6917) );
  OAI22_X1 U19943 ( .A1(n25313), .A2(n25351), .B1(n25311), .B2(n20443), .ZN(
        n6918) );
  OAI22_X1 U19944 ( .A1(n25313), .A2(n25354), .B1(n25311), .B2(n20442), .ZN(
        n6919) );
  OAI22_X1 U19945 ( .A1(n25313), .A2(n25357), .B1(n25311), .B2(n20441), .ZN(
        n6920) );
  OAI22_X1 U19946 ( .A1(n25314), .A2(n25360), .B1(n25311), .B2(n20440), .ZN(
        n6921) );
  OAI22_X1 U19947 ( .A1(n25314), .A2(n25363), .B1(n25311), .B2(n20439), .ZN(
        n6922) );
  OAI22_X1 U19948 ( .A1(n25314), .A2(n25366), .B1(n25311), .B2(n20438), .ZN(
        n6923) );
  OAI22_X1 U19949 ( .A1(n25314), .A2(n25369), .B1(n25311), .B2(n20437), .ZN(
        n6924) );
  OAI22_X1 U19950 ( .A1(n25314), .A2(n25372), .B1(n25311), .B2(n20436), .ZN(
        n6925) );
  OAI22_X1 U19951 ( .A1(n25315), .A2(n25375), .B1(n25311), .B2(n20435), .ZN(
        n6926) );
  OAI22_X1 U19952 ( .A1(n25315), .A2(n25378), .B1(n25311), .B2(n20434), .ZN(
        n6927) );
  OAI22_X1 U19953 ( .A1(n25315), .A2(n25381), .B1(n25312), .B2(n20433), .ZN(
        n6928) );
  OAI22_X1 U19954 ( .A1(n25315), .A2(n25384), .B1(n25312), .B2(n20432), .ZN(
        n6929) );
  OAI22_X1 U19955 ( .A1(n25315), .A2(n25387), .B1(n25312), .B2(n20431), .ZN(
        n6930) );
  OAI22_X1 U19956 ( .A1(n25316), .A2(n25390), .B1(n25312), .B2(n20430), .ZN(
        n6931) );
  OAI22_X1 U19957 ( .A1(n25316), .A2(n25393), .B1(n25312), .B2(n20429), .ZN(
        n6932) );
  OAI22_X1 U19958 ( .A1(n25316), .A2(n25396), .B1(n25312), .B2(n20428), .ZN(
        n6933) );
  OAI22_X1 U19959 ( .A1(n25316), .A2(n25399), .B1(n25312), .B2(n20427), .ZN(
        n6934) );
  OAI22_X1 U19960 ( .A1(n25316), .A2(n25402), .B1(n25312), .B2(n20426), .ZN(
        n6935) );
  OAI22_X1 U19961 ( .A1(n25317), .A2(n25405), .B1(n25312), .B2(n20425), .ZN(
        n6936) );
  OAI22_X1 U19962 ( .A1(n25317), .A2(n25408), .B1(n25312), .B2(n20424), .ZN(
        n6937) );
  OAI22_X1 U19963 ( .A1(n25317), .A2(n25411), .B1(n25312), .B2(n20423), .ZN(
        n6938) );
  OAI22_X1 U19964 ( .A1(n25317), .A2(n25414), .B1(n25312), .B2(n20422), .ZN(
        n6939) );
  OAI22_X1 U19965 ( .A1(n25194), .A2(n25345), .B1(n25192), .B2(n20421), .ZN(
        n6468) );
  OAI22_X1 U19966 ( .A1(n25194), .A2(n25348), .B1(n25192), .B2(n20420), .ZN(
        n6469) );
  OAI22_X1 U19967 ( .A1(n25194), .A2(n25351), .B1(n25192), .B2(n20419), .ZN(
        n6470) );
  OAI22_X1 U19968 ( .A1(n25194), .A2(n25354), .B1(n25192), .B2(n20418), .ZN(
        n6471) );
  OAI22_X1 U19969 ( .A1(n25194), .A2(n25357), .B1(n25192), .B2(n20417), .ZN(
        n6472) );
  OAI22_X1 U19970 ( .A1(n25195), .A2(n25360), .B1(n25192), .B2(n20416), .ZN(
        n6473) );
  OAI22_X1 U19971 ( .A1(n25195), .A2(n25363), .B1(n25192), .B2(n20415), .ZN(
        n6474) );
  OAI22_X1 U19972 ( .A1(n25195), .A2(n25366), .B1(n25192), .B2(n20414), .ZN(
        n6475) );
  OAI22_X1 U19973 ( .A1(n25195), .A2(n25369), .B1(n25192), .B2(n20413), .ZN(
        n6476) );
  OAI22_X1 U19974 ( .A1(n25195), .A2(n25372), .B1(n25192), .B2(n20412), .ZN(
        n6477) );
  OAI22_X1 U19975 ( .A1(n25196), .A2(n25375), .B1(n25192), .B2(n20411), .ZN(
        n6478) );
  OAI22_X1 U19976 ( .A1(n25196), .A2(n25378), .B1(n25192), .B2(n20410), .ZN(
        n6479) );
  OAI22_X1 U19977 ( .A1(n25196), .A2(n25381), .B1(n25193), .B2(n20409), .ZN(
        n6480) );
  OAI22_X1 U19978 ( .A1(n25196), .A2(n25384), .B1(n25193), .B2(n20408), .ZN(
        n6481) );
  OAI22_X1 U19979 ( .A1(n25196), .A2(n25387), .B1(n25193), .B2(n20407), .ZN(
        n6482) );
  OAI22_X1 U19980 ( .A1(n25197), .A2(n25390), .B1(n25193), .B2(n20406), .ZN(
        n6483) );
  OAI22_X1 U19981 ( .A1(n25197), .A2(n25393), .B1(n25193), .B2(n20405), .ZN(
        n6484) );
  OAI22_X1 U19982 ( .A1(n25197), .A2(n25396), .B1(n25193), .B2(n20404), .ZN(
        n6485) );
  OAI22_X1 U19983 ( .A1(n25197), .A2(n25399), .B1(n25193), .B2(n20403), .ZN(
        n6486) );
  OAI22_X1 U19984 ( .A1(n25197), .A2(n25402), .B1(n25193), .B2(n20402), .ZN(
        n6487) );
  OAI22_X1 U19985 ( .A1(n25198), .A2(n25405), .B1(n25193), .B2(n20401), .ZN(
        n6488) );
  OAI22_X1 U19986 ( .A1(n25198), .A2(n25408), .B1(n25193), .B2(n20400), .ZN(
        n6489) );
  OAI22_X1 U19987 ( .A1(n25198), .A2(n25411), .B1(n25193), .B2(n20399), .ZN(
        n6490) );
  OAI22_X1 U19988 ( .A1(n25198), .A2(n25414), .B1(n25193), .B2(n20398), .ZN(
        n6491) );
  OAI22_X1 U19989 ( .A1(n25296), .A2(n25345), .B1(n25294), .B2(n20397), .ZN(
        n6852) );
  OAI22_X1 U19990 ( .A1(n25296), .A2(n25348), .B1(n25294), .B2(n20396), .ZN(
        n6853) );
  OAI22_X1 U19991 ( .A1(n25296), .A2(n25351), .B1(n25294), .B2(n20395), .ZN(
        n6854) );
  OAI22_X1 U19992 ( .A1(n25296), .A2(n25354), .B1(n25294), .B2(n20394), .ZN(
        n6855) );
  OAI22_X1 U19993 ( .A1(n25296), .A2(n25357), .B1(n25294), .B2(n20393), .ZN(
        n6856) );
  OAI22_X1 U19994 ( .A1(n25297), .A2(n25360), .B1(n25294), .B2(n20392), .ZN(
        n6857) );
  OAI22_X1 U19995 ( .A1(n25297), .A2(n25363), .B1(n25294), .B2(n20391), .ZN(
        n6858) );
  OAI22_X1 U19996 ( .A1(n25297), .A2(n25366), .B1(n25294), .B2(n20390), .ZN(
        n6859) );
  OAI22_X1 U19997 ( .A1(n25297), .A2(n25369), .B1(n25294), .B2(n20389), .ZN(
        n6860) );
  OAI22_X1 U19998 ( .A1(n25297), .A2(n25372), .B1(n25294), .B2(n20388), .ZN(
        n6861) );
  OAI22_X1 U19999 ( .A1(n25298), .A2(n25375), .B1(n25294), .B2(n20387), .ZN(
        n6862) );
  OAI22_X1 U20000 ( .A1(n25298), .A2(n25378), .B1(n25294), .B2(n20386), .ZN(
        n6863) );
  OAI22_X1 U20001 ( .A1(n25298), .A2(n25381), .B1(n25295), .B2(n20385), .ZN(
        n6864) );
  OAI22_X1 U20002 ( .A1(n25298), .A2(n25384), .B1(n25295), .B2(n20384), .ZN(
        n6865) );
  OAI22_X1 U20003 ( .A1(n25298), .A2(n25387), .B1(n25295), .B2(n20383), .ZN(
        n6866) );
  OAI22_X1 U20004 ( .A1(n25299), .A2(n25390), .B1(n25295), .B2(n20382), .ZN(
        n6867) );
  OAI22_X1 U20005 ( .A1(n25299), .A2(n25393), .B1(n25295), .B2(n20381), .ZN(
        n6868) );
  OAI22_X1 U20006 ( .A1(n25299), .A2(n25396), .B1(n25295), .B2(n20380), .ZN(
        n6869) );
  OAI22_X1 U20007 ( .A1(n25299), .A2(n25399), .B1(n25295), .B2(n20379), .ZN(
        n6870) );
  OAI22_X1 U20008 ( .A1(n25299), .A2(n25402), .B1(n25295), .B2(n20378), .ZN(
        n6871) );
  OAI22_X1 U20009 ( .A1(n25300), .A2(n25405), .B1(n25295), .B2(n20377), .ZN(
        n6872) );
  OAI22_X1 U20010 ( .A1(n25300), .A2(n25408), .B1(n25295), .B2(n20376), .ZN(
        n6873) );
  OAI22_X1 U20011 ( .A1(n25300), .A2(n25411), .B1(n25295), .B2(n20375), .ZN(
        n6874) );
  OAI22_X1 U20012 ( .A1(n25300), .A2(n25414), .B1(n25295), .B2(n20374), .ZN(
        n6875) );
  OAI22_X1 U20013 ( .A1(n24871), .A2(n25347), .B1(n24869), .B2(n19737), .ZN(
        n5252) );
  OAI22_X1 U20014 ( .A1(n24871), .A2(n25350), .B1(n24869), .B2(n19736), .ZN(
        n5253) );
  OAI22_X1 U20015 ( .A1(n24871), .A2(n25353), .B1(n24869), .B2(n19735), .ZN(
        n5254) );
  OAI22_X1 U20016 ( .A1(n24871), .A2(n25356), .B1(n24869), .B2(n19734), .ZN(
        n5255) );
  OAI22_X1 U20017 ( .A1(n24871), .A2(n25359), .B1(n24869), .B2(n19733), .ZN(
        n5256) );
  OAI22_X1 U20018 ( .A1(n24872), .A2(n25362), .B1(n24869), .B2(n19732), .ZN(
        n5257) );
  OAI22_X1 U20019 ( .A1(n24872), .A2(n25365), .B1(n24869), .B2(n19731), .ZN(
        n5258) );
  OAI22_X1 U20020 ( .A1(n24872), .A2(n25368), .B1(n24869), .B2(n19730), .ZN(
        n5259) );
  OAI22_X1 U20021 ( .A1(n24872), .A2(n25371), .B1(n24869), .B2(n19729), .ZN(
        n5260) );
  OAI22_X1 U20022 ( .A1(n24872), .A2(n25374), .B1(n24869), .B2(n19728), .ZN(
        n5261) );
  OAI22_X1 U20023 ( .A1(n24873), .A2(n25377), .B1(n24869), .B2(n19727), .ZN(
        n5262) );
  OAI22_X1 U20024 ( .A1(n24873), .A2(n25380), .B1(n24869), .B2(n19726), .ZN(
        n5263) );
  OAI22_X1 U20025 ( .A1(n24873), .A2(n25383), .B1(n24870), .B2(n19725), .ZN(
        n5264) );
  OAI22_X1 U20026 ( .A1(n24873), .A2(n25386), .B1(n24870), .B2(n19724), .ZN(
        n5265) );
  OAI22_X1 U20027 ( .A1(n24873), .A2(n25389), .B1(n24870), .B2(n19723), .ZN(
        n5266) );
  OAI22_X1 U20028 ( .A1(n24874), .A2(n25392), .B1(n24870), .B2(n19722), .ZN(
        n5267) );
  OAI22_X1 U20029 ( .A1(n24874), .A2(n25395), .B1(n24870), .B2(n19721), .ZN(
        n5268) );
  OAI22_X1 U20030 ( .A1(n24874), .A2(n25398), .B1(n24870), .B2(n19720), .ZN(
        n5269) );
  OAI22_X1 U20031 ( .A1(n24874), .A2(n25401), .B1(n24870), .B2(n19719), .ZN(
        n5270) );
  OAI22_X1 U20032 ( .A1(n24874), .A2(n25404), .B1(n24870), .B2(n19718), .ZN(
        n5271) );
  OAI22_X1 U20033 ( .A1(n24875), .A2(n25407), .B1(n24870), .B2(n19717), .ZN(
        n5272) );
  OAI22_X1 U20034 ( .A1(n24875), .A2(n25410), .B1(n24870), .B2(n19716), .ZN(
        n5273) );
  OAI22_X1 U20035 ( .A1(n24875), .A2(n25413), .B1(n24870), .B2(n19715), .ZN(
        n5274) );
  OAI22_X1 U20036 ( .A1(n24875), .A2(n25416), .B1(n24870), .B2(n19714), .ZN(
        n5275) );
  OAI22_X1 U20037 ( .A1(n24939), .A2(n25347), .B1(n24937), .B2(n19707), .ZN(
        n5508) );
  OAI22_X1 U20038 ( .A1(n24939), .A2(n25350), .B1(n24937), .B2(n19706), .ZN(
        n5509) );
  OAI22_X1 U20039 ( .A1(n24939), .A2(n25353), .B1(n24937), .B2(n19705), .ZN(
        n5510) );
  OAI22_X1 U20040 ( .A1(n24939), .A2(n25356), .B1(n24937), .B2(n19704), .ZN(
        n5511) );
  OAI22_X1 U20041 ( .A1(n24939), .A2(n25359), .B1(n24937), .B2(n19703), .ZN(
        n5512) );
  OAI22_X1 U20042 ( .A1(n24940), .A2(n25362), .B1(n24937), .B2(n19702), .ZN(
        n5513) );
  OAI22_X1 U20043 ( .A1(n24940), .A2(n25365), .B1(n24937), .B2(n19701), .ZN(
        n5514) );
  OAI22_X1 U20044 ( .A1(n24940), .A2(n25368), .B1(n24937), .B2(n19700), .ZN(
        n5515) );
  OAI22_X1 U20045 ( .A1(n24940), .A2(n25371), .B1(n24937), .B2(n19699), .ZN(
        n5516) );
  OAI22_X1 U20046 ( .A1(n24940), .A2(n25374), .B1(n24937), .B2(n19698), .ZN(
        n5517) );
  OAI22_X1 U20047 ( .A1(n24941), .A2(n25377), .B1(n24937), .B2(n19697), .ZN(
        n5518) );
  OAI22_X1 U20048 ( .A1(n24941), .A2(n25380), .B1(n24937), .B2(n19696), .ZN(
        n5519) );
  OAI22_X1 U20049 ( .A1(n24941), .A2(n25383), .B1(n24938), .B2(n19695), .ZN(
        n5520) );
  OAI22_X1 U20050 ( .A1(n24941), .A2(n25386), .B1(n24938), .B2(n19694), .ZN(
        n5521) );
  OAI22_X1 U20051 ( .A1(n24941), .A2(n25389), .B1(n24938), .B2(n19693), .ZN(
        n5522) );
  OAI22_X1 U20052 ( .A1(n24942), .A2(n25392), .B1(n24938), .B2(n19692), .ZN(
        n5523) );
  OAI22_X1 U20053 ( .A1(n24942), .A2(n25395), .B1(n24938), .B2(n19691), .ZN(
        n5524) );
  OAI22_X1 U20054 ( .A1(n24942), .A2(n25398), .B1(n24938), .B2(n19690), .ZN(
        n5525) );
  OAI22_X1 U20055 ( .A1(n24942), .A2(n25401), .B1(n24938), .B2(n19689), .ZN(
        n5526) );
  OAI22_X1 U20056 ( .A1(n24942), .A2(n25404), .B1(n24938), .B2(n19688), .ZN(
        n5527) );
  OAI22_X1 U20057 ( .A1(n24943), .A2(n25407), .B1(n24938), .B2(n19687), .ZN(
        n5528) );
  OAI22_X1 U20058 ( .A1(n24943), .A2(n25410), .B1(n24938), .B2(n19686), .ZN(
        n5529) );
  OAI22_X1 U20059 ( .A1(n24943), .A2(n25413), .B1(n24938), .B2(n19685), .ZN(
        n5530) );
  OAI22_X1 U20060 ( .A1(n24943), .A2(n25416), .B1(n24938), .B2(n19684), .ZN(
        n5531) );
  OAI22_X1 U20061 ( .A1(n25279), .A2(n25345), .B1(n25277), .B2(n19395), .ZN(
        n6788) );
  OAI22_X1 U20062 ( .A1(n25279), .A2(n25348), .B1(n25277), .B2(n19394), .ZN(
        n6789) );
  OAI22_X1 U20063 ( .A1(n25279), .A2(n25351), .B1(n25277), .B2(n19393), .ZN(
        n6790) );
  OAI22_X1 U20064 ( .A1(n25279), .A2(n25354), .B1(n25277), .B2(n19392), .ZN(
        n6791) );
  OAI22_X1 U20065 ( .A1(n25279), .A2(n25357), .B1(n25277), .B2(n19391), .ZN(
        n6792) );
  OAI22_X1 U20066 ( .A1(n25280), .A2(n25360), .B1(n25277), .B2(n19390), .ZN(
        n6793) );
  OAI22_X1 U20067 ( .A1(n25280), .A2(n25363), .B1(n25277), .B2(n19389), .ZN(
        n6794) );
  OAI22_X1 U20068 ( .A1(n25280), .A2(n25366), .B1(n25277), .B2(n19388), .ZN(
        n6795) );
  OAI22_X1 U20069 ( .A1(n25280), .A2(n25369), .B1(n25277), .B2(n19387), .ZN(
        n6796) );
  OAI22_X1 U20070 ( .A1(n25280), .A2(n25372), .B1(n25277), .B2(n19386), .ZN(
        n6797) );
  OAI22_X1 U20071 ( .A1(n25281), .A2(n25375), .B1(n25277), .B2(n19385), .ZN(
        n6798) );
  OAI22_X1 U20072 ( .A1(n25281), .A2(n25378), .B1(n25277), .B2(n19384), .ZN(
        n6799) );
  OAI22_X1 U20073 ( .A1(n25281), .A2(n25381), .B1(n25278), .B2(n19383), .ZN(
        n6800) );
  OAI22_X1 U20074 ( .A1(n25281), .A2(n25384), .B1(n25278), .B2(n19382), .ZN(
        n6801) );
  OAI22_X1 U20075 ( .A1(n25281), .A2(n25387), .B1(n25278), .B2(n19381), .ZN(
        n6802) );
  OAI22_X1 U20076 ( .A1(n25282), .A2(n25390), .B1(n25278), .B2(n19380), .ZN(
        n6803) );
  OAI22_X1 U20077 ( .A1(n25282), .A2(n25393), .B1(n25278), .B2(n19379), .ZN(
        n6804) );
  OAI22_X1 U20078 ( .A1(n25282), .A2(n25396), .B1(n25278), .B2(n19378), .ZN(
        n6805) );
  OAI22_X1 U20079 ( .A1(n25282), .A2(n25399), .B1(n25278), .B2(n19377), .ZN(
        n6806) );
  OAI22_X1 U20080 ( .A1(n25282), .A2(n25402), .B1(n25278), .B2(n19376), .ZN(
        n6807) );
  OAI22_X1 U20081 ( .A1(n25283), .A2(n25405), .B1(n25278), .B2(n19375), .ZN(
        n6808) );
  OAI22_X1 U20082 ( .A1(n25283), .A2(n25408), .B1(n25278), .B2(n19374), .ZN(
        n6809) );
  OAI22_X1 U20083 ( .A1(n25283), .A2(n25411), .B1(n25278), .B2(n19373), .ZN(
        n6810) );
  OAI22_X1 U20084 ( .A1(n25283), .A2(n25414), .B1(n25278), .B2(n19372), .ZN(
        n6811) );
  OAI22_X1 U20085 ( .A1(n25537), .A2(n25345), .B1(n25535), .B2(n19331), .ZN(
        n7044) );
  OAI22_X1 U20086 ( .A1(n25537), .A2(n25348), .B1(n25535), .B2(n19330), .ZN(
        n7045) );
  OAI22_X1 U20087 ( .A1(n25537), .A2(n25351), .B1(n25535), .B2(n19329), .ZN(
        n7046) );
  OAI22_X1 U20088 ( .A1(n25537), .A2(n25354), .B1(n25535), .B2(n19328), .ZN(
        n7047) );
  OAI22_X1 U20089 ( .A1(n25537), .A2(n25357), .B1(n25535), .B2(n19327), .ZN(
        n7048) );
  OAI22_X1 U20090 ( .A1(n25538), .A2(n25360), .B1(n25535), .B2(n19326), .ZN(
        n7049) );
  OAI22_X1 U20091 ( .A1(n25538), .A2(n25363), .B1(n25535), .B2(n19325), .ZN(
        n7050) );
  OAI22_X1 U20092 ( .A1(n25538), .A2(n25366), .B1(n25535), .B2(n19324), .ZN(
        n7051) );
  OAI22_X1 U20093 ( .A1(n25538), .A2(n25369), .B1(n25535), .B2(n19323), .ZN(
        n7052) );
  OAI22_X1 U20094 ( .A1(n25538), .A2(n25372), .B1(n25535), .B2(n19322), .ZN(
        n7053) );
  OAI22_X1 U20095 ( .A1(n25539), .A2(n25375), .B1(n25535), .B2(n19321), .ZN(
        n7054) );
  OAI22_X1 U20096 ( .A1(n25539), .A2(n25378), .B1(n25535), .B2(n19320), .ZN(
        n7055) );
  OAI22_X1 U20097 ( .A1(n25539), .A2(n25381), .B1(n25536), .B2(n19319), .ZN(
        n7056) );
  OAI22_X1 U20098 ( .A1(n25539), .A2(n25384), .B1(n25536), .B2(n19318), .ZN(
        n7057) );
  OAI22_X1 U20099 ( .A1(n25539), .A2(n25387), .B1(n25536), .B2(n19317), .ZN(
        n7058) );
  OAI22_X1 U20100 ( .A1(n25540), .A2(n25390), .B1(n25536), .B2(n19316), .ZN(
        n7059) );
  OAI22_X1 U20101 ( .A1(n25540), .A2(n25393), .B1(n25536), .B2(n19315), .ZN(
        n7060) );
  OAI22_X1 U20102 ( .A1(n25540), .A2(n25396), .B1(n25536), .B2(n19314), .ZN(
        n7061) );
  OAI22_X1 U20103 ( .A1(n25540), .A2(n25399), .B1(n25536), .B2(n19313), .ZN(
        n7062) );
  OAI22_X1 U20104 ( .A1(n25540), .A2(n25402), .B1(n25536), .B2(n19312), .ZN(
        n7063) );
  OAI22_X1 U20105 ( .A1(n25541), .A2(n25405), .B1(n25536), .B2(n19311), .ZN(
        n7064) );
  OAI22_X1 U20106 ( .A1(n25541), .A2(n25408), .B1(n25536), .B2(n19310), .ZN(
        n7065) );
  OAI22_X1 U20107 ( .A1(n25541), .A2(n25411), .B1(n25536), .B2(n19309), .ZN(
        n7066) );
  OAI22_X1 U20108 ( .A1(n25541), .A2(n25414), .B1(n25536), .B2(n19308), .ZN(
        n7067) );
  OAI22_X1 U20109 ( .A1(n24994), .A2(n25418), .B1(n24988), .B2(n21050), .ZN(
        n5724) );
  OAI22_X1 U20110 ( .A1(n24995), .A2(n25421), .B1(n24989), .B2(n21049), .ZN(
        n5725) );
  OAI22_X1 U20111 ( .A1(n24995), .A2(n25424), .B1(n24987), .B2(n21048), .ZN(
        n5726) );
  OAI22_X1 U20112 ( .A1(n24995), .A2(n25427), .B1(n24988), .B2(n21047), .ZN(
        n5727) );
  OAI22_X1 U20113 ( .A1(n24995), .A2(n25430), .B1(n24989), .B2(n21046), .ZN(
        n5728) );
  OAI22_X1 U20114 ( .A1(n24995), .A2(n25433), .B1(n24987), .B2(n21045), .ZN(
        n5729) );
  OAI22_X1 U20115 ( .A1(n24996), .A2(n25436), .B1(n24988), .B2(n21044), .ZN(
        n5730) );
  OAI22_X1 U20116 ( .A1(n24996), .A2(n25439), .B1(n24989), .B2(n21043), .ZN(
        n5731) );
  OAI22_X1 U20117 ( .A1(n24996), .A2(n25442), .B1(n24987), .B2(n21042), .ZN(
        n5732) );
  OAI22_X1 U20118 ( .A1(n24996), .A2(n25445), .B1(n24988), .B2(n21041), .ZN(
        n5733) );
  OAI22_X1 U20119 ( .A1(n24996), .A2(n25448), .B1(n24989), .B2(n21040), .ZN(
        n5734) );
  OAI22_X1 U20120 ( .A1(n24997), .A2(n25451), .B1(n24987), .B2(n21039), .ZN(
        n5735) );
  OAI22_X1 U20121 ( .A1(n24997), .A2(n25454), .B1(n21285), .B2(n21038), .ZN(
        n5736) );
  OAI22_X1 U20122 ( .A1(n24997), .A2(n25457), .B1(n24987), .B2(n21037), .ZN(
        n5737) );
  OAI22_X1 U20123 ( .A1(n24997), .A2(n25460), .B1(n21285), .B2(n21036), .ZN(
        n5738) );
  OAI22_X1 U20124 ( .A1(n24997), .A2(n25463), .B1(n24987), .B2(n21035), .ZN(
        n5739) );
  OAI22_X1 U20125 ( .A1(n24998), .A2(n25466), .B1(n21285), .B2(n21034), .ZN(
        n5740) );
  OAI22_X1 U20126 ( .A1(n24998), .A2(n25469), .B1(n24987), .B2(n21033), .ZN(
        n5741) );
  OAI22_X1 U20127 ( .A1(n24998), .A2(n25472), .B1(n24988), .B2(n21032), .ZN(
        n5742) );
  OAI22_X1 U20128 ( .A1(n24998), .A2(n25475), .B1(n24989), .B2(n21031), .ZN(
        n5743) );
  OAI22_X1 U20129 ( .A1(n24998), .A2(n25478), .B1(n24987), .B2(n21030), .ZN(
        n5744) );
  OAI22_X1 U20130 ( .A1(n24999), .A2(n25481), .B1(n24987), .B2(n21029), .ZN(
        n5745) );
  OAI22_X1 U20131 ( .A1(n24999), .A2(n25484), .B1(n24988), .B2(n21028), .ZN(
        n5746) );
  OAI22_X1 U20132 ( .A1(n24999), .A2(n25487), .B1(n24989), .B2(n21027), .ZN(
        n5747) );
  OAI22_X1 U20133 ( .A1(n24999), .A2(n25490), .B1(n24987), .B2(n21026), .ZN(
        n5748) );
  OAI22_X1 U20134 ( .A1(n24999), .A2(n25493), .B1(n24987), .B2(n21025), .ZN(
        n5749) );
  OAI22_X1 U20135 ( .A1(n25000), .A2(n25496), .B1(n21285), .B2(n21024), .ZN(
        n5750) );
  OAI22_X1 U20136 ( .A1(n25000), .A2(n25499), .B1(n24987), .B2(n21023), .ZN(
        n5751) );
  OAI22_X1 U20137 ( .A1(n25000), .A2(n25502), .B1(n21285), .B2(n21022), .ZN(
        n5752) );
  OAI22_X1 U20138 ( .A1(n25000), .A2(n25505), .B1(n24987), .B2(n21021), .ZN(
        n5753) );
  OAI22_X1 U20139 ( .A1(n25000), .A2(n25508), .B1(n21285), .B2(n21020), .ZN(
        n5754) );
  OAI22_X1 U20140 ( .A1(n25001), .A2(n25511), .B1(n24987), .B2(n21019), .ZN(
        n5755) );
  OAI22_X1 U20141 ( .A1(n25001), .A2(n25514), .B1(n21285), .B2(n21018), .ZN(
        n5756) );
  OAI22_X1 U20142 ( .A1(n25001), .A2(n25517), .B1(n24987), .B2(n21017), .ZN(
        n5757) );
  OAI22_X1 U20143 ( .A1(n25001), .A2(n25520), .B1(n21285), .B2(n21016), .ZN(
        n5758) );
  OAI22_X1 U20144 ( .A1(n25001), .A2(n25523), .B1(n24987), .B2(n21015), .ZN(
        n5759) );
  OAI22_X1 U20145 ( .A1(n25232), .A2(n25417), .B1(n25226), .B2(n21014), .ZN(
        n6620) );
  OAI22_X1 U20146 ( .A1(n25233), .A2(n25420), .B1(n25227), .B2(n21013), .ZN(
        n6621) );
  OAI22_X1 U20147 ( .A1(n25233), .A2(n25423), .B1(n25225), .B2(n21012), .ZN(
        n6622) );
  OAI22_X1 U20148 ( .A1(n25233), .A2(n25426), .B1(n25226), .B2(n21011), .ZN(
        n6623) );
  OAI22_X1 U20149 ( .A1(n25233), .A2(n25429), .B1(n25227), .B2(n21010), .ZN(
        n6624) );
  OAI22_X1 U20150 ( .A1(n25233), .A2(n25432), .B1(n25225), .B2(n21009), .ZN(
        n6625) );
  OAI22_X1 U20151 ( .A1(n25234), .A2(n25435), .B1(n25226), .B2(n21008), .ZN(
        n6626) );
  OAI22_X1 U20152 ( .A1(n25234), .A2(n25438), .B1(n25227), .B2(n21007), .ZN(
        n6627) );
  OAI22_X1 U20153 ( .A1(n25234), .A2(n25441), .B1(n25225), .B2(n21006), .ZN(
        n6628) );
  OAI22_X1 U20154 ( .A1(n25234), .A2(n25444), .B1(n25226), .B2(n21005), .ZN(
        n6629) );
  OAI22_X1 U20155 ( .A1(n25234), .A2(n25447), .B1(n25227), .B2(n21004), .ZN(
        n6630) );
  OAI22_X1 U20156 ( .A1(n25235), .A2(n25450), .B1(n25225), .B2(n21003), .ZN(
        n6631) );
  OAI22_X1 U20157 ( .A1(n25235), .A2(n25453), .B1(n21267), .B2(n21002), .ZN(
        n6632) );
  OAI22_X1 U20158 ( .A1(n25235), .A2(n25456), .B1(n25225), .B2(n21001), .ZN(
        n6633) );
  OAI22_X1 U20159 ( .A1(n25235), .A2(n25459), .B1(n21267), .B2(n21000), .ZN(
        n6634) );
  OAI22_X1 U20160 ( .A1(n25235), .A2(n25462), .B1(n25225), .B2(n20999), .ZN(
        n6635) );
  OAI22_X1 U20161 ( .A1(n25236), .A2(n25465), .B1(n21267), .B2(n20998), .ZN(
        n6636) );
  OAI22_X1 U20162 ( .A1(n25236), .A2(n25468), .B1(n25225), .B2(n20997), .ZN(
        n6637) );
  OAI22_X1 U20163 ( .A1(n25236), .A2(n25471), .B1(n25226), .B2(n20996), .ZN(
        n6638) );
  OAI22_X1 U20164 ( .A1(n25236), .A2(n25474), .B1(n25227), .B2(n20995), .ZN(
        n6639) );
  OAI22_X1 U20165 ( .A1(n25236), .A2(n25477), .B1(n25225), .B2(n20994), .ZN(
        n6640) );
  OAI22_X1 U20166 ( .A1(n25237), .A2(n25480), .B1(n25225), .B2(n20993), .ZN(
        n6641) );
  OAI22_X1 U20167 ( .A1(n25237), .A2(n25483), .B1(n25226), .B2(n20992), .ZN(
        n6642) );
  OAI22_X1 U20168 ( .A1(n25237), .A2(n25486), .B1(n25227), .B2(n20991), .ZN(
        n6643) );
  OAI22_X1 U20169 ( .A1(n25237), .A2(n25489), .B1(n25225), .B2(n20990), .ZN(
        n6644) );
  OAI22_X1 U20170 ( .A1(n25237), .A2(n25492), .B1(n25225), .B2(n20989), .ZN(
        n6645) );
  OAI22_X1 U20171 ( .A1(n25238), .A2(n25495), .B1(n21267), .B2(n20988), .ZN(
        n6646) );
  OAI22_X1 U20172 ( .A1(n25238), .A2(n25498), .B1(n25225), .B2(n20987), .ZN(
        n6647) );
  OAI22_X1 U20173 ( .A1(n25238), .A2(n25501), .B1(n21267), .B2(n20986), .ZN(
        n6648) );
  OAI22_X1 U20174 ( .A1(n25238), .A2(n25504), .B1(n25225), .B2(n20985), .ZN(
        n6649) );
  OAI22_X1 U20175 ( .A1(n25238), .A2(n25507), .B1(n21267), .B2(n20984), .ZN(
        n6650) );
  OAI22_X1 U20176 ( .A1(n25239), .A2(n25510), .B1(n25225), .B2(n20983), .ZN(
        n6651) );
  OAI22_X1 U20177 ( .A1(n25239), .A2(n25513), .B1(n21267), .B2(n20982), .ZN(
        n6652) );
  OAI22_X1 U20178 ( .A1(n25239), .A2(n25516), .B1(n25225), .B2(n20981), .ZN(
        n6653) );
  OAI22_X1 U20179 ( .A1(n25239), .A2(n25519), .B1(n21267), .B2(n20980), .ZN(
        n6654) );
  OAI22_X1 U20180 ( .A1(n25239), .A2(n25522), .B1(n25225), .B2(n20979), .ZN(
        n6655) );
  OAI22_X1 U20181 ( .A1(n25215), .A2(n25417), .B1(n25209), .B2(n20978), .ZN(
        n6556) );
  OAI22_X1 U20182 ( .A1(n25216), .A2(n25420), .B1(n25210), .B2(n20977), .ZN(
        n6557) );
  OAI22_X1 U20183 ( .A1(n25216), .A2(n25423), .B1(n25208), .B2(n20976), .ZN(
        n6558) );
  OAI22_X1 U20184 ( .A1(n25216), .A2(n25426), .B1(n25209), .B2(n20975), .ZN(
        n6559) );
  OAI22_X1 U20185 ( .A1(n25216), .A2(n25429), .B1(n25210), .B2(n20974), .ZN(
        n6560) );
  OAI22_X1 U20186 ( .A1(n25216), .A2(n25432), .B1(n25208), .B2(n20973), .ZN(
        n6561) );
  OAI22_X1 U20187 ( .A1(n25217), .A2(n25435), .B1(n25209), .B2(n20972), .ZN(
        n6562) );
  OAI22_X1 U20188 ( .A1(n25217), .A2(n25438), .B1(n25210), .B2(n20971), .ZN(
        n6563) );
  OAI22_X1 U20189 ( .A1(n25217), .A2(n25441), .B1(n25208), .B2(n20970), .ZN(
        n6564) );
  OAI22_X1 U20190 ( .A1(n25217), .A2(n25444), .B1(n25209), .B2(n20969), .ZN(
        n6565) );
  OAI22_X1 U20191 ( .A1(n25217), .A2(n25447), .B1(n25210), .B2(n20968), .ZN(
        n6566) );
  OAI22_X1 U20192 ( .A1(n25218), .A2(n25450), .B1(n25208), .B2(n20967), .ZN(
        n6567) );
  OAI22_X1 U20193 ( .A1(n25218), .A2(n25453), .B1(n21270), .B2(n20966), .ZN(
        n6568) );
  OAI22_X1 U20194 ( .A1(n25218), .A2(n25456), .B1(n25208), .B2(n20965), .ZN(
        n6569) );
  OAI22_X1 U20195 ( .A1(n25218), .A2(n25459), .B1(n21270), .B2(n20964), .ZN(
        n6570) );
  OAI22_X1 U20196 ( .A1(n25218), .A2(n25462), .B1(n25208), .B2(n20963), .ZN(
        n6571) );
  OAI22_X1 U20197 ( .A1(n25219), .A2(n25465), .B1(n21270), .B2(n20962), .ZN(
        n6572) );
  OAI22_X1 U20198 ( .A1(n25219), .A2(n25468), .B1(n25208), .B2(n20961), .ZN(
        n6573) );
  OAI22_X1 U20199 ( .A1(n25219), .A2(n25471), .B1(n25209), .B2(n20960), .ZN(
        n6574) );
  OAI22_X1 U20200 ( .A1(n25219), .A2(n25474), .B1(n25210), .B2(n20959), .ZN(
        n6575) );
  OAI22_X1 U20201 ( .A1(n25219), .A2(n25477), .B1(n25208), .B2(n20958), .ZN(
        n6576) );
  OAI22_X1 U20202 ( .A1(n25220), .A2(n25480), .B1(n25208), .B2(n20957), .ZN(
        n6577) );
  OAI22_X1 U20203 ( .A1(n25220), .A2(n25483), .B1(n25209), .B2(n20956), .ZN(
        n6578) );
  OAI22_X1 U20204 ( .A1(n25220), .A2(n25486), .B1(n25210), .B2(n20955), .ZN(
        n6579) );
  OAI22_X1 U20205 ( .A1(n25220), .A2(n25489), .B1(n25208), .B2(n20954), .ZN(
        n6580) );
  OAI22_X1 U20206 ( .A1(n25220), .A2(n25492), .B1(n25208), .B2(n20953), .ZN(
        n6581) );
  OAI22_X1 U20207 ( .A1(n25221), .A2(n25495), .B1(n21270), .B2(n20952), .ZN(
        n6582) );
  OAI22_X1 U20208 ( .A1(n25221), .A2(n25498), .B1(n25208), .B2(n20951), .ZN(
        n6583) );
  OAI22_X1 U20209 ( .A1(n25221), .A2(n25501), .B1(n21270), .B2(n20950), .ZN(
        n6584) );
  OAI22_X1 U20210 ( .A1(n25221), .A2(n25504), .B1(n25208), .B2(n20949), .ZN(
        n6585) );
  OAI22_X1 U20211 ( .A1(n25221), .A2(n25507), .B1(n21270), .B2(n20948), .ZN(
        n6586) );
  OAI22_X1 U20212 ( .A1(n25222), .A2(n25510), .B1(n25208), .B2(n20947), .ZN(
        n6587) );
  OAI22_X1 U20213 ( .A1(n25222), .A2(n25513), .B1(n21270), .B2(n20946), .ZN(
        n6588) );
  OAI22_X1 U20214 ( .A1(n25222), .A2(n25516), .B1(n25208), .B2(n20945), .ZN(
        n6589) );
  OAI22_X1 U20215 ( .A1(n25222), .A2(n25519), .B1(n21270), .B2(n20944), .ZN(
        n6590) );
  OAI22_X1 U20216 ( .A1(n25222), .A2(n25522), .B1(n25208), .B2(n20943), .ZN(
        n6591) );
  OAI22_X1 U20217 ( .A1(n25147), .A2(n25418), .B1(n25141), .B2(n20942), .ZN(
        n6300) );
  OAI22_X1 U20218 ( .A1(n25148), .A2(n25421), .B1(n25142), .B2(n20941), .ZN(
        n6301) );
  OAI22_X1 U20219 ( .A1(n25148), .A2(n25424), .B1(n25140), .B2(n20940), .ZN(
        n6302) );
  OAI22_X1 U20220 ( .A1(n25148), .A2(n25427), .B1(n25141), .B2(n20939), .ZN(
        n6303) );
  OAI22_X1 U20221 ( .A1(n25148), .A2(n25430), .B1(n25142), .B2(n20938), .ZN(
        n6304) );
  OAI22_X1 U20222 ( .A1(n25148), .A2(n25433), .B1(n25140), .B2(n20937), .ZN(
        n6305) );
  OAI22_X1 U20223 ( .A1(n25149), .A2(n25436), .B1(n25141), .B2(n20936), .ZN(
        n6306) );
  OAI22_X1 U20224 ( .A1(n25149), .A2(n25439), .B1(n25142), .B2(n20935), .ZN(
        n6307) );
  OAI22_X1 U20225 ( .A1(n25149), .A2(n25442), .B1(n25140), .B2(n20934), .ZN(
        n6308) );
  OAI22_X1 U20226 ( .A1(n25149), .A2(n25445), .B1(n25141), .B2(n20933), .ZN(
        n6309) );
  OAI22_X1 U20227 ( .A1(n25149), .A2(n25448), .B1(n25142), .B2(n20932), .ZN(
        n6310) );
  OAI22_X1 U20228 ( .A1(n25150), .A2(n25451), .B1(n25140), .B2(n20931), .ZN(
        n6311) );
  OAI22_X1 U20229 ( .A1(n25150), .A2(n25454), .B1(n21275), .B2(n20930), .ZN(
        n6312) );
  OAI22_X1 U20230 ( .A1(n25150), .A2(n25457), .B1(n25140), .B2(n20929), .ZN(
        n6313) );
  OAI22_X1 U20231 ( .A1(n25150), .A2(n25460), .B1(n21275), .B2(n20928), .ZN(
        n6314) );
  OAI22_X1 U20232 ( .A1(n25150), .A2(n25463), .B1(n25140), .B2(n20927), .ZN(
        n6315) );
  OAI22_X1 U20233 ( .A1(n25151), .A2(n25466), .B1(n21275), .B2(n20926), .ZN(
        n6316) );
  OAI22_X1 U20234 ( .A1(n25151), .A2(n25469), .B1(n25140), .B2(n20925), .ZN(
        n6317) );
  OAI22_X1 U20235 ( .A1(n25151), .A2(n25472), .B1(n25141), .B2(n20924), .ZN(
        n6318) );
  OAI22_X1 U20236 ( .A1(n25151), .A2(n25475), .B1(n25142), .B2(n20923), .ZN(
        n6319) );
  OAI22_X1 U20237 ( .A1(n25151), .A2(n25478), .B1(n25140), .B2(n20922), .ZN(
        n6320) );
  OAI22_X1 U20238 ( .A1(n25152), .A2(n25481), .B1(n25140), .B2(n20921), .ZN(
        n6321) );
  OAI22_X1 U20239 ( .A1(n25152), .A2(n25484), .B1(n25141), .B2(n20920), .ZN(
        n6322) );
  OAI22_X1 U20240 ( .A1(n25152), .A2(n25487), .B1(n25142), .B2(n20919), .ZN(
        n6323) );
  OAI22_X1 U20241 ( .A1(n25152), .A2(n25490), .B1(n25140), .B2(n20918), .ZN(
        n6324) );
  OAI22_X1 U20242 ( .A1(n25152), .A2(n25493), .B1(n25140), .B2(n20917), .ZN(
        n6325) );
  OAI22_X1 U20243 ( .A1(n25153), .A2(n25496), .B1(n21275), .B2(n20916), .ZN(
        n6326) );
  OAI22_X1 U20244 ( .A1(n25153), .A2(n25499), .B1(n25140), .B2(n20915), .ZN(
        n6327) );
  OAI22_X1 U20245 ( .A1(n25153), .A2(n25502), .B1(n21275), .B2(n20914), .ZN(
        n6328) );
  OAI22_X1 U20246 ( .A1(n25153), .A2(n25505), .B1(n25140), .B2(n20913), .ZN(
        n6329) );
  OAI22_X1 U20247 ( .A1(n25153), .A2(n25508), .B1(n21275), .B2(n20912), .ZN(
        n6330) );
  OAI22_X1 U20248 ( .A1(n25154), .A2(n25511), .B1(n25140), .B2(n20911), .ZN(
        n6331) );
  OAI22_X1 U20249 ( .A1(n25154), .A2(n25514), .B1(n21275), .B2(n20910), .ZN(
        n6332) );
  OAI22_X1 U20250 ( .A1(n25154), .A2(n25517), .B1(n25140), .B2(n20909), .ZN(
        n6333) );
  OAI22_X1 U20251 ( .A1(n25154), .A2(n25520), .B1(n21275), .B2(n20908), .ZN(
        n6334) );
  OAI22_X1 U20252 ( .A1(n25154), .A2(n25523), .B1(n25140), .B2(n20907), .ZN(
        n6335) );
  OAI22_X1 U20253 ( .A1(n25249), .A2(n25417), .B1(n25243), .B2(n20726), .ZN(
        n6684) );
  OAI22_X1 U20254 ( .A1(n25250), .A2(n25420), .B1(n25244), .B2(n20725), .ZN(
        n6685) );
  OAI22_X1 U20255 ( .A1(n25250), .A2(n25423), .B1(n25242), .B2(n20724), .ZN(
        n6686) );
  OAI22_X1 U20256 ( .A1(n25250), .A2(n25426), .B1(n25243), .B2(n20723), .ZN(
        n6687) );
  OAI22_X1 U20257 ( .A1(n25250), .A2(n25429), .B1(n25244), .B2(n20722), .ZN(
        n6688) );
  OAI22_X1 U20258 ( .A1(n25250), .A2(n25432), .B1(n25242), .B2(n20721), .ZN(
        n6689) );
  OAI22_X1 U20259 ( .A1(n25251), .A2(n25435), .B1(n25243), .B2(n20720), .ZN(
        n6690) );
  OAI22_X1 U20260 ( .A1(n25251), .A2(n25438), .B1(n25244), .B2(n20719), .ZN(
        n6691) );
  OAI22_X1 U20261 ( .A1(n25251), .A2(n25441), .B1(n25242), .B2(n20718), .ZN(
        n6692) );
  OAI22_X1 U20262 ( .A1(n25251), .A2(n25444), .B1(n25243), .B2(n20717), .ZN(
        n6693) );
  OAI22_X1 U20263 ( .A1(n25251), .A2(n25447), .B1(n25244), .B2(n20716), .ZN(
        n6694) );
  OAI22_X1 U20264 ( .A1(n25252), .A2(n25450), .B1(n25242), .B2(n20715), .ZN(
        n6695) );
  OAI22_X1 U20265 ( .A1(n25252), .A2(n25453), .B1(n21265), .B2(n20714), .ZN(
        n6696) );
  OAI22_X1 U20266 ( .A1(n25252), .A2(n25456), .B1(n25242), .B2(n20713), .ZN(
        n6697) );
  OAI22_X1 U20267 ( .A1(n25252), .A2(n25459), .B1(n21265), .B2(n20712), .ZN(
        n6698) );
  OAI22_X1 U20268 ( .A1(n25252), .A2(n25462), .B1(n25242), .B2(n20711), .ZN(
        n6699) );
  OAI22_X1 U20269 ( .A1(n25253), .A2(n25465), .B1(n21265), .B2(n20710), .ZN(
        n6700) );
  OAI22_X1 U20270 ( .A1(n25253), .A2(n25468), .B1(n25242), .B2(n20709), .ZN(
        n6701) );
  OAI22_X1 U20271 ( .A1(n25253), .A2(n25471), .B1(n25243), .B2(n20708), .ZN(
        n6702) );
  OAI22_X1 U20272 ( .A1(n25253), .A2(n25474), .B1(n25244), .B2(n20707), .ZN(
        n6703) );
  OAI22_X1 U20273 ( .A1(n25253), .A2(n25477), .B1(n25242), .B2(n20706), .ZN(
        n6704) );
  OAI22_X1 U20274 ( .A1(n25254), .A2(n25480), .B1(n25242), .B2(n20705), .ZN(
        n6705) );
  OAI22_X1 U20275 ( .A1(n25254), .A2(n25483), .B1(n25243), .B2(n20704), .ZN(
        n6706) );
  OAI22_X1 U20276 ( .A1(n25254), .A2(n25486), .B1(n25244), .B2(n20703), .ZN(
        n6707) );
  OAI22_X1 U20277 ( .A1(n25254), .A2(n25489), .B1(n25242), .B2(n20702), .ZN(
        n6708) );
  OAI22_X1 U20278 ( .A1(n25254), .A2(n25492), .B1(n25242), .B2(n20701), .ZN(
        n6709) );
  OAI22_X1 U20279 ( .A1(n25255), .A2(n25495), .B1(n21265), .B2(n20700), .ZN(
        n6710) );
  OAI22_X1 U20280 ( .A1(n25255), .A2(n25498), .B1(n25242), .B2(n20699), .ZN(
        n6711) );
  OAI22_X1 U20281 ( .A1(n25255), .A2(n25501), .B1(n21265), .B2(n20698), .ZN(
        n6712) );
  OAI22_X1 U20282 ( .A1(n25255), .A2(n25504), .B1(n25242), .B2(n20697), .ZN(
        n6713) );
  OAI22_X1 U20283 ( .A1(n25255), .A2(n25507), .B1(n21265), .B2(n20696), .ZN(
        n6714) );
  OAI22_X1 U20284 ( .A1(n25256), .A2(n25510), .B1(n25242), .B2(n20695), .ZN(
        n6715) );
  OAI22_X1 U20285 ( .A1(n25256), .A2(n25513), .B1(n21265), .B2(n20694), .ZN(
        n6716) );
  OAI22_X1 U20286 ( .A1(n25256), .A2(n25516), .B1(n25242), .B2(n20693), .ZN(
        n6717) );
  OAI22_X1 U20287 ( .A1(n25256), .A2(n25519), .B1(n21265), .B2(n20692), .ZN(
        n6718) );
  OAI22_X1 U20288 ( .A1(n25256), .A2(n25522), .B1(n25242), .B2(n20691), .ZN(
        n6719) );
  OAI22_X1 U20289 ( .A1(n25079), .A2(n25418), .B1(n25073), .B2(n20690), .ZN(
        n6044) );
  OAI22_X1 U20290 ( .A1(n25080), .A2(n25421), .B1(n25074), .B2(n20689), .ZN(
        n6045) );
  OAI22_X1 U20291 ( .A1(n25080), .A2(n25424), .B1(n25072), .B2(n20688), .ZN(
        n6046) );
  OAI22_X1 U20292 ( .A1(n25080), .A2(n25427), .B1(n25073), .B2(n20687), .ZN(
        n6047) );
  OAI22_X1 U20293 ( .A1(n25080), .A2(n25430), .B1(n25074), .B2(n20686), .ZN(
        n6048) );
  OAI22_X1 U20294 ( .A1(n25080), .A2(n25433), .B1(n25072), .B2(n20685), .ZN(
        n6049) );
  OAI22_X1 U20295 ( .A1(n25081), .A2(n25436), .B1(n25073), .B2(n20684), .ZN(
        n6050) );
  OAI22_X1 U20296 ( .A1(n25081), .A2(n25439), .B1(n25074), .B2(n20683), .ZN(
        n6051) );
  OAI22_X1 U20297 ( .A1(n25081), .A2(n25442), .B1(n25072), .B2(n20682), .ZN(
        n6052) );
  OAI22_X1 U20298 ( .A1(n25081), .A2(n25445), .B1(n25073), .B2(n20681), .ZN(
        n6053) );
  OAI22_X1 U20299 ( .A1(n25081), .A2(n25448), .B1(n25074), .B2(n20680), .ZN(
        n6054) );
  OAI22_X1 U20300 ( .A1(n25082), .A2(n25451), .B1(n25072), .B2(n20679), .ZN(
        n6055) );
  OAI22_X1 U20301 ( .A1(n25082), .A2(n25454), .B1(n21279), .B2(n20678), .ZN(
        n6056) );
  OAI22_X1 U20302 ( .A1(n25082), .A2(n25457), .B1(n25072), .B2(n20677), .ZN(
        n6057) );
  OAI22_X1 U20303 ( .A1(n25082), .A2(n25460), .B1(n21279), .B2(n20676), .ZN(
        n6058) );
  OAI22_X1 U20304 ( .A1(n25082), .A2(n25463), .B1(n25072), .B2(n20675), .ZN(
        n6059) );
  OAI22_X1 U20305 ( .A1(n25083), .A2(n25466), .B1(n21279), .B2(n20674), .ZN(
        n6060) );
  OAI22_X1 U20306 ( .A1(n25083), .A2(n25469), .B1(n25072), .B2(n20673), .ZN(
        n6061) );
  OAI22_X1 U20307 ( .A1(n25083), .A2(n25472), .B1(n25073), .B2(n20672), .ZN(
        n6062) );
  OAI22_X1 U20308 ( .A1(n25083), .A2(n25475), .B1(n25074), .B2(n20671), .ZN(
        n6063) );
  OAI22_X1 U20309 ( .A1(n25083), .A2(n25478), .B1(n25072), .B2(n20670), .ZN(
        n6064) );
  OAI22_X1 U20310 ( .A1(n25084), .A2(n25481), .B1(n25072), .B2(n20669), .ZN(
        n6065) );
  OAI22_X1 U20311 ( .A1(n25084), .A2(n25484), .B1(n25073), .B2(n20668), .ZN(
        n6066) );
  OAI22_X1 U20312 ( .A1(n25084), .A2(n25487), .B1(n25074), .B2(n20667), .ZN(
        n6067) );
  OAI22_X1 U20313 ( .A1(n25084), .A2(n25490), .B1(n25072), .B2(n20666), .ZN(
        n6068) );
  OAI22_X1 U20314 ( .A1(n25084), .A2(n25493), .B1(n25072), .B2(n20665), .ZN(
        n6069) );
  OAI22_X1 U20315 ( .A1(n25085), .A2(n25496), .B1(n21279), .B2(n20664), .ZN(
        n6070) );
  OAI22_X1 U20316 ( .A1(n25085), .A2(n25499), .B1(n25072), .B2(n20663), .ZN(
        n6071) );
  OAI22_X1 U20317 ( .A1(n25085), .A2(n25502), .B1(n21279), .B2(n20662), .ZN(
        n6072) );
  OAI22_X1 U20318 ( .A1(n25085), .A2(n25505), .B1(n25072), .B2(n20661), .ZN(
        n6073) );
  OAI22_X1 U20319 ( .A1(n25085), .A2(n25508), .B1(n21279), .B2(n20660), .ZN(
        n6074) );
  OAI22_X1 U20320 ( .A1(n25086), .A2(n25511), .B1(n25072), .B2(n20659), .ZN(
        n6075) );
  OAI22_X1 U20321 ( .A1(n25086), .A2(n25514), .B1(n21279), .B2(n20658), .ZN(
        n6076) );
  OAI22_X1 U20322 ( .A1(n25086), .A2(n25517), .B1(n25072), .B2(n20657), .ZN(
        n6077) );
  OAI22_X1 U20323 ( .A1(n25086), .A2(n25520), .B1(n21279), .B2(n20656), .ZN(
        n6078) );
  OAI22_X1 U20324 ( .A1(n25086), .A2(n25523), .B1(n25072), .B2(n20655), .ZN(
        n6079) );
  OAI22_X1 U20325 ( .A1(n25011), .A2(n25418), .B1(n25005), .B2(n20654), .ZN(
        n5788) );
  OAI22_X1 U20326 ( .A1(n25012), .A2(n25421), .B1(n25006), .B2(n20653), .ZN(
        n5789) );
  OAI22_X1 U20327 ( .A1(n25012), .A2(n25424), .B1(n25004), .B2(n20652), .ZN(
        n5790) );
  OAI22_X1 U20328 ( .A1(n25012), .A2(n25427), .B1(n25005), .B2(n20651), .ZN(
        n5791) );
  OAI22_X1 U20329 ( .A1(n25012), .A2(n25430), .B1(n25006), .B2(n20650), .ZN(
        n5792) );
  OAI22_X1 U20330 ( .A1(n25012), .A2(n25433), .B1(n25004), .B2(n20649), .ZN(
        n5793) );
  OAI22_X1 U20331 ( .A1(n25013), .A2(n25436), .B1(n25005), .B2(n20648), .ZN(
        n5794) );
  OAI22_X1 U20332 ( .A1(n25013), .A2(n25439), .B1(n25006), .B2(n20647), .ZN(
        n5795) );
  OAI22_X1 U20333 ( .A1(n25013), .A2(n25442), .B1(n25004), .B2(n20646), .ZN(
        n5796) );
  OAI22_X1 U20334 ( .A1(n25013), .A2(n25445), .B1(n25005), .B2(n20645), .ZN(
        n5797) );
  OAI22_X1 U20335 ( .A1(n25013), .A2(n25448), .B1(n25006), .B2(n20644), .ZN(
        n5798) );
  OAI22_X1 U20336 ( .A1(n25014), .A2(n25451), .B1(n25004), .B2(n20643), .ZN(
        n5799) );
  OAI22_X1 U20337 ( .A1(n25014), .A2(n25454), .B1(n21284), .B2(n20642), .ZN(
        n5800) );
  OAI22_X1 U20338 ( .A1(n25014), .A2(n25457), .B1(n25004), .B2(n20641), .ZN(
        n5801) );
  OAI22_X1 U20339 ( .A1(n25014), .A2(n25460), .B1(n21284), .B2(n20640), .ZN(
        n5802) );
  OAI22_X1 U20340 ( .A1(n25014), .A2(n25463), .B1(n25004), .B2(n20639), .ZN(
        n5803) );
  OAI22_X1 U20341 ( .A1(n25015), .A2(n25466), .B1(n21284), .B2(n20638), .ZN(
        n5804) );
  OAI22_X1 U20342 ( .A1(n25015), .A2(n25469), .B1(n25004), .B2(n20637), .ZN(
        n5805) );
  OAI22_X1 U20343 ( .A1(n25015), .A2(n25472), .B1(n25005), .B2(n20636), .ZN(
        n5806) );
  OAI22_X1 U20344 ( .A1(n25015), .A2(n25475), .B1(n25006), .B2(n20635), .ZN(
        n5807) );
  OAI22_X1 U20345 ( .A1(n25015), .A2(n25478), .B1(n25004), .B2(n20634), .ZN(
        n5808) );
  OAI22_X1 U20346 ( .A1(n25016), .A2(n25481), .B1(n25004), .B2(n20633), .ZN(
        n5809) );
  OAI22_X1 U20347 ( .A1(n25016), .A2(n25484), .B1(n25005), .B2(n20632), .ZN(
        n5810) );
  OAI22_X1 U20348 ( .A1(n25016), .A2(n25487), .B1(n25006), .B2(n20631), .ZN(
        n5811) );
  OAI22_X1 U20349 ( .A1(n25016), .A2(n25490), .B1(n25004), .B2(n20630), .ZN(
        n5812) );
  OAI22_X1 U20350 ( .A1(n25016), .A2(n25493), .B1(n25004), .B2(n20629), .ZN(
        n5813) );
  OAI22_X1 U20351 ( .A1(n25017), .A2(n25496), .B1(n21284), .B2(n20628), .ZN(
        n5814) );
  OAI22_X1 U20352 ( .A1(n25017), .A2(n25499), .B1(n25004), .B2(n20627), .ZN(
        n5815) );
  OAI22_X1 U20353 ( .A1(n25017), .A2(n25502), .B1(n21284), .B2(n20626), .ZN(
        n5816) );
  OAI22_X1 U20354 ( .A1(n25017), .A2(n25505), .B1(n25004), .B2(n20625), .ZN(
        n5817) );
  OAI22_X1 U20355 ( .A1(n25017), .A2(n25508), .B1(n21284), .B2(n20624), .ZN(
        n5818) );
  OAI22_X1 U20356 ( .A1(n25018), .A2(n25511), .B1(n25004), .B2(n20623), .ZN(
        n5819) );
  OAI22_X1 U20357 ( .A1(n25018), .A2(n25514), .B1(n21284), .B2(n20622), .ZN(
        n5820) );
  OAI22_X1 U20358 ( .A1(n25018), .A2(n25517), .B1(n25004), .B2(n20621), .ZN(
        n5821) );
  OAI22_X1 U20359 ( .A1(n25018), .A2(n25520), .B1(n21284), .B2(n20620), .ZN(
        n5822) );
  OAI22_X1 U20360 ( .A1(n25018), .A2(n25523), .B1(n25004), .B2(n20619), .ZN(
        n5823) );
  OAI22_X1 U20361 ( .A1(n24909), .A2(n25419), .B1(n24903), .B2(n20618), .ZN(
        n5404) );
  OAI22_X1 U20362 ( .A1(n24910), .A2(n25422), .B1(n24904), .B2(n20617), .ZN(
        n5405) );
  OAI22_X1 U20363 ( .A1(n24910), .A2(n25425), .B1(n24902), .B2(n20616), .ZN(
        n5406) );
  OAI22_X1 U20364 ( .A1(n24910), .A2(n25428), .B1(n24903), .B2(n20615), .ZN(
        n5407) );
  OAI22_X1 U20365 ( .A1(n24910), .A2(n25431), .B1(n24904), .B2(n20614), .ZN(
        n5408) );
  OAI22_X1 U20366 ( .A1(n24910), .A2(n25434), .B1(n24902), .B2(n20613), .ZN(
        n5409) );
  OAI22_X1 U20367 ( .A1(n24911), .A2(n25437), .B1(n24903), .B2(n20612), .ZN(
        n5410) );
  OAI22_X1 U20368 ( .A1(n24911), .A2(n25440), .B1(n24904), .B2(n20611), .ZN(
        n5411) );
  OAI22_X1 U20369 ( .A1(n24911), .A2(n25443), .B1(n24902), .B2(n20610), .ZN(
        n5412) );
  OAI22_X1 U20370 ( .A1(n24911), .A2(n25446), .B1(n24903), .B2(n20609), .ZN(
        n5413) );
  OAI22_X1 U20371 ( .A1(n24911), .A2(n25449), .B1(n24904), .B2(n20608), .ZN(
        n5414) );
  OAI22_X1 U20372 ( .A1(n24912), .A2(n25452), .B1(n24902), .B2(n20607), .ZN(
        n5415) );
  OAI22_X1 U20373 ( .A1(n24912), .A2(n25455), .B1(n21291), .B2(n20606), .ZN(
        n5416) );
  OAI22_X1 U20374 ( .A1(n24912), .A2(n25458), .B1(n24902), .B2(n20605), .ZN(
        n5417) );
  OAI22_X1 U20375 ( .A1(n24912), .A2(n25461), .B1(n21291), .B2(n20604), .ZN(
        n5418) );
  OAI22_X1 U20376 ( .A1(n24912), .A2(n25464), .B1(n24902), .B2(n20603), .ZN(
        n5419) );
  OAI22_X1 U20377 ( .A1(n24913), .A2(n25467), .B1(n21291), .B2(n20602), .ZN(
        n5420) );
  OAI22_X1 U20378 ( .A1(n24913), .A2(n25470), .B1(n24902), .B2(n20601), .ZN(
        n5421) );
  OAI22_X1 U20379 ( .A1(n24913), .A2(n25473), .B1(n24903), .B2(n20600), .ZN(
        n5422) );
  OAI22_X1 U20380 ( .A1(n24913), .A2(n25476), .B1(n24904), .B2(n20599), .ZN(
        n5423) );
  OAI22_X1 U20381 ( .A1(n24913), .A2(n25479), .B1(n24902), .B2(n20598), .ZN(
        n5424) );
  OAI22_X1 U20382 ( .A1(n24914), .A2(n25482), .B1(n24902), .B2(n20597), .ZN(
        n5425) );
  OAI22_X1 U20383 ( .A1(n24914), .A2(n25485), .B1(n24903), .B2(n20596), .ZN(
        n5426) );
  OAI22_X1 U20384 ( .A1(n24914), .A2(n25488), .B1(n24904), .B2(n20595), .ZN(
        n5427) );
  OAI22_X1 U20385 ( .A1(n24914), .A2(n25491), .B1(n24902), .B2(n20594), .ZN(
        n5428) );
  OAI22_X1 U20386 ( .A1(n24914), .A2(n25494), .B1(n24902), .B2(n20593), .ZN(
        n5429) );
  OAI22_X1 U20387 ( .A1(n24915), .A2(n25497), .B1(n21291), .B2(n20592), .ZN(
        n5430) );
  OAI22_X1 U20388 ( .A1(n24915), .A2(n25500), .B1(n24902), .B2(n20591), .ZN(
        n5431) );
  OAI22_X1 U20389 ( .A1(n24915), .A2(n25503), .B1(n21291), .B2(n20590), .ZN(
        n5432) );
  OAI22_X1 U20390 ( .A1(n24915), .A2(n25506), .B1(n24902), .B2(n20589), .ZN(
        n5433) );
  OAI22_X1 U20391 ( .A1(n24915), .A2(n25509), .B1(n21291), .B2(n20588), .ZN(
        n5434) );
  OAI22_X1 U20392 ( .A1(n24916), .A2(n25512), .B1(n24902), .B2(n20587), .ZN(
        n5435) );
  OAI22_X1 U20393 ( .A1(n24916), .A2(n25515), .B1(n21291), .B2(n20586), .ZN(
        n5436) );
  OAI22_X1 U20394 ( .A1(n24916), .A2(n25518), .B1(n24902), .B2(n20585), .ZN(
        n5437) );
  OAI22_X1 U20395 ( .A1(n24916), .A2(n25521), .B1(n21291), .B2(n20584), .ZN(
        n5438) );
  OAI22_X1 U20396 ( .A1(n24916), .A2(n25524), .B1(n24902), .B2(n20583), .ZN(
        n5439) );
  OAI22_X1 U20397 ( .A1(n24841), .A2(n25419), .B1(n24835), .B2(n20582), .ZN(
        n5148) );
  OAI22_X1 U20398 ( .A1(n24842), .A2(n25422), .B1(n24836), .B2(n20581), .ZN(
        n5149) );
  OAI22_X1 U20399 ( .A1(n24842), .A2(n25425), .B1(n24834), .B2(n20580), .ZN(
        n5150) );
  OAI22_X1 U20400 ( .A1(n24842), .A2(n25428), .B1(n24835), .B2(n20579), .ZN(
        n5151) );
  OAI22_X1 U20401 ( .A1(n24842), .A2(n25431), .B1(n24836), .B2(n20578), .ZN(
        n5152) );
  OAI22_X1 U20402 ( .A1(n24842), .A2(n25434), .B1(n24834), .B2(n20577), .ZN(
        n5153) );
  OAI22_X1 U20403 ( .A1(n24843), .A2(n25437), .B1(n24835), .B2(n20576), .ZN(
        n5154) );
  OAI22_X1 U20404 ( .A1(n24843), .A2(n25440), .B1(n24836), .B2(n20575), .ZN(
        n5155) );
  OAI22_X1 U20405 ( .A1(n24843), .A2(n25443), .B1(n24834), .B2(n20574), .ZN(
        n5156) );
  OAI22_X1 U20406 ( .A1(n24843), .A2(n25446), .B1(n24835), .B2(n20573), .ZN(
        n5157) );
  OAI22_X1 U20407 ( .A1(n24843), .A2(n25449), .B1(n24836), .B2(n20572), .ZN(
        n5158) );
  OAI22_X1 U20408 ( .A1(n24844), .A2(n25452), .B1(n24834), .B2(n20571), .ZN(
        n5159) );
  OAI22_X1 U20409 ( .A1(n24844), .A2(n25455), .B1(n21295), .B2(n20570), .ZN(
        n5160) );
  OAI22_X1 U20410 ( .A1(n24844), .A2(n25458), .B1(n24834), .B2(n20569), .ZN(
        n5161) );
  OAI22_X1 U20411 ( .A1(n24844), .A2(n25461), .B1(n21295), .B2(n20568), .ZN(
        n5162) );
  OAI22_X1 U20412 ( .A1(n24844), .A2(n25464), .B1(n24834), .B2(n20567), .ZN(
        n5163) );
  OAI22_X1 U20413 ( .A1(n24845), .A2(n25467), .B1(n21295), .B2(n20566), .ZN(
        n5164) );
  OAI22_X1 U20414 ( .A1(n24845), .A2(n25470), .B1(n24834), .B2(n20565), .ZN(
        n5165) );
  OAI22_X1 U20415 ( .A1(n24845), .A2(n25473), .B1(n24835), .B2(n20564), .ZN(
        n5166) );
  OAI22_X1 U20416 ( .A1(n24845), .A2(n25476), .B1(n24836), .B2(n20563), .ZN(
        n5167) );
  OAI22_X1 U20417 ( .A1(n24845), .A2(n25479), .B1(n24834), .B2(n20562), .ZN(
        n5168) );
  OAI22_X1 U20418 ( .A1(n24846), .A2(n25482), .B1(n24834), .B2(n20561), .ZN(
        n5169) );
  OAI22_X1 U20419 ( .A1(n24846), .A2(n25485), .B1(n24835), .B2(n20560), .ZN(
        n5170) );
  OAI22_X1 U20420 ( .A1(n24846), .A2(n25488), .B1(n24836), .B2(n20559), .ZN(
        n5171) );
  OAI22_X1 U20421 ( .A1(n24846), .A2(n25491), .B1(n24834), .B2(n20558), .ZN(
        n5172) );
  OAI22_X1 U20422 ( .A1(n24846), .A2(n25494), .B1(n24834), .B2(n20557), .ZN(
        n5173) );
  OAI22_X1 U20423 ( .A1(n24847), .A2(n25497), .B1(n21295), .B2(n20556), .ZN(
        n5174) );
  OAI22_X1 U20424 ( .A1(n24847), .A2(n25500), .B1(n24834), .B2(n20555), .ZN(
        n5175) );
  OAI22_X1 U20425 ( .A1(n24847), .A2(n25503), .B1(n21295), .B2(n20554), .ZN(
        n5176) );
  OAI22_X1 U20426 ( .A1(n24847), .A2(n25506), .B1(n24834), .B2(n20553), .ZN(
        n5177) );
  OAI22_X1 U20427 ( .A1(n24847), .A2(n25509), .B1(n21295), .B2(n20552), .ZN(
        n5178) );
  OAI22_X1 U20428 ( .A1(n24848), .A2(n25512), .B1(n24834), .B2(n20551), .ZN(
        n5179) );
  OAI22_X1 U20429 ( .A1(n24848), .A2(n25515), .B1(n21295), .B2(n20550), .ZN(
        n5180) );
  OAI22_X1 U20430 ( .A1(n24848), .A2(n25518), .B1(n24834), .B2(n20549), .ZN(
        n5181) );
  OAI22_X1 U20431 ( .A1(n24848), .A2(n25521), .B1(n21295), .B2(n20548), .ZN(
        n5182) );
  OAI22_X1 U20432 ( .A1(n24848), .A2(n25524), .B1(n24834), .B2(n20547), .ZN(
        n5183) );
  OAI22_X1 U20433 ( .A1(n25062), .A2(n25418), .B1(n25056), .B2(n20481), .ZN(
        n5980) );
  OAI22_X1 U20434 ( .A1(n25063), .A2(n25421), .B1(n25057), .B2(n20480), .ZN(
        n5981) );
  OAI22_X1 U20435 ( .A1(n25063), .A2(n25424), .B1(n25055), .B2(n20479), .ZN(
        n5982) );
  OAI22_X1 U20436 ( .A1(n25063), .A2(n25427), .B1(n25056), .B2(n20478), .ZN(
        n5983) );
  OAI22_X1 U20437 ( .A1(n25063), .A2(n25430), .B1(n25057), .B2(n20477), .ZN(
        n5984) );
  OAI22_X1 U20438 ( .A1(n25063), .A2(n25433), .B1(n25055), .B2(n20476), .ZN(
        n5985) );
  OAI22_X1 U20439 ( .A1(n25064), .A2(n25436), .B1(n25056), .B2(n20475), .ZN(
        n5986) );
  OAI22_X1 U20440 ( .A1(n25064), .A2(n25439), .B1(n25057), .B2(n20474), .ZN(
        n5987) );
  OAI22_X1 U20441 ( .A1(n25064), .A2(n25442), .B1(n25055), .B2(n20473), .ZN(
        n5988) );
  OAI22_X1 U20442 ( .A1(n25064), .A2(n25445), .B1(n25056), .B2(n20472), .ZN(
        n5989) );
  OAI22_X1 U20443 ( .A1(n25064), .A2(n25448), .B1(n25057), .B2(n20471), .ZN(
        n5990) );
  OAI22_X1 U20444 ( .A1(n25065), .A2(n25451), .B1(n25055), .B2(n20470), .ZN(
        n5991) );
  OAI22_X1 U20445 ( .A1(n25065), .A2(n25454), .B1(n21281), .B2(n20469), .ZN(
        n5992) );
  OAI22_X1 U20446 ( .A1(n25065), .A2(n25457), .B1(n25055), .B2(n20468), .ZN(
        n5993) );
  OAI22_X1 U20447 ( .A1(n25065), .A2(n25460), .B1(n21281), .B2(n20467), .ZN(
        n5994) );
  OAI22_X1 U20448 ( .A1(n25065), .A2(n25463), .B1(n25055), .B2(n20466), .ZN(
        n5995) );
  OAI22_X1 U20449 ( .A1(n25066), .A2(n25466), .B1(n21281), .B2(n20465), .ZN(
        n5996) );
  OAI22_X1 U20450 ( .A1(n25066), .A2(n25469), .B1(n25055), .B2(n20464), .ZN(
        n5997) );
  OAI22_X1 U20451 ( .A1(n25066), .A2(n25472), .B1(n25056), .B2(n20463), .ZN(
        n5998) );
  OAI22_X1 U20452 ( .A1(n25066), .A2(n25475), .B1(n25057), .B2(n20462), .ZN(
        n5999) );
  OAI22_X1 U20453 ( .A1(n25066), .A2(n25478), .B1(n25055), .B2(n20461), .ZN(
        n6000) );
  OAI22_X1 U20454 ( .A1(n25067), .A2(n25481), .B1(n25055), .B2(n20460), .ZN(
        n6001) );
  OAI22_X1 U20455 ( .A1(n25067), .A2(n25484), .B1(n25056), .B2(n20459), .ZN(
        n6002) );
  OAI22_X1 U20456 ( .A1(n25067), .A2(n25487), .B1(n25057), .B2(n20458), .ZN(
        n6003) );
  OAI22_X1 U20457 ( .A1(n25067), .A2(n25490), .B1(n25055), .B2(n20457), .ZN(
        n6004) );
  OAI22_X1 U20458 ( .A1(n25067), .A2(n25493), .B1(n25055), .B2(n20456), .ZN(
        n6005) );
  OAI22_X1 U20459 ( .A1(n25068), .A2(n25496), .B1(n21281), .B2(n20455), .ZN(
        n6006) );
  OAI22_X1 U20460 ( .A1(n25068), .A2(n25499), .B1(n25055), .B2(n20454), .ZN(
        n6007) );
  OAI22_X1 U20461 ( .A1(n25068), .A2(n25502), .B1(n21281), .B2(n20453), .ZN(
        n6008) );
  OAI22_X1 U20462 ( .A1(n25068), .A2(n25505), .B1(n25055), .B2(n20452), .ZN(
        n6009) );
  OAI22_X1 U20463 ( .A1(n25068), .A2(n25508), .B1(n21281), .B2(n20451), .ZN(
        n6010) );
  OAI22_X1 U20464 ( .A1(n25069), .A2(n25511), .B1(n25055), .B2(n20450), .ZN(
        n6011) );
  OAI22_X1 U20465 ( .A1(n25069), .A2(n25514), .B1(n21281), .B2(n20449), .ZN(
        n6012) );
  OAI22_X1 U20466 ( .A1(n25069), .A2(n25517), .B1(n25055), .B2(n20448), .ZN(
        n6013) );
  OAI22_X1 U20467 ( .A1(n25069), .A2(n25520), .B1(n21281), .B2(n20447), .ZN(
        n6014) );
  OAI22_X1 U20468 ( .A1(n25069), .A2(n25523), .B1(n25055), .B2(n20446), .ZN(
        n6015) );
  OAI22_X1 U20469 ( .A1(n25317), .A2(n25417), .B1(n25311), .B2(n20373), .ZN(
        n6940) );
  OAI22_X1 U20470 ( .A1(n25318), .A2(n25420), .B1(n25312), .B2(n20372), .ZN(
        n6941) );
  OAI22_X1 U20471 ( .A1(n25318), .A2(n25423), .B1(n25310), .B2(n20371), .ZN(
        n6942) );
  OAI22_X1 U20472 ( .A1(n25318), .A2(n25426), .B1(n25311), .B2(n20370), .ZN(
        n6943) );
  OAI22_X1 U20473 ( .A1(n25318), .A2(n25429), .B1(n25312), .B2(n20369), .ZN(
        n6944) );
  OAI22_X1 U20474 ( .A1(n25318), .A2(n25432), .B1(n25310), .B2(n20368), .ZN(
        n6945) );
  OAI22_X1 U20475 ( .A1(n25319), .A2(n25435), .B1(n25311), .B2(n20367), .ZN(
        n6946) );
  OAI22_X1 U20476 ( .A1(n25319), .A2(n25438), .B1(n25312), .B2(n20366), .ZN(
        n6947) );
  OAI22_X1 U20477 ( .A1(n25319), .A2(n25441), .B1(n25310), .B2(n20365), .ZN(
        n6948) );
  OAI22_X1 U20478 ( .A1(n25319), .A2(n25444), .B1(n25311), .B2(n20364), .ZN(
        n6949) );
  OAI22_X1 U20479 ( .A1(n25319), .A2(n25447), .B1(n25312), .B2(n20363), .ZN(
        n6950) );
  OAI22_X1 U20480 ( .A1(n25320), .A2(n25450), .B1(n25310), .B2(n20362), .ZN(
        n6951) );
  OAI22_X1 U20481 ( .A1(n25320), .A2(n25453), .B1(n21257), .B2(n20361), .ZN(
        n6952) );
  OAI22_X1 U20482 ( .A1(n25320), .A2(n25456), .B1(n25310), .B2(n20360), .ZN(
        n6953) );
  OAI22_X1 U20483 ( .A1(n25320), .A2(n25459), .B1(n21257), .B2(n20359), .ZN(
        n6954) );
  OAI22_X1 U20484 ( .A1(n25320), .A2(n25462), .B1(n25310), .B2(n20358), .ZN(
        n6955) );
  OAI22_X1 U20485 ( .A1(n25321), .A2(n25465), .B1(n21257), .B2(n20357), .ZN(
        n6956) );
  OAI22_X1 U20486 ( .A1(n25321), .A2(n25468), .B1(n25310), .B2(n20356), .ZN(
        n6957) );
  OAI22_X1 U20487 ( .A1(n25321), .A2(n25471), .B1(n25311), .B2(n20355), .ZN(
        n6958) );
  OAI22_X1 U20488 ( .A1(n25321), .A2(n25474), .B1(n25312), .B2(n20354), .ZN(
        n6959) );
  OAI22_X1 U20489 ( .A1(n25321), .A2(n25477), .B1(n25310), .B2(n20353), .ZN(
        n6960) );
  OAI22_X1 U20490 ( .A1(n25322), .A2(n25480), .B1(n25310), .B2(n20352), .ZN(
        n6961) );
  OAI22_X1 U20491 ( .A1(n25322), .A2(n25483), .B1(n25311), .B2(n20351), .ZN(
        n6962) );
  OAI22_X1 U20492 ( .A1(n25322), .A2(n25486), .B1(n25312), .B2(n20350), .ZN(
        n6963) );
  OAI22_X1 U20493 ( .A1(n25322), .A2(n25489), .B1(n25310), .B2(n20349), .ZN(
        n6964) );
  OAI22_X1 U20494 ( .A1(n25322), .A2(n25492), .B1(n25310), .B2(n20348), .ZN(
        n6965) );
  OAI22_X1 U20495 ( .A1(n25323), .A2(n25495), .B1(n21257), .B2(n20347), .ZN(
        n6966) );
  OAI22_X1 U20496 ( .A1(n25323), .A2(n25498), .B1(n25310), .B2(n20346), .ZN(
        n6967) );
  OAI22_X1 U20497 ( .A1(n25323), .A2(n25501), .B1(n21257), .B2(n20345), .ZN(
        n6968) );
  OAI22_X1 U20498 ( .A1(n25323), .A2(n25504), .B1(n25310), .B2(n20344), .ZN(
        n6969) );
  OAI22_X1 U20499 ( .A1(n25323), .A2(n25507), .B1(n21257), .B2(n20343), .ZN(
        n6970) );
  OAI22_X1 U20500 ( .A1(n25324), .A2(n25510), .B1(n25310), .B2(n20342), .ZN(
        n6971) );
  OAI22_X1 U20501 ( .A1(n25324), .A2(n25513), .B1(n21257), .B2(n20341), .ZN(
        n6972) );
  OAI22_X1 U20502 ( .A1(n25324), .A2(n25516), .B1(n25310), .B2(n20340), .ZN(
        n6973) );
  OAI22_X1 U20503 ( .A1(n25324), .A2(n25519), .B1(n21257), .B2(n20339), .ZN(
        n6974) );
  OAI22_X1 U20504 ( .A1(n25324), .A2(n25522), .B1(n25310), .B2(n20338), .ZN(
        n6975) );
  OAI22_X1 U20505 ( .A1(n25198), .A2(n25417), .B1(n25192), .B2(n20337), .ZN(
        n6492) );
  OAI22_X1 U20506 ( .A1(n25199), .A2(n25420), .B1(n25193), .B2(n20336), .ZN(
        n6493) );
  OAI22_X1 U20507 ( .A1(n25199), .A2(n25423), .B1(n25191), .B2(n20335), .ZN(
        n6494) );
  OAI22_X1 U20508 ( .A1(n25199), .A2(n25426), .B1(n25192), .B2(n20334), .ZN(
        n6495) );
  OAI22_X1 U20509 ( .A1(n25199), .A2(n25429), .B1(n25193), .B2(n20333), .ZN(
        n6496) );
  OAI22_X1 U20510 ( .A1(n25199), .A2(n25432), .B1(n25191), .B2(n20332), .ZN(
        n6497) );
  OAI22_X1 U20511 ( .A1(n25200), .A2(n25435), .B1(n25192), .B2(n20331), .ZN(
        n6498) );
  OAI22_X1 U20512 ( .A1(n25200), .A2(n25438), .B1(n25193), .B2(n20330), .ZN(
        n6499) );
  OAI22_X1 U20513 ( .A1(n25200), .A2(n25441), .B1(n25191), .B2(n20329), .ZN(
        n6500) );
  OAI22_X1 U20514 ( .A1(n25200), .A2(n25444), .B1(n25192), .B2(n20328), .ZN(
        n6501) );
  OAI22_X1 U20515 ( .A1(n25200), .A2(n25447), .B1(n25193), .B2(n20327), .ZN(
        n6502) );
  OAI22_X1 U20516 ( .A1(n25201), .A2(n25450), .B1(n25191), .B2(n20326), .ZN(
        n6503) );
  OAI22_X1 U20517 ( .A1(n25201), .A2(n25453), .B1(n21272), .B2(n20325), .ZN(
        n6504) );
  OAI22_X1 U20518 ( .A1(n25201), .A2(n25456), .B1(n25191), .B2(n20324), .ZN(
        n6505) );
  OAI22_X1 U20519 ( .A1(n25201), .A2(n25459), .B1(n21272), .B2(n20323), .ZN(
        n6506) );
  OAI22_X1 U20520 ( .A1(n25201), .A2(n25462), .B1(n25191), .B2(n20322), .ZN(
        n6507) );
  OAI22_X1 U20521 ( .A1(n25202), .A2(n25465), .B1(n21272), .B2(n20321), .ZN(
        n6508) );
  OAI22_X1 U20522 ( .A1(n25202), .A2(n25468), .B1(n25191), .B2(n20320), .ZN(
        n6509) );
  OAI22_X1 U20523 ( .A1(n25202), .A2(n25471), .B1(n25192), .B2(n20319), .ZN(
        n6510) );
  OAI22_X1 U20524 ( .A1(n25202), .A2(n25474), .B1(n25193), .B2(n20318), .ZN(
        n6511) );
  OAI22_X1 U20525 ( .A1(n25202), .A2(n25477), .B1(n25191), .B2(n20317), .ZN(
        n6512) );
  OAI22_X1 U20526 ( .A1(n25203), .A2(n25480), .B1(n25191), .B2(n20316), .ZN(
        n6513) );
  OAI22_X1 U20527 ( .A1(n25203), .A2(n25483), .B1(n25192), .B2(n20315), .ZN(
        n6514) );
  OAI22_X1 U20528 ( .A1(n25203), .A2(n25486), .B1(n25193), .B2(n20314), .ZN(
        n6515) );
  OAI22_X1 U20529 ( .A1(n25203), .A2(n25489), .B1(n25191), .B2(n20313), .ZN(
        n6516) );
  OAI22_X1 U20530 ( .A1(n25203), .A2(n25492), .B1(n25191), .B2(n20312), .ZN(
        n6517) );
  OAI22_X1 U20531 ( .A1(n25204), .A2(n25495), .B1(n21272), .B2(n20311), .ZN(
        n6518) );
  OAI22_X1 U20532 ( .A1(n25204), .A2(n25498), .B1(n25191), .B2(n20310), .ZN(
        n6519) );
  OAI22_X1 U20533 ( .A1(n25204), .A2(n25501), .B1(n21272), .B2(n20309), .ZN(
        n6520) );
  OAI22_X1 U20534 ( .A1(n25204), .A2(n25504), .B1(n25191), .B2(n20308), .ZN(
        n6521) );
  OAI22_X1 U20535 ( .A1(n25204), .A2(n25507), .B1(n21272), .B2(n20307), .ZN(
        n6522) );
  OAI22_X1 U20536 ( .A1(n25205), .A2(n25510), .B1(n25191), .B2(n20306), .ZN(
        n6523) );
  OAI22_X1 U20537 ( .A1(n25205), .A2(n25513), .B1(n21272), .B2(n20305), .ZN(
        n6524) );
  OAI22_X1 U20538 ( .A1(n25205), .A2(n25516), .B1(n25191), .B2(n20304), .ZN(
        n6525) );
  OAI22_X1 U20539 ( .A1(n25205), .A2(n25519), .B1(n21272), .B2(n20303), .ZN(
        n6526) );
  OAI22_X1 U20540 ( .A1(n25205), .A2(n25522), .B1(n25191), .B2(n20302), .ZN(
        n6527) );
  OAI22_X1 U20541 ( .A1(n25300), .A2(n25417), .B1(n25294), .B2(n20301), .ZN(
        n6876) );
  OAI22_X1 U20542 ( .A1(n25301), .A2(n25420), .B1(n25295), .B2(n20300), .ZN(
        n6877) );
  OAI22_X1 U20543 ( .A1(n25301), .A2(n25423), .B1(n25293), .B2(n20299), .ZN(
        n6878) );
  OAI22_X1 U20544 ( .A1(n25301), .A2(n25426), .B1(n25294), .B2(n20298), .ZN(
        n6879) );
  OAI22_X1 U20545 ( .A1(n25301), .A2(n25429), .B1(n25295), .B2(n20297), .ZN(
        n6880) );
  OAI22_X1 U20546 ( .A1(n25301), .A2(n25432), .B1(n25293), .B2(n20296), .ZN(
        n6881) );
  OAI22_X1 U20547 ( .A1(n25302), .A2(n25435), .B1(n25294), .B2(n20295), .ZN(
        n6882) );
  OAI22_X1 U20548 ( .A1(n25302), .A2(n25438), .B1(n25295), .B2(n20294), .ZN(
        n6883) );
  OAI22_X1 U20549 ( .A1(n25302), .A2(n25441), .B1(n25293), .B2(n20293), .ZN(
        n6884) );
  OAI22_X1 U20550 ( .A1(n25302), .A2(n25444), .B1(n25294), .B2(n20292), .ZN(
        n6885) );
  OAI22_X1 U20551 ( .A1(n25302), .A2(n25447), .B1(n25295), .B2(n20291), .ZN(
        n6886) );
  OAI22_X1 U20552 ( .A1(n25303), .A2(n25450), .B1(n25293), .B2(n20290), .ZN(
        n6887) );
  OAI22_X1 U20553 ( .A1(n25303), .A2(n25453), .B1(n21259), .B2(n20289), .ZN(
        n6888) );
  OAI22_X1 U20554 ( .A1(n25303), .A2(n25456), .B1(n25293), .B2(n20288), .ZN(
        n6889) );
  OAI22_X1 U20555 ( .A1(n25303), .A2(n25459), .B1(n21259), .B2(n20287), .ZN(
        n6890) );
  OAI22_X1 U20556 ( .A1(n25303), .A2(n25462), .B1(n25293), .B2(n20286), .ZN(
        n6891) );
  OAI22_X1 U20557 ( .A1(n25304), .A2(n25465), .B1(n21259), .B2(n20285), .ZN(
        n6892) );
  OAI22_X1 U20558 ( .A1(n25304), .A2(n25468), .B1(n25293), .B2(n20284), .ZN(
        n6893) );
  OAI22_X1 U20559 ( .A1(n25304), .A2(n25471), .B1(n25294), .B2(n20283), .ZN(
        n6894) );
  OAI22_X1 U20560 ( .A1(n25304), .A2(n25474), .B1(n25295), .B2(n20282), .ZN(
        n6895) );
  OAI22_X1 U20561 ( .A1(n25304), .A2(n25477), .B1(n25293), .B2(n20281), .ZN(
        n6896) );
  OAI22_X1 U20562 ( .A1(n25305), .A2(n25480), .B1(n25293), .B2(n20280), .ZN(
        n6897) );
  OAI22_X1 U20563 ( .A1(n25305), .A2(n25483), .B1(n25294), .B2(n20279), .ZN(
        n6898) );
  OAI22_X1 U20564 ( .A1(n25305), .A2(n25486), .B1(n25295), .B2(n20278), .ZN(
        n6899) );
  OAI22_X1 U20565 ( .A1(n25305), .A2(n25489), .B1(n25293), .B2(n20277), .ZN(
        n6900) );
  OAI22_X1 U20566 ( .A1(n25305), .A2(n25492), .B1(n25293), .B2(n20276), .ZN(
        n6901) );
  OAI22_X1 U20567 ( .A1(n25306), .A2(n25495), .B1(n21259), .B2(n20275), .ZN(
        n6902) );
  OAI22_X1 U20568 ( .A1(n25306), .A2(n25498), .B1(n25293), .B2(n20274), .ZN(
        n6903) );
  OAI22_X1 U20569 ( .A1(n25306), .A2(n25501), .B1(n21259), .B2(n20273), .ZN(
        n6904) );
  OAI22_X1 U20570 ( .A1(n25306), .A2(n25504), .B1(n25293), .B2(n20272), .ZN(
        n6905) );
  OAI22_X1 U20571 ( .A1(n25306), .A2(n25507), .B1(n21259), .B2(n20271), .ZN(
        n6906) );
  OAI22_X1 U20572 ( .A1(n25307), .A2(n25510), .B1(n25293), .B2(n20270), .ZN(
        n6907) );
  OAI22_X1 U20573 ( .A1(n25307), .A2(n25513), .B1(n21259), .B2(n20269), .ZN(
        n6908) );
  OAI22_X1 U20574 ( .A1(n25307), .A2(n25516), .B1(n25293), .B2(n20268), .ZN(
        n6909) );
  OAI22_X1 U20575 ( .A1(n25307), .A2(n25519), .B1(n21259), .B2(n20267), .ZN(
        n6910) );
  OAI22_X1 U20576 ( .A1(n25307), .A2(n25522), .B1(n25293), .B2(n20266), .ZN(
        n6911) );
  OAI22_X1 U20577 ( .A1(n24877), .A2(n25437), .B1(n24868), .B2(n20186), .ZN(
        n5282) );
  OAI22_X1 U20578 ( .A1(n24877), .A2(n25440), .B1(n24868), .B2(n20185), .ZN(
        n5283) );
  OAI22_X1 U20579 ( .A1(n24877), .A2(n25443), .B1(n21293), .B2(n20184), .ZN(
        n5284) );
  OAI22_X1 U20580 ( .A1(n24877), .A2(n25446), .B1(n24868), .B2(n20183), .ZN(
        n5285) );
  OAI22_X1 U20581 ( .A1(n24877), .A2(n25449), .B1(n21293), .B2(n20182), .ZN(
        n5286) );
  OAI22_X1 U20582 ( .A1(n24878), .A2(n25452), .B1(n24868), .B2(n20181), .ZN(
        n5287) );
  OAI22_X1 U20583 ( .A1(n24878), .A2(n25455), .B1(n24869), .B2(n20180), .ZN(
        n5288) );
  OAI22_X1 U20584 ( .A1(n24878), .A2(n25458), .B1(n24870), .B2(n20179), .ZN(
        n5289) );
  OAI22_X1 U20585 ( .A1(n24878), .A2(n25461), .B1(n24868), .B2(n20178), .ZN(
        n5290) );
  OAI22_X1 U20586 ( .A1(n24878), .A2(n25464), .B1(n24869), .B2(n20177), .ZN(
        n5291) );
  OAI22_X1 U20587 ( .A1(n24879), .A2(n25467), .B1(n24870), .B2(n20176), .ZN(
        n5292) );
  OAI22_X1 U20588 ( .A1(n24879), .A2(n25470), .B1(n24868), .B2(n20175), .ZN(
        n5293) );
  OAI22_X1 U20589 ( .A1(n24879), .A2(n25473), .B1(n24869), .B2(n20174), .ZN(
        n5294) );
  OAI22_X1 U20590 ( .A1(n24879), .A2(n25476), .B1(n24870), .B2(n20173), .ZN(
        n5295) );
  OAI22_X1 U20591 ( .A1(n24879), .A2(n25479), .B1(n24868), .B2(n20172), .ZN(
        n5296) );
  OAI22_X1 U20592 ( .A1(n24880), .A2(n25482), .B1(n24869), .B2(n20171), .ZN(
        n5297) );
  OAI22_X1 U20593 ( .A1(n24880), .A2(n25485), .B1(n24870), .B2(n20170), .ZN(
        n5298) );
  OAI22_X1 U20594 ( .A1(n24880), .A2(n25488), .B1(n24868), .B2(n20169), .ZN(
        n5299) );
  OAI22_X1 U20595 ( .A1(n24880), .A2(n25491), .B1(n21293), .B2(n20168), .ZN(
        n5300) );
  OAI22_X1 U20596 ( .A1(n24880), .A2(n25494), .B1(n24868), .B2(n20167), .ZN(
        n5301) );
  OAI22_X1 U20597 ( .A1(n24881), .A2(n25497), .B1(n21293), .B2(n20166), .ZN(
        n5302) );
  OAI22_X1 U20598 ( .A1(n24881), .A2(n25500), .B1(n24868), .B2(n20165), .ZN(
        n5303) );
  OAI22_X1 U20599 ( .A1(n24881), .A2(n25503), .B1(n21293), .B2(n20164), .ZN(
        n5304) );
  OAI22_X1 U20600 ( .A1(n24881), .A2(n25506), .B1(n24868), .B2(n20163), .ZN(
        n5305) );
  OAI22_X1 U20601 ( .A1(n24881), .A2(n25509), .B1(n24869), .B2(n20162), .ZN(
        n5306) );
  OAI22_X1 U20602 ( .A1(n24882), .A2(n25512), .B1(n24870), .B2(n20161), .ZN(
        n5307) );
  OAI22_X1 U20603 ( .A1(n24882), .A2(n25515), .B1(n24868), .B2(n20160), .ZN(
        n5308) );
  OAI22_X1 U20604 ( .A1(n24882), .A2(n25518), .B1(n24868), .B2(n20159), .ZN(
        n5309) );
  OAI22_X1 U20605 ( .A1(n24882), .A2(n25521), .B1(n24869), .B2(n20158), .ZN(
        n5310) );
  OAI22_X1 U20606 ( .A1(n24882), .A2(n25524), .B1(n24870), .B2(n20157), .ZN(
        n5311) );
  OAI22_X1 U20607 ( .A1(n24875), .A2(n25419), .B1(n21293), .B2(n19713), .ZN(
        n5276) );
  OAI22_X1 U20608 ( .A1(n24876), .A2(n25422), .B1(n24868), .B2(n19712), .ZN(
        n5277) );
  OAI22_X1 U20609 ( .A1(n24876), .A2(n25425), .B1(n21293), .B2(n19711), .ZN(
        n5278) );
  OAI22_X1 U20610 ( .A1(n24876), .A2(n25428), .B1(n24868), .B2(n19710), .ZN(
        n5279) );
  OAI22_X1 U20611 ( .A1(n24876), .A2(n25431), .B1(n21293), .B2(n19709), .ZN(
        n5280) );
  OAI22_X1 U20612 ( .A1(n24876), .A2(n25434), .B1(n24868), .B2(n19708), .ZN(
        n5281) );
  OAI22_X1 U20613 ( .A1(n24943), .A2(n25419), .B1(n24937), .B2(n19683), .ZN(
        n5532) );
  OAI22_X1 U20614 ( .A1(n24944), .A2(n25422), .B1(n24938), .B2(n19682), .ZN(
        n5533) );
  OAI22_X1 U20615 ( .A1(n24944), .A2(n25425), .B1(n24936), .B2(n19681), .ZN(
        n5534) );
  OAI22_X1 U20616 ( .A1(n24944), .A2(n25428), .B1(n24937), .B2(n19680), .ZN(
        n5535) );
  OAI22_X1 U20617 ( .A1(n24944), .A2(n25431), .B1(n24938), .B2(n19679), .ZN(
        n5536) );
  OAI22_X1 U20618 ( .A1(n24944), .A2(n25434), .B1(n24936), .B2(n19678), .ZN(
        n5537) );
  OAI22_X1 U20619 ( .A1(n24945), .A2(n25437), .B1(n24937), .B2(n19677), .ZN(
        n5538) );
  OAI22_X1 U20620 ( .A1(n24945), .A2(n25440), .B1(n24938), .B2(n19676), .ZN(
        n5539) );
  OAI22_X1 U20621 ( .A1(n24945), .A2(n25443), .B1(n24936), .B2(n19675), .ZN(
        n5540) );
  OAI22_X1 U20622 ( .A1(n24945), .A2(n25446), .B1(n24937), .B2(n19674), .ZN(
        n5541) );
  OAI22_X1 U20623 ( .A1(n24945), .A2(n25449), .B1(n24938), .B2(n19673), .ZN(
        n5542) );
  OAI22_X1 U20624 ( .A1(n24946), .A2(n25452), .B1(n24936), .B2(n19672), .ZN(
        n5543) );
  OAI22_X1 U20625 ( .A1(n24946), .A2(n25455), .B1(n21288), .B2(n19671), .ZN(
        n5544) );
  OAI22_X1 U20626 ( .A1(n24946), .A2(n25458), .B1(n24936), .B2(n19670), .ZN(
        n5545) );
  OAI22_X1 U20627 ( .A1(n24946), .A2(n25461), .B1(n21288), .B2(n19669), .ZN(
        n5546) );
  OAI22_X1 U20628 ( .A1(n24946), .A2(n25464), .B1(n24936), .B2(n19668), .ZN(
        n5547) );
  OAI22_X1 U20629 ( .A1(n24947), .A2(n25467), .B1(n21288), .B2(n19667), .ZN(
        n5548) );
  OAI22_X1 U20630 ( .A1(n24947), .A2(n25470), .B1(n24936), .B2(n19666), .ZN(
        n5549) );
  OAI22_X1 U20631 ( .A1(n24947), .A2(n25473), .B1(n24937), .B2(n19665), .ZN(
        n5550) );
  OAI22_X1 U20632 ( .A1(n24947), .A2(n25476), .B1(n24938), .B2(n19664), .ZN(
        n5551) );
  OAI22_X1 U20633 ( .A1(n24947), .A2(n25479), .B1(n24936), .B2(n19663), .ZN(
        n5552) );
  OAI22_X1 U20634 ( .A1(n24948), .A2(n25482), .B1(n24936), .B2(n19662), .ZN(
        n5553) );
  OAI22_X1 U20635 ( .A1(n24948), .A2(n25485), .B1(n24937), .B2(n19661), .ZN(
        n5554) );
  OAI22_X1 U20636 ( .A1(n24948), .A2(n25488), .B1(n24938), .B2(n19660), .ZN(
        n5555) );
  OAI22_X1 U20637 ( .A1(n24948), .A2(n25491), .B1(n24936), .B2(n19659), .ZN(
        n5556) );
  OAI22_X1 U20638 ( .A1(n24948), .A2(n25494), .B1(n24936), .B2(n19658), .ZN(
        n5557) );
  OAI22_X1 U20639 ( .A1(n24949), .A2(n25497), .B1(n21288), .B2(n19657), .ZN(
        n5558) );
  OAI22_X1 U20640 ( .A1(n24949), .A2(n25500), .B1(n24936), .B2(n19656), .ZN(
        n5559) );
  OAI22_X1 U20641 ( .A1(n24949), .A2(n25503), .B1(n21288), .B2(n19655), .ZN(
        n5560) );
  OAI22_X1 U20642 ( .A1(n24949), .A2(n25506), .B1(n24936), .B2(n19654), .ZN(
        n5561) );
  OAI22_X1 U20643 ( .A1(n24949), .A2(n25509), .B1(n21288), .B2(n19653), .ZN(
        n5562) );
  OAI22_X1 U20644 ( .A1(n24950), .A2(n25512), .B1(n24936), .B2(n19652), .ZN(
        n5563) );
  OAI22_X1 U20645 ( .A1(n24950), .A2(n25515), .B1(n21288), .B2(n19651), .ZN(
        n5564) );
  OAI22_X1 U20646 ( .A1(n24950), .A2(n25518), .B1(n24936), .B2(n19650), .ZN(
        n5565) );
  OAI22_X1 U20647 ( .A1(n24950), .A2(n25521), .B1(n21288), .B2(n19649), .ZN(
        n5566) );
  OAI22_X1 U20648 ( .A1(n24950), .A2(n25524), .B1(n24936), .B2(n19648), .ZN(
        n5567) );
  OAI22_X1 U20649 ( .A1(n25283), .A2(n25417), .B1(n25277), .B2(n19371), .ZN(
        n6812) );
  OAI22_X1 U20650 ( .A1(n25284), .A2(n25420), .B1(n25278), .B2(n19370), .ZN(
        n6813) );
  OAI22_X1 U20651 ( .A1(n25284), .A2(n25423), .B1(n25276), .B2(n19369), .ZN(
        n6814) );
  OAI22_X1 U20652 ( .A1(n25284), .A2(n25426), .B1(n25277), .B2(n19368), .ZN(
        n6815) );
  OAI22_X1 U20653 ( .A1(n25284), .A2(n25429), .B1(n25278), .B2(n19367), .ZN(
        n6816) );
  OAI22_X1 U20654 ( .A1(n25284), .A2(n25432), .B1(n25276), .B2(n19366), .ZN(
        n6817) );
  OAI22_X1 U20655 ( .A1(n25285), .A2(n25435), .B1(n25277), .B2(n19365), .ZN(
        n6818) );
  OAI22_X1 U20656 ( .A1(n25285), .A2(n25438), .B1(n25278), .B2(n19364), .ZN(
        n6819) );
  OAI22_X1 U20657 ( .A1(n25285), .A2(n25441), .B1(n25276), .B2(n19363), .ZN(
        n6820) );
  OAI22_X1 U20658 ( .A1(n25285), .A2(n25444), .B1(n25277), .B2(n19362), .ZN(
        n6821) );
  OAI22_X1 U20659 ( .A1(n25285), .A2(n25447), .B1(n25278), .B2(n19361), .ZN(
        n6822) );
  OAI22_X1 U20660 ( .A1(n25286), .A2(n25450), .B1(n25276), .B2(n19360), .ZN(
        n6823) );
  OAI22_X1 U20661 ( .A1(n25286), .A2(n25453), .B1(n21261), .B2(n19359), .ZN(
        n6824) );
  OAI22_X1 U20662 ( .A1(n25286), .A2(n25456), .B1(n25276), .B2(n19358), .ZN(
        n6825) );
  OAI22_X1 U20663 ( .A1(n25286), .A2(n25459), .B1(n21261), .B2(n19357), .ZN(
        n6826) );
  OAI22_X1 U20664 ( .A1(n25286), .A2(n25462), .B1(n25276), .B2(n19356), .ZN(
        n6827) );
  OAI22_X1 U20665 ( .A1(n25287), .A2(n25465), .B1(n21261), .B2(n19355), .ZN(
        n6828) );
  OAI22_X1 U20666 ( .A1(n25287), .A2(n25468), .B1(n25276), .B2(n19354), .ZN(
        n6829) );
  OAI22_X1 U20667 ( .A1(n25287), .A2(n25471), .B1(n25277), .B2(n19353), .ZN(
        n6830) );
  OAI22_X1 U20668 ( .A1(n25287), .A2(n25474), .B1(n25278), .B2(n19352), .ZN(
        n6831) );
  OAI22_X1 U20669 ( .A1(n25287), .A2(n25477), .B1(n25276), .B2(n19351), .ZN(
        n6832) );
  OAI22_X1 U20670 ( .A1(n25288), .A2(n25480), .B1(n25276), .B2(n19350), .ZN(
        n6833) );
  OAI22_X1 U20671 ( .A1(n25288), .A2(n25483), .B1(n25277), .B2(n19349), .ZN(
        n6834) );
  OAI22_X1 U20672 ( .A1(n25288), .A2(n25486), .B1(n25278), .B2(n19348), .ZN(
        n6835) );
  OAI22_X1 U20673 ( .A1(n25288), .A2(n25489), .B1(n25276), .B2(n19347), .ZN(
        n6836) );
  OAI22_X1 U20674 ( .A1(n25288), .A2(n25492), .B1(n25276), .B2(n19346), .ZN(
        n6837) );
  OAI22_X1 U20675 ( .A1(n25289), .A2(n25495), .B1(n21261), .B2(n19345), .ZN(
        n6838) );
  OAI22_X1 U20676 ( .A1(n25289), .A2(n25498), .B1(n25276), .B2(n19344), .ZN(
        n6839) );
  OAI22_X1 U20677 ( .A1(n25289), .A2(n25501), .B1(n21261), .B2(n19343), .ZN(
        n6840) );
  OAI22_X1 U20678 ( .A1(n25289), .A2(n25504), .B1(n25276), .B2(n19342), .ZN(
        n6841) );
  OAI22_X1 U20679 ( .A1(n25289), .A2(n25507), .B1(n21261), .B2(n19341), .ZN(
        n6842) );
  OAI22_X1 U20680 ( .A1(n25290), .A2(n25510), .B1(n25276), .B2(n19340), .ZN(
        n6843) );
  OAI22_X1 U20681 ( .A1(n25290), .A2(n25513), .B1(n21261), .B2(n19339), .ZN(
        n6844) );
  OAI22_X1 U20682 ( .A1(n25290), .A2(n25516), .B1(n25276), .B2(n19338), .ZN(
        n6845) );
  OAI22_X1 U20683 ( .A1(n25290), .A2(n25519), .B1(n21261), .B2(n19337), .ZN(
        n6846) );
  OAI22_X1 U20684 ( .A1(n25290), .A2(n25522), .B1(n25276), .B2(n19336), .ZN(
        n6847) );
  OAI22_X1 U20685 ( .A1(n25541), .A2(n25417), .B1(n25535), .B2(n19307), .ZN(
        n7068) );
  OAI22_X1 U20686 ( .A1(n25542), .A2(n25420), .B1(n25536), .B2(n19306), .ZN(
        n7069) );
  OAI22_X1 U20687 ( .A1(n25542), .A2(n25423), .B1(n25534), .B2(n19305), .ZN(
        n7070) );
  OAI22_X1 U20688 ( .A1(n25542), .A2(n25426), .B1(n25535), .B2(n19304), .ZN(
        n7071) );
  OAI22_X1 U20689 ( .A1(n25542), .A2(n25429), .B1(n25536), .B2(n19303), .ZN(
        n7072) );
  OAI22_X1 U20690 ( .A1(n25542), .A2(n25432), .B1(n25534), .B2(n19302), .ZN(
        n7073) );
  OAI22_X1 U20691 ( .A1(n25543), .A2(n25435), .B1(n25535), .B2(n19301), .ZN(
        n7074) );
  OAI22_X1 U20692 ( .A1(n25543), .A2(n25438), .B1(n25536), .B2(n19300), .ZN(
        n7075) );
  OAI22_X1 U20693 ( .A1(n25543), .A2(n25441), .B1(n25534), .B2(n19299), .ZN(
        n7076) );
  OAI22_X1 U20694 ( .A1(n25543), .A2(n25444), .B1(n25535), .B2(n19298), .ZN(
        n7077) );
  OAI22_X1 U20695 ( .A1(n25543), .A2(n25447), .B1(n25536), .B2(n19297), .ZN(
        n7078) );
  OAI22_X1 U20696 ( .A1(n25544), .A2(n25450), .B1(n25534), .B2(n19296), .ZN(
        n7079) );
  OAI22_X1 U20697 ( .A1(n25544), .A2(n25453), .B1(n21189), .B2(n19295), .ZN(
        n7080) );
  OAI22_X1 U20698 ( .A1(n25544), .A2(n25456), .B1(n25534), .B2(n19294), .ZN(
        n7081) );
  OAI22_X1 U20699 ( .A1(n25544), .A2(n25459), .B1(n21189), .B2(n19293), .ZN(
        n7082) );
  OAI22_X1 U20700 ( .A1(n25544), .A2(n25462), .B1(n25534), .B2(n19292), .ZN(
        n7083) );
  OAI22_X1 U20701 ( .A1(n25545), .A2(n25465), .B1(n21189), .B2(n19291), .ZN(
        n7084) );
  OAI22_X1 U20702 ( .A1(n25545), .A2(n25468), .B1(n25534), .B2(n19290), .ZN(
        n7085) );
  OAI22_X1 U20703 ( .A1(n25545), .A2(n25471), .B1(n25535), .B2(n19289), .ZN(
        n7086) );
  OAI22_X1 U20704 ( .A1(n25545), .A2(n25474), .B1(n25536), .B2(n19288), .ZN(
        n7087) );
  OAI22_X1 U20705 ( .A1(n25545), .A2(n25477), .B1(n25534), .B2(n19287), .ZN(
        n7088) );
  OAI22_X1 U20706 ( .A1(n25546), .A2(n25480), .B1(n25534), .B2(n19286), .ZN(
        n7089) );
  OAI22_X1 U20707 ( .A1(n25546), .A2(n25483), .B1(n25535), .B2(n19285), .ZN(
        n7090) );
  OAI22_X1 U20708 ( .A1(n25546), .A2(n25486), .B1(n25536), .B2(n19284), .ZN(
        n7091) );
  OAI22_X1 U20709 ( .A1(n25546), .A2(n25489), .B1(n25534), .B2(n19283), .ZN(
        n7092) );
  OAI22_X1 U20710 ( .A1(n25546), .A2(n25492), .B1(n25534), .B2(n19282), .ZN(
        n7093) );
  OAI22_X1 U20711 ( .A1(n25547), .A2(n25495), .B1(n21189), .B2(n19281), .ZN(
        n7094) );
  OAI22_X1 U20712 ( .A1(n25547), .A2(n25498), .B1(n25534), .B2(n19280), .ZN(
        n7095) );
  OAI22_X1 U20713 ( .A1(n25547), .A2(n25501), .B1(n21189), .B2(n19279), .ZN(
        n7096) );
  OAI22_X1 U20714 ( .A1(n25547), .A2(n25504), .B1(n25534), .B2(n19278), .ZN(
        n7097) );
  OAI22_X1 U20715 ( .A1(n25547), .A2(n25507), .B1(n21189), .B2(n19277), .ZN(
        n7098) );
  OAI22_X1 U20716 ( .A1(n25548), .A2(n25510), .B1(n25534), .B2(n19276), .ZN(
        n7099) );
  OAI22_X1 U20717 ( .A1(n25548), .A2(n25513), .B1(n21189), .B2(n19275), .ZN(
        n7100) );
  OAI22_X1 U20718 ( .A1(n25548), .A2(n25516), .B1(n25534), .B2(n19274), .ZN(
        n7101) );
  OAI22_X1 U20719 ( .A1(n25548), .A2(n25519), .B1(n21189), .B2(n19273), .ZN(
        n7102) );
  OAI22_X1 U20720 ( .A1(n25548), .A2(n25522), .B1(n25534), .B2(n19272), .ZN(
        n7103) );
  OAI22_X1 U20721 ( .A1(n25330), .A2(n25348), .B1(n21255), .B2(n21147), .ZN(
        n6981) );
  OAI22_X1 U20722 ( .A1(n25002), .A2(n25526), .B1(n21285), .B2(n20546), .ZN(
        n5760) );
  OAI22_X1 U20723 ( .A1(n25002), .A2(n25529), .B1(n21285), .B2(n20545), .ZN(
        n5761) );
  OAI22_X1 U20724 ( .A1(n25002), .A2(n25532), .B1(n24987), .B2(n20544), .ZN(
        n5762) );
  OAI22_X1 U20725 ( .A1(n25002), .A2(n25552), .B1(n21285), .B2(n20543), .ZN(
        n5763) );
  OAI22_X1 U20726 ( .A1(n25240), .A2(n25525), .B1(n21267), .B2(n20542), .ZN(
        n6656) );
  OAI22_X1 U20727 ( .A1(n25240), .A2(n25528), .B1(n21267), .B2(n20541), .ZN(
        n6657) );
  OAI22_X1 U20728 ( .A1(n25240), .A2(n25531), .B1(n25225), .B2(n20540), .ZN(
        n6658) );
  OAI22_X1 U20729 ( .A1(n25240), .A2(n25551), .B1(n21267), .B2(n20539), .ZN(
        n6659) );
  OAI22_X1 U20730 ( .A1(n25223), .A2(n25525), .B1(n21270), .B2(n20538), .ZN(
        n6592) );
  OAI22_X1 U20731 ( .A1(n25223), .A2(n25528), .B1(n21270), .B2(n20537), .ZN(
        n6593) );
  OAI22_X1 U20732 ( .A1(n25223), .A2(n25531), .B1(n25208), .B2(n20536), .ZN(
        n6594) );
  OAI22_X1 U20733 ( .A1(n25223), .A2(n25551), .B1(n21270), .B2(n20535), .ZN(
        n6595) );
  OAI22_X1 U20734 ( .A1(n25155), .A2(n25526), .B1(n21275), .B2(n20534), .ZN(
        n6336) );
  OAI22_X1 U20735 ( .A1(n25155), .A2(n25529), .B1(n21275), .B2(n20533), .ZN(
        n6337) );
  OAI22_X1 U20736 ( .A1(n25155), .A2(n25532), .B1(n25140), .B2(n20532), .ZN(
        n6338) );
  OAI22_X1 U20737 ( .A1(n25155), .A2(n25552), .B1(n21275), .B2(n20531), .ZN(
        n6339) );
  OAI22_X1 U20738 ( .A1(n25257), .A2(n25525), .B1(n21265), .B2(n20525), .ZN(
        n6720) );
  OAI22_X1 U20739 ( .A1(n25257), .A2(n25528), .B1(n21265), .B2(n20524), .ZN(
        n6721) );
  OAI22_X1 U20740 ( .A1(n25257), .A2(n25531), .B1(n25242), .B2(n20523), .ZN(
        n6722) );
  OAI22_X1 U20741 ( .A1(n25257), .A2(n25551), .B1(n21265), .B2(n20522), .ZN(
        n6723) );
  OAI22_X1 U20742 ( .A1(n25087), .A2(n25526), .B1(n21279), .B2(n20521), .ZN(
        n6080) );
  OAI22_X1 U20743 ( .A1(n25087), .A2(n25529), .B1(n21279), .B2(n20520), .ZN(
        n6081) );
  OAI22_X1 U20744 ( .A1(n25087), .A2(n25532), .B1(n25072), .B2(n20519), .ZN(
        n6082) );
  OAI22_X1 U20745 ( .A1(n25087), .A2(n25552), .B1(n21279), .B2(n20518), .ZN(
        n6083) );
  OAI22_X1 U20746 ( .A1(n25019), .A2(n25526), .B1(n21284), .B2(n20517), .ZN(
        n5824) );
  OAI22_X1 U20747 ( .A1(n25019), .A2(n25529), .B1(n21284), .B2(n20516), .ZN(
        n5825) );
  OAI22_X1 U20748 ( .A1(n25019), .A2(n25532), .B1(n25004), .B2(n20515), .ZN(
        n5826) );
  OAI22_X1 U20749 ( .A1(n25019), .A2(n25552), .B1(n21284), .B2(n20514), .ZN(
        n5827) );
  OAI22_X1 U20750 ( .A1(n24917), .A2(n25527), .B1(n21291), .B2(n20513), .ZN(
        n5440) );
  OAI22_X1 U20751 ( .A1(n24917), .A2(n25530), .B1(n21291), .B2(n20512), .ZN(
        n5441) );
  OAI22_X1 U20752 ( .A1(n24917), .A2(n25533), .B1(n24902), .B2(n20511), .ZN(
        n5442) );
  OAI22_X1 U20753 ( .A1(n24917), .A2(n25553), .B1(n21291), .B2(n20510), .ZN(
        n5443) );
  OAI22_X1 U20754 ( .A1(n24849), .A2(n25527), .B1(n21295), .B2(n20509), .ZN(
        n5184) );
  OAI22_X1 U20755 ( .A1(n24849), .A2(n25530), .B1(n21295), .B2(n20508), .ZN(
        n5185) );
  OAI22_X1 U20756 ( .A1(n24849), .A2(n25533), .B1(n24834), .B2(n20507), .ZN(
        n5186) );
  OAI22_X1 U20757 ( .A1(n24849), .A2(n25553), .B1(n21295), .B2(n20506), .ZN(
        n5187) );
  OAI22_X1 U20758 ( .A1(n25070), .A2(n25526), .B1(n21281), .B2(n20265), .ZN(
        n6016) );
  OAI22_X1 U20759 ( .A1(n25070), .A2(n25529), .B1(n21281), .B2(n20264), .ZN(
        n6017) );
  OAI22_X1 U20760 ( .A1(n25070), .A2(n25532), .B1(n25055), .B2(n20263), .ZN(
        n6018) );
  OAI22_X1 U20761 ( .A1(n25070), .A2(n25552), .B1(n21281), .B2(n20262), .ZN(
        n6019) );
  OAI22_X1 U20762 ( .A1(n25325), .A2(n25525), .B1(n21257), .B2(n20261), .ZN(
        n6976) );
  OAI22_X1 U20763 ( .A1(n25325), .A2(n25528), .B1(n21257), .B2(n20260), .ZN(
        n6977) );
  OAI22_X1 U20764 ( .A1(n25325), .A2(n25531), .B1(n25310), .B2(n20259), .ZN(
        n6978) );
  OAI22_X1 U20765 ( .A1(n25325), .A2(n25551), .B1(n21257), .B2(n20258), .ZN(
        n6979) );
  OAI22_X1 U20766 ( .A1(n25206), .A2(n25525), .B1(n21272), .B2(n20257), .ZN(
        n6528) );
  OAI22_X1 U20767 ( .A1(n25206), .A2(n25528), .B1(n21272), .B2(n20256), .ZN(
        n6529) );
  OAI22_X1 U20768 ( .A1(n25206), .A2(n25531), .B1(n25191), .B2(n20255), .ZN(
        n6530) );
  OAI22_X1 U20769 ( .A1(n25206), .A2(n25551), .B1(n21272), .B2(n20254), .ZN(
        n6531) );
  OAI22_X1 U20770 ( .A1(n25308), .A2(n25525), .B1(n21259), .B2(n20253), .ZN(
        n6912) );
  OAI22_X1 U20771 ( .A1(n25308), .A2(n25528), .B1(n21259), .B2(n20252), .ZN(
        n6913) );
  OAI22_X1 U20772 ( .A1(n25308), .A2(n25531), .B1(n25293), .B2(n20251), .ZN(
        n6914) );
  OAI22_X1 U20773 ( .A1(n25308), .A2(n25551), .B1(n21259), .B2(n20250), .ZN(
        n6915) );
  OAI22_X1 U20774 ( .A1(n24951), .A2(n25527), .B1(n21288), .B2(n20152), .ZN(
        n5568) );
  OAI22_X1 U20775 ( .A1(n24951), .A2(n25530), .B1(n21288), .B2(n20151), .ZN(
        n5569) );
  OAI22_X1 U20776 ( .A1(n24951), .A2(n25533), .B1(n24936), .B2(n20150), .ZN(
        n5570) );
  OAI22_X1 U20777 ( .A1(n24951), .A2(n25553), .B1(n21288), .B2(n20149), .ZN(
        n5571) );
  OAI22_X1 U20778 ( .A1(n24883), .A2(n25527), .B1(n21293), .B2(n20148), .ZN(
        n5312) );
  OAI22_X1 U20779 ( .A1(n24883), .A2(n25530), .B1(n21293), .B2(n20147), .ZN(
        n5313) );
  OAI22_X1 U20780 ( .A1(n24883), .A2(n25533), .B1(n24868), .B2(n20146), .ZN(
        n5314) );
  OAI22_X1 U20781 ( .A1(n24883), .A2(n25553), .B1(n21293), .B2(n20145), .ZN(
        n5315) );
  OAI22_X1 U20782 ( .A1(n25291), .A2(n25525), .B1(n21261), .B2(n19335), .ZN(
        n6848) );
  OAI22_X1 U20783 ( .A1(n25291), .A2(n25528), .B1(n21261), .B2(n19334), .ZN(
        n6849) );
  OAI22_X1 U20784 ( .A1(n25291), .A2(n25531), .B1(n25276), .B2(n19333), .ZN(
        n6850) );
  OAI22_X1 U20785 ( .A1(n25291), .A2(n25551), .B1(n21261), .B2(n19332), .ZN(
        n6851) );
  OAI22_X1 U20786 ( .A1(n25549), .A2(n25525), .B1(n21189), .B2(n19271), .ZN(
        n7104) );
  OAI22_X1 U20787 ( .A1(n25549), .A2(n25528), .B1(n21189), .B2(n19270), .ZN(
        n7105) );
  OAI22_X1 U20788 ( .A1(n25549), .A2(n25531), .B1(n25534), .B2(n19269), .ZN(
        n7106) );
  OAI22_X1 U20789 ( .A1(n25549), .A2(n25551), .B1(n21189), .B2(n19268), .ZN(
        n7107) );
  NOR3_X1 U20790 ( .A1(n19203), .A2(n19199), .A3(n19200), .ZN(n23739) );
  BUF_X1 U20791 ( .A(n21298), .Z(n24802) );
  BUF_X1 U20792 ( .A(n21298), .Z(n24801) );
  BUF_X1 U20793 ( .A(n21298), .Z(n24799) );
  BUF_X1 U20794 ( .A(n21298), .Z(n24798) );
  BUF_X1 U20795 ( .A(n21298), .Z(n24800) );
  BUF_X1 U20796 ( .A(n22608), .Z(n24409) );
  BUF_X1 U20797 ( .A(n22608), .Z(n24412) );
  BUF_X1 U20798 ( .A(n22608), .Z(n24411) );
  BUF_X1 U20799 ( .A(n22608), .Z(n24410) );
  BUF_X1 U20800 ( .A(n21297), .Z(n24805) );
  BUF_X1 U20801 ( .A(n21297), .Z(n24806) );
  BUF_X1 U20802 ( .A(n21297), .Z(n24807) );
  BUF_X1 U20803 ( .A(n21297), .Z(n24808) );
  NAND2_X1 U20804 ( .A1(n22542), .A2(n22554), .ZN(n21339) );
  NAND2_X1 U20805 ( .A1(n22542), .A2(n22553), .ZN(n21340) );
  NAND2_X1 U20806 ( .A1(n23748), .A2(n23744), .ZN(n22610) );
  NAND2_X1 U20807 ( .A1(n23742), .A2(n23747), .ZN(n22584) );
  NOR2_X1 U20808 ( .A1(n19202), .A2(n19201), .ZN(n23755) );
  BUF_X1 U20809 ( .A(n21252), .Z(n25346) );
  BUF_X1 U20810 ( .A(n21251), .Z(n25349) );
  BUF_X1 U20811 ( .A(n21250), .Z(n25352) );
  BUF_X1 U20812 ( .A(n21249), .Z(n25355) );
  BUF_X1 U20813 ( .A(n21248), .Z(n25358) );
  BUF_X1 U20814 ( .A(n21247), .Z(n25361) );
  BUF_X1 U20815 ( .A(n21246), .Z(n25364) );
  BUF_X1 U20816 ( .A(n21245), .Z(n25367) );
  BUF_X1 U20817 ( .A(n21244), .Z(n25370) );
  BUF_X1 U20818 ( .A(n21243), .Z(n25373) );
  BUF_X1 U20819 ( .A(n21242), .Z(n25376) );
  BUF_X1 U20820 ( .A(n21241), .Z(n25379) );
  BUF_X1 U20821 ( .A(n21240), .Z(n25382) );
  BUF_X1 U20822 ( .A(n21239), .Z(n25385) );
  BUF_X1 U20823 ( .A(n21238), .Z(n25388) );
  BUF_X1 U20824 ( .A(n21237), .Z(n25391) );
  BUF_X1 U20825 ( .A(n21236), .Z(n25394) );
  BUF_X1 U20826 ( .A(n21235), .Z(n25397) );
  BUF_X1 U20827 ( .A(n21234), .Z(n25400) );
  BUF_X1 U20828 ( .A(n21233), .Z(n25403) );
  BUF_X1 U20829 ( .A(n21232), .Z(n25406) );
  BUF_X1 U20830 ( .A(n21231), .Z(n25409) );
  BUF_X1 U20831 ( .A(n21230), .Z(n25412) );
  BUF_X1 U20832 ( .A(n21229), .Z(n25415) );
  BUF_X1 U20833 ( .A(n21228), .Z(n25418) );
  BUF_X1 U20834 ( .A(n21227), .Z(n25421) );
  BUF_X1 U20835 ( .A(n21226), .Z(n25424) );
  BUF_X1 U20836 ( .A(n21225), .Z(n25427) );
  BUF_X1 U20837 ( .A(n21224), .Z(n25430) );
  BUF_X1 U20838 ( .A(n21223), .Z(n25433) );
  BUF_X1 U20839 ( .A(n21222), .Z(n25436) );
  BUF_X1 U20840 ( .A(n21221), .Z(n25439) );
  BUF_X1 U20841 ( .A(n21220), .Z(n25442) );
  BUF_X1 U20842 ( .A(n21219), .Z(n25445) );
  BUF_X1 U20843 ( .A(n21218), .Z(n25448) );
  BUF_X1 U20844 ( .A(n21217), .Z(n25451) );
  BUF_X1 U20845 ( .A(n21216), .Z(n25454) );
  BUF_X1 U20846 ( .A(n21215), .Z(n25457) );
  BUF_X1 U20847 ( .A(n21214), .Z(n25460) );
  BUF_X1 U20848 ( .A(n21213), .Z(n25463) );
  BUF_X1 U20849 ( .A(n21212), .Z(n25466) );
  BUF_X1 U20850 ( .A(n21211), .Z(n25469) );
  BUF_X1 U20851 ( .A(n21210), .Z(n25472) );
  BUF_X1 U20852 ( .A(n21209), .Z(n25475) );
  BUF_X1 U20853 ( .A(n21208), .Z(n25478) );
  BUF_X1 U20854 ( .A(n21207), .Z(n25481) );
  BUF_X1 U20855 ( .A(n21206), .Z(n25484) );
  BUF_X1 U20856 ( .A(n21205), .Z(n25487) );
  BUF_X1 U20857 ( .A(n21204), .Z(n25490) );
  BUF_X1 U20858 ( .A(n21203), .Z(n25493) );
  BUF_X1 U20859 ( .A(n21202), .Z(n25496) );
  BUF_X1 U20860 ( .A(n21201), .Z(n25499) );
  BUF_X1 U20861 ( .A(n21200), .Z(n25502) );
  BUF_X1 U20862 ( .A(n21199), .Z(n25505) );
  BUF_X1 U20863 ( .A(n21198), .Z(n25508) );
  BUF_X1 U20864 ( .A(n21197), .Z(n25511) );
  BUF_X1 U20865 ( .A(n21196), .Z(n25514) );
  BUF_X1 U20866 ( .A(n21195), .Z(n25517) );
  BUF_X1 U20867 ( .A(n21194), .Z(n25520) );
  BUF_X1 U20868 ( .A(n21193), .Z(n25523) );
  BUF_X1 U20869 ( .A(n21192), .Z(n25526) );
  BUF_X1 U20870 ( .A(n21191), .Z(n25529) );
  BUF_X1 U20871 ( .A(n21190), .Z(n25532) );
  BUF_X1 U20872 ( .A(n21188), .Z(n25552) );
  BUF_X1 U20873 ( .A(n21252), .Z(n25345) );
  BUF_X1 U20874 ( .A(n21251), .Z(n25348) );
  BUF_X1 U20875 ( .A(n21250), .Z(n25351) );
  BUF_X1 U20876 ( .A(n21249), .Z(n25354) );
  BUF_X1 U20877 ( .A(n21248), .Z(n25357) );
  BUF_X1 U20878 ( .A(n21247), .Z(n25360) );
  BUF_X1 U20879 ( .A(n21246), .Z(n25363) );
  BUF_X1 U20880 ( .A(n21245), .Z(n25366) );
  BUF_X1 U20881 ( .A(n21244), .Z(n25369) );
  BUF_X1 U20882 ( .A(n21243), .Z(n25372) );
  BUF_X1 U20883 ( .A(n21242), .Z(n25375) );
  BUF_X1 U20884 ( .A(n21241), .Z(n25378) );
  BUF_X1 U20885 ( .A(n21240), .Z(n25381) );
  BUF_X1 U20886 ( .A(n21239), .Z(n25384) );
  BUF_X1 U20887 ( .A(n21238), .Z(n25387) );
  BUF_X1 U20888 ( .A(n21237), .Z(n25390) );
  BUF_X1 U20889 ( .A(n21236), .Z(n25393) );
  BUF_X1 U20890 ( .A(n21235), .Z(n25396) );
  BUF_X1 U20891 ( .A(n21234), .Z(n25399) );
  BUF_X1 U20892 ( .A(n21233), .Z(n25402) );
  BUF_X1 U20893 ( .A(n21232), .Z(n25405) );
  BUF_X1 U20894 ( .A(n21231), .Z(n25408) );
  BUF_X1 U20895 ( .A(n21230), .Z(n25411) );
  BUF_X1 U20896 ( .A(n21229), .Z(n25414) );
  BUF_X1 U20897 ( .A(n21228), .Z(n25417) );
  BUF_X1 U20898 ( .A(n21227), .Z(n25420) );
  BUF_X1 U20899 ( .A(n21226), .Z(n25423) );
  BUF_X1 U20900 ( .A(n21225), .Z(n25426) );
  BUF_X1 U20901 ( .A(n21224), .Z(n25429) );
  BUF_X1 U20902 ( .A(n21223), .Z(n25432) );
  BUF_X1 U20903 ( .A(n21222), .Z(n25435) );
  BUF_X1 U20904 ( .A(n21221), .Z(n25438) );
  BUF_X1 U20905 ( .A(n21220), .Z(n25441) );
  BUF_X1 U20906 ( .A(n21219), .Z(n25444) );
  BUF_X1 U20907 ( .A(n21218), .Z(n25447) );
  BUF_X1 U20908 ( .A(n21217), .Z(n25450) );
  BUF_X1 U20909 ( .A(n21216), .Z(n25453) );
  BUF_X1 U20910 ( .A(n21215), .Z(n25456) );
  BUF_X1 U20911 ( .A(n21214), .Z(n25459) );
  BUF_X1 U20912 ( .A(n21213), .Z(n25462) );
  BUF_X1 U20913 ( .A(n21212), .Z(n25465) );
  BUF_X1 U20914 ( .A(n21211), .Z(n25468) );
  BUF_X1 U20915 ( .A(n21210), .Z(n25471) );
  BUF_X1 U20916 ( .A(n21209), .Z(n25474) );
  BUF_X1 U20917 ( .A(n21208), .Z(n25477) );
  BUF_X1 U20918 ( .A(n21207), .Z(n25480) );
  BUF_X1 U20919 ( .A(n21206), .Z(n25483) );
  BUF_X1 U20920 ( .A(n21205), .Z(n25486) );
  BUF_X1 U20921 ( .A(n21204), .Z(n25489) );
  BUF_X1 U20922 ( .A(n21203), .Z(n25492) );
  BUF_X1 U20923 ( .A(n21202), .Z(n25495) );
  BUF_X1 U20924 ( .A(n21201), .Z(n25498) );
  BUF_X1 U20925 ( .A(n21200), .Z(n25501) );
  BUF_X1 U20926 ( .A(n21199), .Z(n25504) );
  BUF_X1 U20927 ( .A(n21198), .Z(n25507) );
  BUF_X1 U20928 ( .A(n21197), .Z(n25510) );
  BUF_X1 U20929 ( .A(n21196), .Z(n25513) );
  BUF_X1 U20930 ( .A(n21195), .Z(n25516) );
  BUF_X1 U20931 ( .A(n21194), .Z(n25519) );
  BUF_X1 U20932 ( .A(n21193), .Z(n25522) );
  BUF_X1 U20933 ( .A(n21192), .Z(n25525) );
  BUF_X1 U20934 ( .A(n21191), .Z(n25528) );
  BUF_X1 U20935 ( .A(n21190), .Z(n25531) );
  BUF_X1 U20936 ( .A(n21188), .Z(n25551) );
  NAND2_X1 U20937 ( .A1(n22554), .A2(n22538), .ZN(n21334) );
  NAND2_X1 U20938 ( .A1(n22539), .A2(n22538), .ZN(n21310) );
  NAND2_X1 U20939 ( .A1(n22537), .A2(n22538), .ZN(n21311) );
  NAND2_X1 U20940 ( .A1(n22546), .A2(n22538), .ZN(n21320) );
  NAND2_X1 U20941 ( .A1(n22545), .A2(n22538), .ZN(n21321) );
  NAND2_X1 U20942 ( .A1(n23756), .A2(n23757), .ZN(n22593) );
  NAND2_X1 U20943 ( .A1(n23754), .A2(n23757), .ZN(n22595) );
  NAND2_X1 U20944 ( .A1(n23754), .A2(n23758), .ZN(n22596) );
  NAND2_X1 U20945 ( .A1(n23756), .A2(n23755), .ZN(n22597) );
  NAND2_X1 U20946 ( .A1(n22538), .A2(n22553), .ZN(n21335) );
  NAND2_X1 U20947 ( .A1(n23740), .A2(n23741), .ZN(n22569) );
  NAND2_X1 U20948 ( .A1(n23747), .A2(n23738), .ZN(n22579) );
  NAND2_X1 U20949 ( .A1(n22558), .A2(n22540), .ZN(n21344) );
  NAND2_X1 U20950 ( .A1(n22557), .A2(n22540), .ZN(n21345) );
  NAND2_X1 U20951 ( .A1(n22558), .A2(n22543), .ZN(n21349) );
  NAND2_X1 U20952 ( .A1(n22557), .A2(n22543), .ZN(n21350) );
  NAND2_X1 U20953 ( .A1(n23740), .A2(n23745), .ZN(n22611) );
  NAND2_X1 U20954 ( .A1(n23740), .A2(n23742), .ZN(n22605) );
  NAND2_X1 U20955 ( .A1(n23737), .A2(n23745), .ZN(n22606) );
  NAND2_X1 U20956 ( .A1(n22539), .A2(n22542), .ZN(n21315) );
  NAND2_X1 U20957 ( .A1(n22537), .A2(n22542), .ZN(n21316) );
  NAND2_X1 U20958 ( .A1(n22546), .A2(n22542), .ZN(n21325) );
  NAND2_X1 U20959 ( .A1(n22545), .A2(n22542), .ZN(n21326) );
  BUF_X1 U20960 ( .A(n22608), .Z(n24408) );
  BUF_X1 U20961 ( .A(n21297), .Z(n24804) );
  BUF_X1 U20962 ( .A(n21192), .Z(n25527) );
  BUF_X1 U20963 ( .A(n21191), .Z(n25530) );
  BUF_X1 U20964 ( .A(n21190), .Z(n25533) );
  BUF_X1 U20965 ( .A(n21188), .Z(n25553) );
  BUF_X1 U20966 ( .A(n21252), .Z(n25347) );
  BUF_X1 U20967 ( .A(n21251), .Z(n25350) );
  BUF_X1 U20968 ( .A(n21250), .Z(n25353) );
  BUF_X1 U20969 ( .A(n21249), .Z(n25356) );
  BUF_X1 U20970 ( .A(n21248), .Z(n25359) );
  BUF_X1 U20971 ( .A(n21247), .Z(n25362) );
  BUF_X1 U20972 ( .A(n21246), .Z(n25365) );
  BUF_X1 U20973 ( .A(n21245), .Z(n25368) );
  BUF_X1 U20974 ( .A(n21244), .Z(n25371) );
  BUF_X1 U20975 ( .A(n21243), .Z(n25374) );
  BUF_X1 U20976 ( .A(n21242), .Z(n25377) );
  BUF_X1 U20977 ( .A(n21241), .Z(n25380) );
  BUF_X1 U20978 ( .A(n21240), .Z(n25383) );
  BUF_X1 U20979 ( .A(n21239), .Z(n25386) );
  BUF_X1 U20980 ( .A(n21238), .Z(n25389) );
  BUF_X1 U20981 ( .A(n21237), .Z(n25392) );
  BUF_X1 U20982 ( .A(n21236), .Z(n25395) );
  BUF_X1 U20983 ( .A(n21235), .Z(n25398) );
  BUF_X1 U20984 ( .A(n21234), .Z(n25401) );
  BUF_X1 U20985 ( .A(n21233), .Z(n25404) );
  BUF_X1 U20986 ( .A(n21232), .Z(n25407) );
  BUF_X1 U20987 ( .A(n21231), .Z(n25410) );
  BUF_X1 U20988 ( .A(n21230), .Z(n25413) );
  BUF_X1 U20989 ( .A(n21229), .Z(n25416) );
  BUF_X1 U20990 ( .A(n21228), .Z(n25419) );
  BUF_X1 U20991 ( .A(n21227), .Z(n25422) );
  BUF_X1 U20992 ( .A(n21226), .Z(n25425) );
  BUF_X1 U20993 ( .A(n21225), .Z(n25428) );
  BUF_X1 U20994 ( .A(n21224), .Z(n25431) );
  BUF_X1 U20995 ( .A(n21223), .Z(n25434) );
  BUF_X1 U20996 ( .A(n21222), .Z(n25437) );
  BUF_X1 U20997 ( .A(n21221), .Z(n25440) );
  BUF_X1 U20998 ( .A(n21220), .Z(n25443) );
  BUF_X1 U20999 ( .A(n21219), .Z(n25446) );
  BUF_X1 U21000 ( .A(n21218), .Z(n25449) );
  BUF_X1 U21001 ( .A(n21217), .Z(n25452) );
  BUF_X1 U21002 ( .A(n21216), .Z(n25455) );
  BUF_X1 U21003 ( .A(n21215), .Z(n25458) );
  BUF_X1 U21004 ( .A(n21214), .Z(n25461) );
  BUF_X1 U21005 ( .A(n21213), .Z(n25464) );
  BUF_X1 U21006 ( .A(n21212), .Z(n25467) );
  BUF_X1 U21007 ( .A(n21211), .Z(n25470) );
  BUF_X1 U21008 ( .A(n21210), .Z(n25473) );
  BUF_X1 U21009 ( .A(n21209), .Z(n25476) );
  BUF_X1 U21010 ( .A(n21208), .Z(n25479) );
  BUF_X1 U21011 ( .A(n21207), .Z(n25482) );
  BUF_X1 U21012 ( .A(n21206), .Z(n25485) );
  BUF_X1 U21013 ( .A(n21205), .Z(n25488) );
  BUF_X1 U21014 ( .A(n21204), .Z(n25491) );
  BUF_X1 U21015 ( .A(n21203), .Z(n25494) );
  BUF_X1 U21016 ( .A(n21202), .Z(n25497) );
  BUF_X1 U21017 ( .A(n21201), .Z(n25500) );
  BUF_X1 U21018 ( .A(n21200), .Z(n25503) );
  BUF_X1 U21019 ( .A(n21199), .Z(n25506) );
  BUF_X1 U21020 ( .A(n21198), .Z(n25509) );
  BUF_X1 U21021 ( .A(n21197), .Z(n25512) );
  BUF_X1 U21022 ( .A(n21196), .Z(n25515) );
  BUF_X1 U21023 ( .A(n21195), .Z(n25518) );
  BUF_X1 U21024 ( .A(n21194), .Z(n25521) );
  BUF_X1 U21025 ( .A(n21193), .Z(n25524) );
  OAI21_X1 U21026 ( .B1(n21268), .B2(n21289), .A(n25564), .ZN(n21296) );
  NAND2_X1 U21027 ( .A1(n23745), .A2(n23744), .ZN(n22573) );
  AND2_X1 U21028 ( .A1(n23758), .A2(n23761), .ZN(n23740) );
  NAND2_X1 U21029 ( .A1(n23742), .A2(n23737), .ZN(n22568) );
  AND2_X1 U21030 ( .A1(n23761), .A2(n23757), .ZN(n23744) );
  AND2_X1 U21031 ( .A1(n23755), .A2(n23761), .ZN(n23737) );
  AND2_X1 U21032 ( .A1(n23759), .A2(n23761), .ZN(n23747) );
  NAND2_X1 U21033 ( .A1(n23737), .A2(n23748), .ZN(n22583) );
  NAND2_X1 U21034 ( .A1(n23740), .A2(n23748), .ZN(n22578) );
  AND2_X1 U21035 ( .A1(n23760), .A2(n19203), .ZN(n23754) );
  OR2_X1 U21036 ( .A1(n24413), .A2(n19190), .ZN(n22598) );
  NAND2_X1 U21037 ( .A1(n23754), .A2(n23759), .ZN(n22601) );
  NAND2_X1 U21038 ( .A1(n23756), .A2(n23758), .ZN(n22599) );
  NAND2_X1 U21039 ( .A1(n23756), .A2(n23759), .ZN(n22600) );
  AND2_X1 U21040 ( .A1(n23748), .A2(n23747), .ZN(n22586) );
  AND2_X1 U21041 ( .A1(n23745), .A2(n23747), .ZN(n22588) );
  AND2_X1 U21042 ( .A1(n23742), .A2(n23744), .ZN(n22582) );
  AND2_X1 U21043 ( .A1(n22543), .A2(n22554), .ZN(n21336) );
  AND2_X1 U21044 ( .A1(n22543), .A2(n22553), .ZN(n21337) );
  AND2_X1 U21045 ( .A1(n22558), .A2(n22542), .ZN(n21346) );
  AND2_X1 U21046 ( .A1(n22557), .A2(n22542), .ZN(n21347) );
  AND2_X1 U21047 ( .A1(n22558), .A2(n22538), .ZN(n21341) );
  AND2_X1 U21048 ( .A1(n22557), .A2(n22538), .ZN(n21342) );
  AND2_X1 U21049 ( .A1(n23738), .A2(n23744), .ZN(n22587) );
  AND2_X1 U21050 ( .A1(n23741), .A2(n23744), .ZN(n22576) );
  AND2_X1 U21051 ( .A1(n23741), .A2(n23747), .ZN(n22581) );
  AND2_X1 U21052 ( .A1(n23741), .A2(n23737), .ZN(n22607) );
  AND2_X1 U21053 ( .A1(n24803), .A2(n19190), .ZN(n21302) );
  AND2_X1 U21054 ( .A1(n22540), .A2(n22553), .ZN(n21332) );
  AND2_X1 U21055 ( .A1(n22539), .A2(n22543), .ZN(n21312) );
  AND2_X1 U21056 ( .A1(n22537), .A2(n22543), .ZN(n21313) );
  AND2_X1 U21057 ( .A1(n22546), .A2(n22543), .ZN(n21322) );
  AND2_X1 U21058 ( .A1(n22545), .A2(n22543), .ZN(n21323) );
  AND2_X1 U21059 ( .A1(n22540), .A2(n22554), .ZN(n21331) );
  AND2_X1 U21060 ( .A1(n23737), .A2(n23738), .ZN(n22572) );
  AND2_X1 U21061 ( .A1(n23740), .A2(n23738), .ZN(n22603) );
  AND2_X1 U21062 ( .A1(n22539), .A2(n22540), .ZN(n21307) );
  AND2_X1 U21063 ( .A1(n22537), .A2(n22540), .ZN(n21308) );
  AND2_X1 U21064 ( .A1(n22546), .A2(n22540), .ZN(n21317) );
  AND2_X1 U21065 ( .A1(n22545), .A2(n22540), .ZN(n21318) );
  AND3_X1 U21066 ( .A1(n19200), .A2(n19199), .A3(n23761), .ZN(n23760) );
  BUF_X1 U21067 ( .A(n21267), .Z(n25225) );
  OAI21_X1 U21068 ( .B1(n21253), .B2(n21268), .A(n25564), .ZN(n21267) );
  BUF_X1 U21069 ( .A(n21265), .Z(n25242) );
  OAI21_X1 U21070 ( .B1(n21253), .B2(n21266), .A(n25564), .ZN(n21265) );
  BUF_X1 U21071 ( .A(n21257), .Z(n25310) );
  OAI21_X1 U21072 ( .B1(n21253), .B2(n21258), .A(n25564), .ZN(n21257) );
  BUF_X1 U21073 ( .A(n21259), .Z(n25293) );
  OAI21_X1 U21074 ( .B1(n21253), .B2(n21260), .A(n25564), .ZN(n21259) );
  BUF_X1 U21075 ( .A(n21255), .Z(n25327) );
  OAI21_X1 U21076 ( .B1(n21253), .B2(n21256), .A(n25564), .ZN(n21255) );
  BUF_X1 U21077 ( .A(n21263), .Z(n25259) );
  OAI21_X1 U21078 ( .B1(n21253), .B2(n21264), .A(n25564), .ZN(n21263) );
  BUF_X1 U21079 ( .A(n21261), .Z(n25276) );
  OAI21_X1 U21080 ( .B1(n21253), .B2(n21262), .A(n25564), .ZN(n21261) );
  BUF_X1 U21081 ( .A(n21285), .Z(n24987) );
  OAI21_X1 U21082 ( .B1(n21264), .B2(n21280), .A(n25563), .ZN(n21285) );
  BUF_X1 U21083 ( .A(n21270), .Z(n25208) );
  OAI21_X1 U21084 ( .B1(n21254), .B2(n21271), .A(n25564), .ZN(n21270) );
  BUF_X1 U21085 ( .A(n21275), .Z(n25140) );
  OAI21_X1 U21086 ( .B1(n21262), .B2(n21271), .A(n25563), .ZN(n21275) );
  BUF_X1 U21087 ( .A(n21292), .Z(n24885) );
  OAI21_X1 U21088 ( .B1(n21260), .B2(n21289), .A(n25562), .ZN(n21292) );
  BUF_X1 U21089 ( .A(n21279), .Z(n25072) );
  OAI21_X1 U21090 ( .B1(n21254), .B2(n21280), .A(n25563), .ZN(n21279) );
  BUF_X1 U21091 ( .A(n21284), .Z(n25004) );
  OAI21_X1 U21092 ( .B1(n21262), .B2(n21280), .A(n25563), .ZN(n21284) );
  BUF_X1 U21093 ( .A(n21291), .Z(n24902) );
  OAI21_X1 U21094 ( .B1(n21258), .B2(n21289), .A(n25562), .ZN(n21291) );
  BUF_X1 U21095 ( .A(n21295), .Z(n24834) );
  OAI21_X1 U21096 ( .B1(n21266), .B2(n21289), .A(n25562), .ZN(n21295) );
  BUF_X1 U21097 ( .A(n21281), .Z(n25055) );
  OAI21_X1 U21098 ( .B1(n21256), .B2(n21280), .A(n25563), .ZN(n21281) );
  BUF_X1 U21099 ( .A(n21272), .Z(n25191) );
  OAI21_X1 U21100 ( .B1(n21256), .B2(n21271), .A(n25564), .ZN(n21272) );
  BUF_X1 U21101 ( .A(n21273), .Z(n25174) );
  OAI21_X1 U21102 ( .B1(n21258), .B2(n21271), .A(n25563), .ZN(n21273) );
  BUF_X1 U21103 ( .A(n21278), .Z(n25089) );
  OAI21_X1 U21104 ( .B1(n21268), .B2(n21271), .A(n25563), .ZN(n21278) );
  BUF_X1 U21105 ( .A(n21282), .Z(n25038) );
  OAI21_X1 U21106 ( .B1(n21258), .B2(n21280), .A(n25563), .ZN(n21282) );
  BUF_X1 U21107 ( .A(n21283), .Z(n25021) );
  OAI21_X1 U21108 ( .B1(n21260), .B2(n21280), .A(n25563), .ZN(n21283) );
  BUF_X1 U21109 ( .A(n21294), .Z(n24851) );
  OAI21_X1 U21110 ( .B1(n21264), .B2(n21289), .A(n25562), .ZN(n21294) );
  BUF_X1 U21111 ( .A(n21293), .Z(n24868) );
  OAI21_X1 U21112 ( .B1(n21262), .B2(n21289), .A(n25562), .ZN(n21293) );
  BUF_X1 U21113 ( .A(n21290), .Z(n24919) );
  OAI21_X1 U21114 ( .B1(n21256), .B2(n21289), .A(n25562), .ZN(n21290) );
  BUF_X1 U21115 ( .A(n21288), .Z(n24936) );
  OAI21_X1 U21116 ( .B1(n21254), .B2(n21289), .A(n25562), .ZN(n21288) );
  BUF_X1 U21117 ( .A(n21287), .Z(n24953) );
  OAI21_X1 U21118 ( .B1(n21268), .B2(n21280), .A(n25562), .ZN(n21287) );
  BUF_X1 U21119 ( .A(n21286), .Z(n24970) );
  OAI21_X1 U21120 ( .B1(n21266), .B2(n21280), .A(n25563), .ZN(n21286) );
  BUF_X1 U21121 ( .A(n21277), .Z(n25106) );
  OAI21_X1 U21122 ( .B1(n21266), .B2(n21271), .A(n25563), .ZN(n21277) );
  BUF_X1 U21123 ( .A(n21276), .Z(n25123) );
  OAI21_X1 U21124 ( .B1(n21264), .B2(n21271), .A(n25563), .ZN(n21276) );
  BUF_X1 U21125 ( .A(n21274), .Z(n25157) );
  OAI21_X1 U21126 ( .B1(n21260), .B2(n21271), .A(n25563), .ZN(n21274) );
  AOI222_X1 U21127 ( .A1(n24513), .A2(n24008), .B1(n24507), .B2(n8629), .C1(
        n24501), .C2(n8501), .ZN(n23019) );
  AOI222_X1 U21128 ( .A1(n24513), .A2(n24009), .B1(n24507), .B2(n8628), .C1(
        n24501), .C2(n8500), .ZN(n23001) );
  AOI222_X1 U21129 ( .A1(n24513), .A2(n24010), .B1(n24507), .B2(n8627), .C1(
        n24501), .C2(n8499), .ZN(n22983) );
  AOI222_X1 U21130 ( .A1(n24513), .A2(n24011), .B1(n24507), .B2(n8626), .C1(
        n24501), .C2(n8498), .ZN(n22965) );
  AOI222_X1 U21131 ( .A1(n24513), .A2(n24012), .B1(n24507), .B2(n8625), .C1(
        n24501), .C2(n8497), .ZN(n22947) );
  AOI222_X1 U21132 ( .A1(n24513), .A2(n24013), .B1(n24507), .B2(n8624), .C1(
        n24501), .C2(n8496), .ZN(n22929) );
  AOI222_X1 U21133 ( .A1(n24513), .A2(n24014), .B1(n24507), .B2(n8623), .C1(
        n24501), .C2(n8495), .ZN(n22911) );
  AOI222_X1 U21134 ( .A1(n24513), .A2(n24015), .B1(n24507), .B2(n8622), .C1(
        n24501), .C2(n8494), .ZN(n22893) );
  AOI222_X1 U21135 ( .A1(n24514), .A2(n24016), .B1(n24508), .B2(n8621), .C1(
        n24502), .C2(n8493), .ZN(n22875) );
  AOI222_X1 U21136 ( .A1(n24514), .A2(n24017), .B1(n24508), .B2(n8620), .C1(
        n24502), .C2(n8492), .ZN(n22857) );
  AOI222_X1 U21137 ( .A1(n24514), .A2(n24018), .B1(n24508), .B2(n8619), .C1(
        n24502), .C2(n8491), .ZN(n22839) );
  AOI222_X1 U21138 ( .A1(n24514), .A2(n24019), .B1(n24508), .B2(n8618), .C1(
        n24502), .C2(n8490), .ZN(n22821) );
  AOI222_X1 U21139 ( .A1(n24514), .A2(n24020), .B1(n24508), .B2(n8617), .C1(
        n24502), .C2(n8489), .ZN(n22803) );
  AOI222_X1 U21140 ( .A1(n24514), .A2(n24021), .B1(n24508), .B2(n8616), .C1(
        n24502), .C2(n8488), .ZN(n22785) );
  AOI222_X1 U21141 ( .A1(n24514), .A2(n24022), .B1(n24508), .B2(n8615), .C1(
        n24502), .C2(n8487), .ZN(n22767) );
  AOI222_X1 U21142 ( .A1(n24514), .A2(n24023), .B1(n24508), .B2(n8614), .C1(
        n24502), .C2(n8486), .ZN(n22749) );
  AOI222_X1 U21143 ( .A1(n24514), .A2(n24024), .B1(n24508), .B2(n8613), .C1(
        n24502), .C2(n8485), .ZN(n22731) );
  AOI222_X1 U21144 ( .A1(n24514), .A2(n24025), .B1(n24508), .B2(n8612), .C1(
        n24502), .C2(n8484), .ZN(n22713) );
  AOI222_X1 U21145 ( .A1(n24514), .A2(n24026), .B1(n24508), .B2(n8611), .C1(
        n24502), .C2(n8483), .ZN(n22695) );
  AOI222_X1 U21146 ( .A1(n24514), .A2(n24027), .B1(n24508), .B2(n8610), .C1(
        n24502), .C2(n8482), .ZN(n22677) );
  AOI222_X1 U21147 ( .A1(n24515), .A2(n24028), .B1(n24509), .B2(n8609), .C1(
        n24503), .C2(n8481), .ZN(n22659) );
  AOI222_X1 U21148 ( .A1(n24515), .A2(n24029), .B1(n24509), .B2(n8608), .C1(
        n24503), .C2(n8480), .ZN(n22641) );
  AOI222_X1 U21149 ( .A1(n24515), .A2(n24030), .B1(n24509), .B2(n8607), .C1(
        n24503), .C2(n8479), .ZN(n22623) );
  AOI222_X1 U21150 ( .A1(n24515), .A2(n24031), .B1(n24509), .B2(n8606), .C1(
        n24503), .C2(n8478), .ZN(n22585) );
  AOI222_X1 U21151 ( .A1(n24510), .A2(n23968), .B1(n24504), .B2(n8669), .C1(
        n24498), .C2(n8541), .ZN(n23749) );
  AOI222_X1 U21152 ( .A1(n24510), .A2(n23969), .B1(n24504), .B2(n8668), .C1(
        n24498), .C2(n8540), .ZN(n23721) );
  AOI222_X1 U21153 ( .A1(n24510), .A2(n23970), .B1(n24504), .B2(n8667), .C1(
        n24498), .C2(n8539), .ZN(n23703) );
  AOI222_X1 U21154 ( .A1(n24510), .A2(n23971), .B1(n24504), .B2(n8666), .C1(
        n24498), .C2(n8538), .ZN(n23685) );
  AOI222_X1 U21155 ( .A1(n24510), .A2(n23972), .B1(n24504), .B2(n8665), .C1(
        n24498), .C2(n8537), .ZN(n23667) );
  AOI222_X1 U21156 ( .A1(n24510), .A2(n23973), .B1(n24504), .B2(n8664), .C1(
        n24498), .C2(n8536), .ZN(n23649) );
  AOI222_X1 U21157 ( .A1(n24510), .A2(n23974), .B1(n24504), .B2(n8663), .C1(
        n24498), .C2(n8535), .ZN(n23631) );
  AOI222_X1 U21158 ( .A1(n24510), .A2(n23975), .B1(n24504), .B2(n8662), .C1(
        n24498), .C2(n8534), .ZN(n23613) );
  AOI222_X1 U21159 ( .A1(n24510), .A2(n23976), .B1(n24504), .B2(n8661), .C1(
        n24498), .C2(n8533), .ZN(n23595) );
  AOI222_X1 U21160 ( .A1(n24510), .A2(n23977), .B1(n24504), .B2(n8660), .C1(
        n24498), .C2(n8532), .ZN(n23577) );
  AOI222_X1 U21161 ( .A1(n24510), .A2(n23978), .B1(n24504), .B2(n8659), .C1(
        n24498), .C2(n8531), .ZN(n23559) );
  AOI222_X1 U21162 ( .A1(n24510), .A2(n23979), .B1(n24504), .B2(n8658), .C1(
        n24498), .C2(n8530), .ZN(n23541) );
  AOI222_X1 U21163 ( .A1(n24511), .A2(n23980), .B1(n24505), .B2(n8657), .C1(
        n24499), .C2(n8529), .ZN(n23523) );
  AOI222_X1 U21164 ( .A1(n24511), .A2(n23981), .B1(n24505), .B2(n8656), .C1(
        n24499), .C2(n8528), .ZN(n23505) );
  AOI222_X1 U21165 ( .A1(n24511), .A2(n23982), .B1(n24505), .B2(n8655), .C1(
        n24499), .C2(n8527), .ZN(n23487) );
  AOI222_X1 U21166 ( .A1(n24511), .A2(n23983), .B1(n24505), .B2(n8654), .C1(
        n24499), .C2(n8526), .ZN(n23469) );
  AOI222_X1 U21167 ( .A1(n24511), .A2(n23984), .B1(n24505), .B2(n8653), .C1(
        n24499), .C2(n8525), .ZN(n23451) );
  AOI222_X1 U21168 ( .A1(n24511), .A2(n23985), .B1(n24505), .B2(n8652), .C1(
        n24499), .C2(n8524), .ZN(n23433) );
  AOI222_X1 U21169 ( .A1(n24511), .A2(n23986), .B1(n24505), .B2(n8651), .C1(
        n24499), .C2(n8523), .ZN(n23415) );
  AOI222_X1 U21170 ( .A1(n24511), .A2(n23987), .B1(n24505), .B2(n8650), .C1(
        n24499), .C2(n8522), .ZN(n23397) );
  AOI222_X1 U21171 ( .A1(n24511), .A2(n23988), .B1(n24505), .B2(n8649), .C1(
        n24499), .C2(n8521), .ZN(n23379) );
  AOI222_X1 U21172 ( .A1(n24511), .A2(n23989), .B1(n24505), .B2(n8648), .C1(
        n24499), .C2(n8520), .ZN(n23361) );
  AOI222_X1 U21173 ( .A1(n24511), .A2(n23990), .B1(n24505), .B2(n8647), .C1(
        n24499), .C2(n8519), .ZN(n23343) );
  AOI222_X1 U21174 ( .A1(n24511), .A2(n23991), .B1(n24505), .B2(n8646), .C1(
        n24499), .C2(n8518), .ZN(n23325) );
  AOI222_X1 U21175 ( .A1(n24512), .A2(n23992), .B1(n24506), .B2(n8645), .C1(
        n24500), .C2(n8517), .ZN(n23307) );
  AOI222_X1 U21176 ( .A1(n24512), .A2(n23993), .B1(n24506), .B2(n8644), .C1(
        n24500), .C2(n8516), .ZN(n23289) );
  AOI222_X1 U21177 ( .A1(n24512), .A2(n23994), .B1(n24506), .B2(n8643), .C1(
        n24500), .C2(n8515), .ZN(n23271) );
  AOI222_X1 U21178 ( .A1(n24512), .A2(n23995), .B1(n24506), .B2(n8642), .C1(
        n24500), .C2(n8514), .ZN(n23253) );
  AOI222_X1 U21179 ( .A1(n24512), .A2(n23996), .B1(n24506), .B2(n8641), .C1(
        n24500), .C2(n8513), .ZN(n23235) );
  AOI222_X1 U21180 ( .A1(n24512), .A2(n23997), .B1(n24506), .B2(n8640), .C1(
        n24500), .C2(n8512), .ZN(n23217) );
  AOI222_X1 U21181 ( .A1(n24512), .A2(n23998), .B1(n24506), .B2(n8639), .C1(
        n24500), .C2(n8511), .ZN(n23199) );
  AOI222_X1 U21182 ( .A1(n24512), .A2(n23999), .B1(n24506), .B2(n8638), .C1(
        n24500), .C2(n8510), .ZN(n23181) );
  AOI222_X1 U21183 ( .A1(n24512), .A2(n24000), .B1(n24506), .B2(n8637), .C1(
        n24500), .C2(n8509), .ZN(n23163) );
  AOI222_X1 U21184 ( .A1(n24512), .A2(n24001), .B1(n24506), .B2(n8636), .C1(
        n24500), .C2(n8508), .ZN(n23145) );
  AOI222_X1 U21185 ( .A1(n24512), .A2(n24002), .B1(n24506), .B2(n8635), .C1(
        n24500), .C2(n8507), .ZN(n23127) );
  AOI222_X1 U21186 ( .A1(n24512), .A2(n24003), .B1(n24506), .B2(n8634), .C1(
        n24500), .C2(n8506), .ZN(n23109) );
  AOI222_X1 U21187 ( .A1(n24513), .A2(n24004), .B1(n24507), .B2(n8633), .C1(
        n24501), .C2(n8505), .ZN(n23091) );
  AOI222_X1 U21188 ( .A1(n24513), .A2(n24005), .B1(n24507), .B2(n8632), .C1(
        n24501), .C2(n8504), .ZN(n23073) );
  AOI222_X1 U21189 ( .A1(n24513), .A2(n24006), .B1(n24507), .B2(n8631), .C1(
        n24501), .C2(n8503), .ZN(n23055) );
  AOI222_X1 U21190 ( .A1(n24513), .A2(n24007), .B1(n24507), .B2(n8630), .C1(
        n24501), .C2(n8502), .ZN(n23037) );
  OAI222_X1 U21191 ( .A1(n20285), .A2(n24459), .B1(n17290), .B2(n24453), .C1(
        n19355), .C2(n24447), .ZN(n23020) );
  OAI222_X1 U21192 ( .A1(n20284), .A2(n24459), .B1(n17287), .B2(n24453), .C1(
        n19354), .C2(n24447), .ZN(n23002) );
  OAI222_X1 U21193 ( .A1(n20283), .A2(n24459), .B1(n17284), .B2(n24453), .C1(
        n19353), .C2(n24447), .ZN(n22984) );
  OAI222_X1 U21194 ( .A1(n20282), .A2(n24459), .B1(n17281), .B2(n24453), .C1(
        n19352), .C2(n24447), .ZN(n22966) );
  OAI222_X1 U21195 ( .A1(n20281), .A2(n24459), .B1(n17278), .B2(n24453), .C1(
        n19351), .C2(n24447), .ZN(n22948) );
  OAI222_X1 U21196 ( .A1(n20280), .A2(n24459), .B1(n17275), .B2(n24453), .C1(
        n19350), .C2(n24447), .ZN(n22930) );
  OAI222_X1 U21197 ( .A1(n20279), .A2(n24459), .B1(n17272), .B2(n24453), .C1(
        n19349), .C2(n24447), .ZN(n22912) );
  OAI222_X1 U21198 ( .A1(n20278), .A2(n24459), .B1(n17269), .B2(n24453), .C1(
        n19348), .C2(n24447), .ZN(n22894) );
  OAI222_X1 U21199 ( .A1(n20277), .A2(n24460), .B1(n17266), .B2(n24454), .C1(
        n19347), .C2(n24448), .ZN(n22876) );
  OAI222_X1 U21200 ( .A1(n20276), .A2(n24460), .B1(n17263), .B2(n24454), .C1(
        n19346), .C2(n24448), .ZN(n22858) );
  OAI222_X1 U21201 ( .A1(n20275), .A2(n24460), .B1(n17260), .B2(n24454), .C1(
        n19345), .C2(n24448), .ZN(n22840) );
  OAI222_X1 U21202 ( .A1(n20274), .A2(n24460), .B1(n17257), .B2(n24454), .C1(
        n19344), .C2(n24448), .ZN(n22822) );
  OAI222_X1 U21203 ( .A1(n20273), .A2(n24460), .B1(n17254), .B2(n24454), .C1(
        n19343), .C2(n24448), .ZN(n22804) );
  OAI222_X1 U21204 ( .A1(n20272), .A2(n24460), .B1(n17251), .B2(n24454), .C1(
        n19342), .C2(n24448), .ZN(n22786) );
  OAI222_X1 U21205 ( .A1(n20271), .A2(n24460), .B1(n17248), .B2(n24454), .C1(
        n19341), .C2(n24448), .ZN(n22768) );
  OAI222_X1 U21206 ( .A1(n20270), .A2(n24460), .B1(n17245), .B2(n24454), .C1(
        n19340), .C2(n24448), .ZN(n22750) );
  OAI222_X1 U21207 ( .A1(n20269), .A2(n24460), .B1(n17242), .B2(n24454), .C1(
        n19339), .C2(n24448), .ZN(n22732) );
  OAI222_X1 U21208 ( .A1(n20268), .A2(n24460), .B1(n17239), .B2(n24454), .C1(
        n19338), .C2(n24448), .ZN(n22714) );
  OAI222_X1 U21209 ( .A1(n20267), .A2(n24460), .B1(n17236), .B2(n24454), .C1(
        n19337), .C2(n24448), .ZN(n22696) );
  OAI222_X1 U21210 ( .A1(n20266), .A2(n24460), .B1(n17233), .B2(n24454), .C1(
        n19336), .C2(n24448), .ZN(n22678) );
  OAI222_X1 U21211 ( .A1(n20397), .A2(n24456), .B1(n17410), .B2(n24450), .C1(
        n19395), .C2(n24444), .ZN(n23750) );
  OAI222_X1 U21212 ( .A1(n20396), .A2(n24456), .B1(n17407), .B2(n24450), .C1(
        n19394), .C2(n24444), .ZN(n23722) );
  OAI222_X1 U21213 ( .A1(n20395), .A2(n24456), .B1(n17404), .B2(n24450), .C1(
        n19393), .C2(n24444), .ZN(n23704) );
  OAI222_X1 U21214 ( .A1(n20394), .A2(n24456), .B1(n17401), .B2(n24450), .C1(
        n19392), .C2(n24444), .ZN(n23686) );
  OAI222_X1 U21215 ( .A1(n20393), .A2(n24456), .B1(n17398), .B2(n24450), .C1(
        n19391), .C2(n24444), .ZN(n23668) );
  OAI222_X1 U21216 ( .A1(n20392), .A2(n24456), .B1(n17395), .B2(n24450), .C1(
        n19390), .C2(n24444), .ZN(n23650) );
  OAI222_X1 U21217 ( .A1(n20391), .A2(n24456), .B1(n17392), .B2(n24450), .C1(
        n19389), .C2(n24444), .ZN(n23632) );
  OAI222_X1 U21218 ( .A1(n20390), .A2(n24456), .B1(n17389), .B2(n24450), .C1(
        n19388), .C2(n24444), .ZN(n23614) );
  OAI222_X1 U21219 ( .A1(n20389), .A2(n24456), .B1(n17386), .B2(n24450), .C1(
        n19387), .C2(n24444), .ZN(n23596) );
  OAI222_X1 U21220 ( .A1(n20388), .A2(n24456), .B1(n17383), .B2(n24450), .C1(
        n19386), .C2(n24444), .ZN(n23578) );
  OAI222_X1 U21221 ( .A1(n20387), .A2(n24456), .B1(n17380), .B2(n24450), .C1(
        n19385), .C2(n24444), .ZN(n23560) );
  OAI222_X1 U21222 ( .A1(n20386), .A2(n24456), .B1(n17377), .B2(n24450), .C1(
        n19384), .C2(n24444), .ZN(n23542) );
  OAI222_X1 U21223 ( .A1(n20385), .A2(n24457), .B1(n17374), .B2(n24451), .C1(
        n19383), .C2(n24445), .ZN(n23524) );
  OAI222_X1 U21224 ( .A1(n20384), .A2(n24457), .B1(n17371), .B2(n24451), .C1(
        n19382), .C2(n24445), .ZN(n23506) );
  OAI222_X1 U21225 ( .A1(n20383), .A2(n24457), .B1(n17368), .B2(n24451), .C1(
        n19381), .C2(n24445), .ZN(n23488) );
  OAI222_X1 U21226 ( .A1(n20382), .A2(n24457), .B1(n17365), .B2(n24451), .C1(
        n19380), .C2(n24445), .ZN(n23470) );
  OAI222_X1 U21227 ( .A1(n20381), .A2(n24457), .B1(n17362), .B2(n24451), .C1(
        n19379), .C2(n24445), .ZN(n23452) );
  OAI222_X1 U21228 ( .A1(n20380), .A2(n24457), .B1(n17359), .B2(n24451), .C1(
        n19378), .C2(n24445), .ZN(n23434) );
  OAI222_X1 U21229 ( .A1(n20379), .A2(n24457), .B1(n17356), .B2(n24451), .C1(
        n19377), .C2(n24445), .ZN(n23416) );
  OAI222_X1 U21230 ( .A1(n20378), .A2(n24457), .B1(n17353), .B2(n24451), .C1(
        n19376), .C2(n24445), .ZN(n23398) );
  OAI222_X1 U21231 ( .A1(n20377), .A2(n24457), .B1(n17350), .B2(n24451), .C1(
        n19375), .C2(n24445), .ZN(n23380) );
  OAI222_X1 U21232 ( .A1(n20376), .A2(n24457), .B1(n17347), .B2(n24451), .C1(
        n19374), .C2(n24445), .ZN(n23362) );
  OAI222_X1 U21233 ( .A1(n20375), .A2(n24457), .B1(n17344), .B2(n24451), .C1(
        n19373), .C2(n24445), .ZN(n23344) );
  OAI222_X1 U21234 ( .A1(n20374), .A2(n24457), .B1(n17341), .B2(n24451), .C1(
        n19372), .C2(n24445), .ZN(n23326) );
  OAI222_X1 U21235 ( .A1(n20301), .A2(n24458), .B1(n17338), .B2(n24452), .C1(
        n19371), .C2(n24446), .ZN(n23308) );
  OAI222_X1 U21236 ( .A1(n20300), .A2(n24458), .B1(n17335), .B2(n24452), .C1(
        n19370), .C2(n24446), .ZN(n23290) );
  OAI222_X1 U21237 ( .A1(n20299), .A2(n24458), .B1(n17332), .B2(n24452), .C1(
        n19369), .C2(n24446), .ZN(n23272) );
  OAI222_X1 U21238 ( .A1(n20298), .A2(n24458), .B1(n17329), .B2(n24452), .C1(
        n19368), .C2(n24446), .ZN(n23254) );
  OAI222_X1 U21239 ( .A1(n20297), .A2(n24458), .B1(n17326), .B2(n24452), .C1(
        n19367), .C2(n24446), .ZN(n23236) );
  OAI222_X1 U21240 ( .A1(n20296), .A2(n24458), .B1(n17323), .B2(n24452), .C1(
        n19366), .C2(n24446), .ZN(n23218) );
  OAI222_X1 U21241 ( .A1(n20295), .A2(n24458), .B1(n17320), .B2(n24452), .C1(
        n19365), .C2(n24446), .ZN(n23200) );
  OAI222_X1 U21242 ( .A1(n20294), .A2(n24458), .B1(n17317), .B2(n24452), .C1(
        n19364), .C2(n24446), .ZN(n23182) );
  OAI222_X1 U21243 ( .A1(n20293), .A2(n24458), .B1(n17314), .B2(n24452), .C1(
        n19363), .C2(n24446), .ZN(n23164) );
  OAI222_X1 U21244 ( .A1(n20292), .A2(n24458), .B1(n17311), .B2(n24452), .C1(
        n19362), .C2(n24446), .ZN(n23146) );
  OAI222_X1 U21245 ( .A1(n20291), .A2(n24458), .B1(n17308), .B2(n24452), .C1(
        n19361), .C2(n24446), .ZN(n23128) );
  OAI222_X1 U21246 ( .A1(n20290), .A2(n24458), .B1(n17305), .B2(n24452), .C1(
        n19360), .C2(n24446), .ZN(n23110) );
  OAI222_X1 U21247 ( .A1(n20289), .A2(n24459), .B1(n17302), .B2(n24453), .C1(
        n19359), .C2(n24447), .ZN(n23092) );
  OAI222_X1 U21248 ( .A1(n20288), .A2(n24459), .B1(n17299), .B2(n24453), .C1(
        n19358), .C2(n24447), .ZN(n23074) );
  OAI222_X1 U21249 ( .A1(n20287), .A2(n24459), .B1(n17296), .B2(n24453), .C1(
        n19357), .C2(n24447), .ZN(n23056) );
  OAI222_X1 U21250 ( .A1(n20286), .A2(n24459), .B1(n17293), .B2(n24453), .C1(
        n19356), .C2(n24447), .ZN(n23038) );
  OAI222_X1 U21251 ( .A1(n20253), .A2(n24461), .B1(n17230), .B2(n24455), .C1(
        n19335), .C2(n24449), .ZN(n22660) );
  OAI222_X1 U21252 ( .A1(n20252), .A2(n24461), .B1(n17227), .B2(n24455), .C1(
        n19334), .C2(n24449), .ZN(n22642) );
  OAI222_X1 U21253 ( .A1(n20251), .A2(n24461), .B1(n17224), .B2(n24455), .C1(
        n19333), .C2(n24449), .ZN(n22624) );
  OAI222_X1 U21254 ( .A1(n20250), .A2(n24461), .B1(n17221), .B2(n24455), .C1(
        n19332), .C2(n24449), .ZN(n22589) );
  NOR4_X1 U21255 ( .A1(n22652), .A2(n22653), .A3(n22654), .A4(n22655), .ZN(
        n22651) );
  OAI221_X1 U21256 ( .B1(n20513), .B2(n24551), .C1(n20517), .C2(n24545), .A(
        n22658), .ZN(n22653) );
  OAI221_X1 U21257 ( .B1(n20265), .B2(n24575), .C1(n7307), .C2(n24569), .A(
        n22657), .ZN(n22654) );
  OAI221_X1 U21258 ( .B1(n20509), .B2(n24527), .C1(n836), .C2(n24521), .A(
        n22659), .ZN(n22652) );
  NOR4_X1 U21259 ( .A1(n22634), .A2(n22635), .A3(n22636), .A4(n22637), .ZN(
        n22633) );
  OAI221_X1 U21260 ( .B1(n20512), .B2(n24551), .C1(n20516), .C2(n24545), .A(
        n22640), .ZN(n22635) );
  OAI221_X1 U21261 ( .B1(n20264), .B2(n24575), .C1(n7305), .C2(n24569), .A(
        n22639), .ZN(n22636) );
  OAI221_X1 U21262 ( .B1(n20508), .B2(n24527), .C1(n835), .C2(n24521), .A(
        n22641), .ZN(n22634) );
  NOR4_X1 U21263 ( .A1(n22616), .A2(n22617), .A3(n22618), .A4(n22619), .ZN(
        n22615) );
  OAI221_X1 U21264 ( .B1(n20511), .B2(n24551), .C1(n20515), .C2(n24545), .A(
        n22622), .ZN(n22617) );
  OAI221_X1 U21265 ( .B1(n20263), .B2(n24575), .C1(n7303), .C2(n24569), .A(
        n22621), .ZN(n22618) );
  OAI221_X1 U21266 ( .B1(n20507), .B2(n24527), .C1(n834), .C2(n24521), .A(
        n22623), .ZN(n22616) );
  NOR4_X1 U21267 ( .A1(n22564), .A2(n22565), .A3(n22566), .A4(n22567), .ZN(
        n22563) );
  OAI221_X1 U21268 ( .B1(n20510), .B2(n24551), .C1(n20514), .C2(n24545), .A(
        n22580), .ZN(n22565) );
  OAI221_X1 U21269 ( .B1(n20262), .B2(n24575), .C1(n7301), .C2(n24569), .A(
        n22575), .ZN(n22566) );
  OAI221_X1 U21270 ( .B1(n20506), .B2(n24527), .C1(n833), .C2(n24521), .A(
        n22585), .ZN(n22564) );
  NOR4_X1 U21271 ( .A1(n23012), .A2(n23013), .A3(n23014), .A4(n23015), .ZN(
        n23011) );
  OAI221_X1 U21272 ( .B1(n20602), .B2(n24549), .C1(n20638), .C2(n24543), .A(
        n23018), .ZN(n23013) );
  OAI221_X1 U21273 ( .B1(n20465), .B2(n24573), .C1(n7347), .C2(n24567), .A(
        n23017), .ZN(n23014) );
  OAI221_X1 U21274 ( .B1(n20566), .B2(n24525), .C1(n856), .C2(n24519), .A(
        n23019), .ZN(n23012) );
  NOR4_X1 U21275 ( .A1(n22994), .A2(n22995), .A3(n22996), .A4(n22997), .ZN(
        n22993) );
  OAI221_X1 U21276 ( .B1(n20601), .B2(n24549), .C1(n20637), .C2(n24543), .A(
        n23000), .ZN(n22995) );
  OAI221_X1 U21277 ( .B1(n20464), .B2(n24573), .C1(n7345), .C2(n24567), .A(
        n22999), .ZN(n22996) );
  OAI221_X1 U21278 ( .B1(n20565), .B2(n24525), .C1(n855), .C2(n24519), .A(
        n23001), .ZN(n22994) );
  NOR4_X1 U21279 ( .A1(n22976), .A2(n22977), .A3(n22978), .A4(n22979), .ZN(
        n22975) );
  OAI221_X1 U21280 ( .B1(n20600), .B2(n24549), .C1(n20636), .C2(n24543), .A(
        n22982), .ZN(n22977) );
  OAI221_X1 U21281 ( .B1(n20463), .B2(n24573), .C1(n7343), .C2(n24567), .A(
        n22981), .ZN(n22978) );
  OAI221_X1 U21282 ( .B1(n20564), .B2(n24525), .C1(n854), .C2(n24519), .A(
        n22983), .ZN(n22976) );
  NOR4_X1 U21283 ( .A1(n22958), .A2(n22959), .A3(n22960), .A4(n22961), .ZN(
        n22957) );
  OAI221_X1 U21284 ( .B1(n20599), .B2(n24549), .C1(n20635), .C2(n24543), .A(
        n22964), .ZN(n22959) );
  OAI221_X1 U21285 ( .B1(n20462), .B2(n24573), .C1(n7341), .C2(n24567), .A(
        n22963), .ZN(n22960) );
  OAI221_X1 U21286 ( .B1(n20563), .B2(n24525), .C1(n853), .C2(n24519), .A(
        n22965), .ZN(n22958) );
  NOR4_X1 U21287 ( .A1(n22940), .A2(n22941), .A3(n22942), .A4(n22943), .ZN(
        n22939) );
  OAI221_X1 U21288 ( .B1(n20598), .B2(n24549), .C1(n20634), .C2(n24543), .A(
        n22946), .ZN(n22941) );
  OAI221_X1 U21289 ( .B1(n20461), .B2(n24573), .C1(n7339), .C2(n24567), .A(
        n22945), .ZN(n22942) );
  OAI221_X1 U21290 ( .B1(n20562), .B2(n24525), .C1(n852), .C2(n24519), .A(
        n22947), .ZN(n22940) );
  NOR4_X1 U21291 ( .A1(n22922), .A2(n22923), .A3(n22924), .A4(n22925), .ZN(
        n22921) );
  OAI221_X1 U21292 ( .B1(n20597), .B2(n24549), .C1(n20633), .C2(n24543), .A(
        n22928), .ZN(n22923) );
  OAI221_X1 U21293 ( .B1(n20460), .B2(n24573), .C1(n7337), .C2(n24567), .A(
        n22927), .ZN(n22924) );
  OAI221_X1 U21294 ( .B1(n20561), .B2(n24525), .C1(n851), .C2(n24519), .A(
        n22929), .ZN(n22922) );
  NOR4_X1 U21295 ( .A1(n22904), .A2(n22905), .A3(n22906), .A4(n22907), .ZN(
        n22903) );
  OAI221_X1 U21296 ( .B1(n20596), .B2(n24549), .C1(n20632), .C2(n24543), .A(
        n22910), .ZN(n22905) );
  OAI221_X1 U21297 ( .B1(n20459), .B2(n24573), .C1(n7335), .C2(n24567), .A(
        n22909), .ZN(n22906) );
  OAI221_X1 U21298 ( .B1(n20560), .B2(n24525), .C1(n850), .C2(n24519), .A(
        n22911), .ZN(n22904) );
  NOR4_X1 U21299 ( .A1(n22886), .A2(n22887), .A3(n22888), .A4(n22889), .ZN(
        n22885) );
  OAI221_X1 U21300 ( .B1(n20595), .B2(n24549), .C1(n20631), .C2(n24543), .A(
        n22892), .ZN(n22887) );
  OAI221_X1 U21301 ( .B1(n20458), .B2(n24573), .C1(n7333), .C2(n24567), .A(
        n22891), .ZN(n22888) );
  OAI221_X1 U21302 ( .B1(n20559), .B2(n24525), .C1(n849), .C2(n24519), .A(
        n22893), .ZN(n22886) );
  NOR4_X1 U21303 ( .A1(n22868), .A2(n22869), .A3(n22870), .A4(n22871), .ZN(
        n22867) );
  OAI221_X1 U21304 ( .B1(n20594), .B2(n24550), .C1(n20630), .C2(n24544), .A(
        n22874), .ZN(n22869) );
  OAI221_X1 U21305 ( .B1(n20457), .B2(n24574), .C1(n7331), .C2(n24568), .A(
        n22873), .ZN(n22870) );
  OAI221_X1 U21306 ( .B1(n20558), .B2(n24526), .C1(n848), .C2(n24520), .A(
        n22875), .ZN(n22868) );
  NOR4_X1 U21307 ( .A1(n22850), .A2(n22851), .A3(n22852), .A4(n22853), .ZN(
        n22849) );
  OAI221_X1 U21308 ( .B1(n20593), .B2(n24550), .C1(n20629), .C2(n24544), .A(
        n22856), .ZN(n22851) );
  OAI221_X1 U21309 ( .B1(n20456), .B2(n24574), .C1(n7329), .C2(n24568), .A(
        n22855), .ZN(n22852) );
  OAI221_X1 U21310 ( .B1(n20557), .B2(n24526), .C1(n847), .C2(n24520), .A(
        n22857), .ZN(n22850) );
  NOR4_X1 U21311 ( .A1(n22832), .A2(n22833), .A3(n22834), .A4(n22835), .ZN(
        n22831) );
  OAI221_X1 U21312 ( .B1(n20592), .B2(n24550), .C1(n20628), .C2(n24544), .A(
        n22838), .ZN(n22833) );
  OAI221_X1 U21313 ( .B1(n20455), .B2(n24574), .C1(n7327), .C2(n24568), .A(
        n22837), .ZN(n22834) );
  OAI221_X1 U21314 ( .B1(n20556), .B2(n24526), .C1(n846), .C2(n24520), .A(
        n22839), .ZN(n22832) );
  NOR4_X1 U21315 ( .A1(n22814), .A2(n22815), .A3(n22816), .A4(n22817), .ZN(
        n22813) );
  OAI221_X1 U21316 ( .B1(n20591), .B2(n24550), .C1(n20627), .C2(n24544), .A(
        n22820), .ZN(n22815) );
  OAI221_X1 U21317 ( .B1(n20454), .B2(n24574), .C1(n7325), .C2(n24568), .A(
        n22819), .ZN(n22816) );
  OAI221_X1 U21318 ( .B1(n20555), .B2(n24526), .C1(n845), .C2(n24520), .A(
        n22821), .ZN(n22814) );
  NOR4_X1 U21319 ( .A1(n22796), .A2(n22797), .A3(n22798), .A4(n22799), .ZN(
        n22795) );
  OAI221_X1 U21320 ( .B1(n20590), .B2(n24550), .C1(n20626), .C2(n24544), .A(
        n22802), .ZN(n22797) );
  OAI221_X1 U21321 ( .B1(n20453), .B2(n24574), .C1(n7323), .C2(n24568), .A(
        n22801), .ZN(n22798) );
  OAI221_X1 U21322 ( .B1(n20554), .B2(n24526), .C1(n844), .C2(n24520), .A(
        n22803), .ZN(n22796) );
  NOR4_X1 U21323 ( .A1(n22778), .A2(n22779), .A3(n22780), .A4(n22781), .ZN(
        n22777) );
  OAI221_X1 U21324 ( .B1(n20589), .B2(n24550), .C1(n20625), .C2(n24544), .A(
        n22784), .ZN(n22779) );
  OAI221_X1 U21325 ( .B1(n20452), .B2(n24574), .C1(n7321), .C2(n24568), .A(
        n22783), .ZN(n22780) );
  OAI221_X1 U21326 ( .B1(n20553), .B2(n24526), .C1(n843), .C2(n24520), .A(
        n22785), .ZN(n22778) );
  NOR4_X1 U21327 ( .A1(n22760), .A2(n22761), .A3(n22762), .A4(n22763), .ZN(
        n22759) );
  OAI221_X1 U21328 ( .B1(n20588), .B2(n24550), .C1(n20624), .C2(n24544), .A(
        n22766), .ZN(n22761) );
  OAI221_X1 U21329 ( .B1(n20451), .B2(n24574), .C1(n7319), .C2(n24568), .A(
        n22765), .ZN(n22762) );
  OAI221_X1 U21330 ( .B1(n20552), .B2(n24526), .C1(n842), .C2(n24520), .A(
        n22767), .ZN(n22760) );
  NOR4_X1 U21331 ( .A1(n22742), .A2(n22743), .A3(n22744), .A4(n22745), .ZN(
        n22741) );
  OAI221_X1 U21332 ( .B1(n20587), .B2(n24550), .C1(n20623), .C2(n24544), .A(
        n22748), .ZN(n22743) );
  OAI221_X1 U21333 ( .B1(n20450), .B2(n24574), .C1(n7317), .C2(n24568), .A(
        n22747), .ZN(n22744) );
  OAI221_X1 U21334 ( .B1(n20551), .B2(n24526), .C1(n841), .C2(n24520), .A(
        n22749), .ZN(n22742) );
  NOR4_X1 U21335 ( .A1(n22724), .A2(n22725), .A3(n22726), .A4(n22727), .ZN(
        n22723) );
  OAI221_X1 U21336 ( .B1(n20586), .B2(n24550), .C1(n20622), .C2(n24544), .A(
        n22730), .ZN(n22725) );
  OAI221_X1 U21337 ( .B1(n20449), .B2(n24574), .C1(n7315), .C2(n24568), .A(
        n22729), .ZN(n22726) );
  OAI221_X1 U21338 ( .B1(n20550), .B2(n24526), .C1(n840), .C2(n24520), .A(
        n22731), .ZN(n22724) );
  NOR4_X1 U21339 ( .A1(n22706), .A2(n22707), .A3(n22708), .A4(n22709), .ZN(
        n22705) );
  OAI221_X1 U21340 ( .B1(n20585), .B2(n24550), .C1(n20621), .C2(n24544), .A(
        n22712), .ZN(n22707) );
  OAI221_X1 U21341 ( .B1(n20448), .B2(n24574), .C1(n7313), .C2(n24568), .A(
        n22711), .ZN(n22708) );
  OAI221_X1 U21342 ( .B1(n20549), .B2(n24526), .C1(n839), .C2(n24520), .A(
        n22713), .ZN(n22706) );
  NOR4_X1 U21343 ( .A1(n22688), .A2(n22689), .A3(n22690), .A4(n22691), .ZN(
        n22687) );
  OAI221_X1 U21344 ( .B1(n20584), .B2(n24550), .C1(n20620), .C2(n24544), .A(
        n22694), .ZN(n22689) );
  OAI221_X1 U21345 ( .B1(n20447), .B2(n24574), .C1(n7311), .C2(n24568), .A(
        n22693), .ZN(n22690) );
  OAI221_X1 U21346 ( .B1(n20548), .B2(n24526), .C1(n838), .C2(n24520), .A(
        n22695), .ZN(n22688) );
  NOR4_X1 U21347 ( .A1(n22670), .A2(n22671), .A3(n22672), .A4(n22673), .ZN(
        n22669) );
  OAI221_X1 U21348 ( .B1(n20583), .B2(n24550), .C1(n20619), .C2(n24544), .A(
        n22676), .ZN(n22671) );
  OAI221_X1 U21349 ( .B1(n20446), .B2(n24574), .C1(n7309), .C2(n24568), .A(
        n22675), .ZN(n22672) );
  OAI221_X1 U21350 ( .B1(n20547), .B2(n24526), .C1(n837), .C2(n24520), .A(
        n22677), .ZN(n22670) );
  NOR4_X1 U21351 ( .A1(n23732), .A2(n23733), .A3(n23734), .A4(n23735), .ZN(
        n23731) );
  OAI221_X1 U21352 ( .B1(n20774), .B2(n24546), .C1(n20798), .C2(n24540), .A(
        n23746), .ZN(n23733) );
  OAI221_X1 U21353 ( .B1(n20505), .B2(n24570), .C1(n7427), .C2(n24564), .A(
        n23743), .ZN(n23734) );
  OAI221_X1 U21354 ( .B1(n20750), .B2(n24522), .C1(n896), .C2(n24516), .A(
        n23749), .ZN(n23732) );
  NOR4_X1 U21355 ( .A1(n23714), .A2(n23715), .A3(n23716), .A4(n23717), .ZN(
        n23713) );
  OAI221_X1 U21356 ( .B1(n20773), .B2(n24546), .C1(n20797), .C2(n24540), .A(
        n23720), .ZN(n23715) );
  OAI221_X1 U21357 ( .B1(n20504), .B2(n24570), .C1(n7425), .C2(n24564), .A(
        n23719), .ZN(n23716) );
  OAI221_X1 U21358 ( .B1(n20749), .B2(n24522), .C1(n895), .C2(n24516), .A(
        n23721), .ZN(n23714) );
  NOR4_X1 U21359 ( .A1(n23696), .A2(n23697), .A3(n23698), .A4(n23699), .ZN(
        n23695) );
  OAI221_X1 U21360 ( .B1(n20772), .B2(n24546), .C1(n20796), .C2(n24540), .A(
        n23702), .ZN(n23697) );
  OAI221_X1 U21361 ( .B1(n20503), .B2(n24570), .C1(n7423), .C2(n24564), .A(
        n23701), .ZN(n23698) );
  OAI221_X1 U21362 ( .B1(n20748), .B2(n24522), .C1(n894), .C2(n24516), .A(
        n23703), .ZN(n23696) );
  NOR4_X1 U21363 ( .A1(n23678), .A2(n23679), .A3(n23680), .A4(n23681), .ZN(
        n23677) );
  OAI221_X1 U21364 ( .B1(n20771), .B2(n24546), .C1(n20795), .C2(n24540), .A(
        n23684), .ZN(n23679) );
  OAI221_X1 U21365 ( .B1(n20502), .B2(n24570), .C1(n7421), .C2(n24564), .A(
        n23683), .ZN(n23680) );
  OAI221_X1 U21366 ( .B1(n20747), .B2(n24522), .C1(n893), .C2(n24516), .A(
        n23685), .ZN(n23678) );
  NOR4_X1 U21367 ( .A1(n23660), .A2(n23661), .A3(n23662), .A4(n23663), .ZN(
        n23659) );
  OAI221_X1 U21368 ( .B1(n20770), .B2(n24546), .C1(n20794), .C2(n24540), .A(
        n23666), .ZN(n23661) );
  OAI221_X1 U21369 ( .B1(n20501), .B2(n24570), .C1(n7419), .C2(n24564), .A(
        n23665), .ZN(n23662) );
  OAI221_X1 U21370 ( .B1(n20746), .B2(n24522), .C1(n892), .C2(n24516), .A(
        n23667), .ZN(n23660) );
  NOR4_X1 U21371 ( .A1(n23642), .A2(n23643), .A3(n23644), .A4(n23645), .ZN(
        n23641) );
  OAI221_X1 U21372 ( .B1(n20769), .B2(n24546), .C1(n20793), .C2(n24540), .A(
        n23648), .ZN(n23643) );
  OAI221_X1 U21373 ( .B1(n20500), .B2(n24570), .C1(n7417), .C2(n24564), .A(
        n23647), .ZN(n23644) );
  OAI221_X1 U21374 ( .B1(n20745), .B2(n24522), .C1(n891), .C2(n24516), .A(
        n23649), .ZN(n23642) );
  NOR4_X1 U21375 ( .A1(n23624), .A2(n23625), .A3(n23626), .A4(n23627), .ZN(
        n23623) );
  OAI221_X1 U21376 ( .B1(n20768), .B2(n24546), .C1(n20792), .C2(n24540), .A(
        n23630), .ZN(n23625) );
  OAI221_X1 U21377 ( .B1(n20499), .B2(n24570), .C1(n7415), .C2(n24564), .A(
        n23629), .ZN(n23626) );
  OAI221_X1 U21378 ( .B1(n20744), .B2(n24522), .C1(n890), .C2(n24516), .A(
        n23631), .ZN(n23624) );
  NOR4_X1 U21379 ( .A1(n23606), .A2(n23607), .A3(n23608), .A4(n23609), .ZN(
        n23605) );
  OAI221_X1 U21380 ( .B1(n20767), .B2(n24546), .C1(n20791), .C2(n24540), .A(
        n23612), .ZN(n23607) );
  OAI221_X1 U21381 ( .B1(n20498), .B2(n24570), .C1(n7413), .C2(n24564), .A(
        n23611), .ZN(n23608) );
  OAI221_X1 U21382 ( .B1(n20743), .B2(n24522), .C1(n889), .C2(n24516), .A(
        n23613), .ZN(n23606) );
  NOR4_X1 U21383 ( .A1(n23588), .A2(n23589), .A3(n23590), .A4(n23591), .ZN(
        n23587) );
  OAI221_X1 U21384 ( .B1(n20766), .B2(n24546), .C1(n20790), .C2(n24540), .A(
        n23594), .ZN(n23589) );
  OAI221_X1 U21385 ( .B1(n20497), .B2(n24570), .C1(n7411), .C2(n24564), .A(
        n23593), .ZN(n23590) );
  OAI221_X1 U21386 ( .B1(n20742), .B2(n24522), .C1(n888), .C2(n24516), .A(
        n23595), .ZN(n23588) );
  NOR4_X1 U21387 ( .A1(n23570), .A2(n23571), .A3(n23572), .A4(n23573), .ZN(
        n23569) );
  OAI221_X1 U21388 ( .B1(n20765), .B2(n24546), .C1(n20789), .C2(n24540), .A(
        n23576), .ZN(n23571) );
  OAI221_X1 U21389 ( .B1(n20496), .B2(n24570), .C1(n7409), .C2(n24564), .A(
        n23575), .ZN(n23572) );
  OAI221_X1 U21390 ( .B1(n20741), .B2(n24522), .C1(n887), .C2(n24516), .A(
        n23577), .ZN(n23570) );
  NOR4_X1 U21391 ( .A1(n23552), .A2(n23553), .A3(n23554), .A4(n23555), .ZN(
        n23551) );
  OAI221_X1 U21392 ( .B1(n20764), .B2(n24546), .C1(n20788), .C2(n24540), .A(
        n23558), .ZN(n23553) );
  OAI221_X1 U21393 ( .B1(n20495), .B2(n24570), .C1(n7407), .C2(n24564), .A(
        n23557), .ZN(n23554) );
  OAI221_X1 U21394 ( .B1(n20740), .B2(n24522), .C1(n886), .C2(n24516), .A(
        n23559), .ZN(n23552) );
  NOR4_X1 U21395 ( .A1(n23534), .A2(n23535), .A3(n23536), .A4(n23537), .ZN(
        n23533) );
  OAI221_X1 U21396 ( .B1(n20763), .B2(n24546), .C1(n20787), .C2(n24540), .A(
        n23540), .ZN(n23535) );
  OAI221_X1 U21397 ( .B1(n20494), .B2(n24570), .C1(n7405), .C2(n24564), .A(
        n23539), .ZN(n23536) );
  OAI221_X1 U21398 ( .B1(n20739), .B2(n24522), .C1(n885), .C2(n24516), .A(
        n23541), .ZN(n23534) );
  NOR4_X1 U21399 ( .A1(n23516), .A2(n23517), .A3(n23518), .A4(n23519), .ZN(
        n23515) );
  OAI221_X1 U21400 ( .B1(n20762), .B2(n24547), .C1(n20786), .C2(n24541), .A(
        n23522), .ZN(n23517) );
  OAI221_X1 U21401 ( .B1(n20493), .B2(n24571), .C1(n7403), .C2(n24565), .A(
        n23521), .ZN(n23518) );
  OAI221_X1 U21402 ( .B1(n20738), .B2(n24523), .C1(n884), .C2(n24517), .A(
        n23523), .ZN(n23516) );
  NOR4_X1 U21403 ( .A1(n23498), .A2(n23499), .A3(n23500), .A4(n23501), .ZN(
        n23497) );
  OAI221_X1 U21404 ( .B1(n20761), .B2(n24547), .C1(n20785), .C2(n24541), .A(
        n23504), .ZN(n23499) );
  OAI221_X1 U21405 ( .B1(n20492), .B2(n24571), .C1(n7401), .C2(n24565), .A(
        n23503), .ZN(n23500) );
  OAI221_X1 U21406 ( .B1(n20737), .B2(n24523), .C1(n883), .C2(n24517), .A(
        n23505), .ZN(n23498) );
  NOR4_X1 U21407 ( .A1(n23480), .A2(n23481), .A3(n23482), .A4(n23483), .ZN(
        n23479) );
  OAI221_X1 U21408 ( .B1(n20760), .B2(n24547), .C1(n20784), .C2(n24541), .A(
        n23486), .ZN(n23481) );
  OAI221_X1 U21409 ( .B1(n20491), .B2(n24571), .C1(n7399), .C2(n24565), .A(
        n23485), .ZN(n23482) );
  OAI221_X1 U21410 ( .B1(n20736), .B2(n24523), .C1(n882), .C2(n24517), .A(
        n23487), .ZN(n23480) );
  NOR4_X1 U21411 ( .A1(n23462), .A2(n23463), .A3(n23464), .A4(n23465), .ZN(
        n23461) );
  OAI221_X1 U21412 ( .B1(n20759), .B2(n24547), .C1(n20783), .C2(n24541), .A(
        n23468), .ZN(n23463) );
  OAI221_X1 U21413 ( .B1(n20490), .B2(n24571), .C1(n7397), .C2(n24565), .A(
        n23467), .ZN(n23464) );
  OAI221_X1 U21414 ( .B1(n20735), .B2(n24523), .C1(n881), .C2(n24517), .A(
        n23469), .ZN(n23462) );
  NOR4_X1 U21415 ( .A1(n23444), .A2(n23445), .A3(n23446), .A4(n23447), .ZN(
        n23443) );
  OAI221_X1 U21416 ( .B1(n20758), .B2(n24547), .C1(n20782), .C2(n24541), .A(
        n23450), .ZN(n23445) );
  OAI221_X1 U21417 ( .B1(n20489), .B2(n24571), .C1(n7395), .C2(n24565), .A(
        n23449), .ZN(n23446) );
  OAI221_X1 U21418 ( .B1(n20734), .B2(n24523), .C1(n880), .C2(n24517), .A(
        n23451), .ZN(n23444) );
  NOR4_X1 U21419 ( .A1(n23426), .A2(n23427), .A3(n23428), .A4(n23429), .ZN(
        n23425) );
  OAI221_X1 U21420 ( .B1(n20757), .B2(n24547), .C1(n20781), .C2(n24541), .A(
        n23432), .ZN(n23427) );
  OAI221_X1 U21421 ( .B1(n20488), .B2(n24571), .C1(n7393), .C2(n24565), .A(
        n23431), .ZN(n23428) );
  OAI221_X1 U21422 ( .B1(n20733), .B2(n24523), .C1(n879), .C2(n24517), .A(
        n23433), .ZN(n23426) );
  NOR4_X1 U21423 ( .A1(n23408), .A2(n23409), .A3(n23410), .A4(n23411), .ZN(
        n23407) );
  OAI221_X1 U21424 ( .B1(n20756), .B2(n24547), .C1(n20780), .C2(n24541), .A(
        n23414), .ZN(n23409) );
  OAI221_X1 U21425 ( .B1(n20487), .B2(n24571), .C1(n7391), .C2(n24565), .A(
        n23413), .ZN(n23410) );
  OAI221_X1 U21426 ( .B1(n20732), .B2(n24523), .C1(n878), .C2(n24517), .A(
        n23415), .ZN(n23408) );
  NOR4_X1 U21427 ( .A1(n23390), .A2(n23391), .A3(n23392), .A4(n23393), .ZN(
        n23389) );
  OAI221_X1 U21428 ( .B1(n20755), .B2(n24547), .C1(n20779), .C2(n24541), .A(
        n23396), .ZN(n23391) );
  OAI221_X1 U21429 ( .B1(n20486), .B2(n24571), .C1(n7389), .C2(n24565), .A(
        n23395), .ZN(n23392) );
  OAI221_X1 U21430 ( .B1(n20731), .B2(n24523), .C1(n877), .C2(n24517), .A(
        n23397), .ZN(n23390) );
  NOR4_X1 U21431 ( .A1(n23372), .A2(n23373), .A3(n23374), .A4(n23375), .ZN(
        n23371) );
  OAI221_X1 U21432 ( .B1(n20754), .B2(n24547), .C1(n20778), .C2(n24541), .A(
        n23378), .ZN(n23373) );
  OAI221_X1 U21433 ( .B1(n20485), .B2(n24571), .C1(n7387), .C2(n24565), .A(
        n23377), .ZN(n23374) );
  OAI221_X1 U21434 ( .B1(n20730), .B2(n24523), .C1(n876), .C2(n24517), .A(
        n23379), .ZN(n23372) );
  NOR4_X1 U21435 ( .A1(n23354), .A2(n23355), .A3(n23356), .A4(n23357), .ZN(
        n23353) );
  OAI221_X1 U21436 ( .B1(n20753), .B2(n24547), .C1(n20777), .C2(n24541), .A(
        n23360), .ZN(n23355) );
  OAI221_X1 U21437 ( .B1(n20484), .B2(n24571), .C1(n7385), .C2(n24565), .A(
        n23359), .ZN(n23356) );
  OAI221_X1 U21438 ( .B1(n20729), .B2(n24523), .C1(n875), .C2(n24517), .A(
        n23361), .ZN(n23354) );
  NOR4_X1 U21439 ( .A1(n23336), .A2(n23337), .A3(n23338), .A4(n23339), .ZN(
        n23335) );
  OAI221_X1 U21440 ( .B1(n20752), .B2(n24547), .C1(n20776), .C2(n24541), .A(
        n23342), .ZN(n23337) );
  OAI221_X1 U21441 ( .B1(n20483), .B2(n24571), .C1(n7383), .C2(n24565), .A(
        n23341), .ZN(n23338) );
  OAI221_X1 U21442 ( .B1(n20728), .B2(n24523), .C1(n874), .C2(n24517), .A(
        n23343), .ZN(n23336) );
  NOR4_X1 U21443 ( .A1(n23318), .A2(n23319), .A3(n23320), .A4(n23321), .ZN(
        n23317) );
  OAI221_X1 U21444 ( .B1(n20751), .B2(n24547), .C1(n20775), .C2(n24541), .A(
        n23324), .ZN(n23319) );
  OAI221_X1 U21445 ( .B1(n20482), .B2(n24571), .C1(n7381), .C2(n24565), .A(
        n23323), .ZN(n23320) );
  OAI221_X1 U21446 ( .B1(n20727), .B2(n24523), .C1(n873), .C2(n24517), .A(
        n23325), .ZN(n23318) );
  NOR4_X1 U21447 ( .A1(n23300), .A2(n23301), .A3(n23302), .A4(n23303), .ZN(
        n23299) );
  OAI221_X1 U21448 ( .B1(n20618), .B2(n24548), .C1(n20654), .C2(n24542), .A(
        n23306), .ZN(n23301) );
  OAI221_X1 U21449 ( .B1(n20481), .B2(n24572), .C1(n7379), .C2(n24566), .A(
        n23305), .ZN(n23302) );
  OAI221_X1 U21450 ( .B1(n20582), .B2(n24524), .C1(n872), .C2(n24518), .A(
        n23307), .ZN(n23300) );
  NOR4_X1 U21451 ( .A1(n23282), .A2(n23283), .A3(n23284), .A4(n23285), .ZN(
        n23281) );
  OAI221_X1 U21452 ( .B1(n20617), .B2(n24548), .C1(n20653), .C2(n24542), .A(
        n23288), .ZN(n23283) );
  OAI221_X1 U21453 ( .B1(n20480), .B2(n24572), .C1(n7377), .C2(n24566), .A(
        n23287), .ZN(n23284) );
  OAI221_X1 U21454 ( .B1(n20581), .B2(n24524), .C1(n871), .C2(n24518), .A(
        n23289), .ZN(n23282) );
  NOR4_X1 U21455 ( .A1(n23264), .A2(n23265), .A3(n23266), .A4(n23267), .ZN(
        n23263) );
  OAI221_X1 U21456 ( .B1(n20616), .B2(n24548), .C1(n20652), .C2(n24542), .A(
        n23270), .ZN(n23265) );
  OAI221_X1 U21457 ( .B1(n20479), .B2(n24572), .C1(n7375), .C2(n24566), .A(
        n23269), .ZN(n23266) );
  OAI221_X1 U21458 ( .B1(n20580), .B2(n24524), .C1(n870), .C2(n24518), .A(
        n23271), .ZN(n23264) );
  NOR4_X1 U21459 ( .A1(n23246), .A2(n23247), .A3(n23248), .A4(n23249), .ZN(
        n23245) );
  OAI221_X1 U21460 ( .B1(n20615), .B2(n24548), .C1(n20651), .C2(n24542), .A(
        n23252), .ZN(n23247) );
  OAI221_X1 U21461 ( .B1(n20478), .B2(n24572), .C1(n7373), .C2(n24566), .A(
        n23251), .ZN(n23248) );
  OAI221_X1 U21462 ( .B1(n20579), .B2(n24524), .C1(n869), .C2(n24518), .A(
        n23253), .ZN(n23246) );
  NOR4_X1 U21463 ( .A1(n23228), .A2(n23229), .A3(n23230), .A4(n23231), .ZN(
        n23227) );
  OAI221_X1 U21464 ( .B1(n20614), .B2(n24548), .C1(n20650), .C2(n24542), .A(
        n23234), .ZN(n23229) );
  OAI221_X1 U21465 ( .B1(n20477), .B2(n24572), .C1(n7371), .C2(n24566), .A(
        n23233), .ZN(n23230) );
  OAI221_X1 U21466 ( .B1(n20578), .B2(n24524), .C1(n868), .C2(n24518), .A(
        n23235), .ZN(n23228) );
  NOR4_X1 U21467 ( .A1(n23210), .A2(n23211), .A3(n23212), .A4(n23213), .ZN(
        n23209) );
  OAI221_X1 U21468 ( .B1(n20613), .B2(n24548), .C1(n20649), .C2(n24542), .A(
        n23216), .ZN(n23211) );
  OAI221_X1 U21469 ( .B1(n20476), .B2(n24572), .C1(n7369), .C2(n24566), .A(
        n23215), .ZN(n23212) );
  OAI221_X1 U21470 ( .B1(n20577), .B2(n24524), .C1(n867), .C2(n24518), .A(
        n23217), .ZN(n23210) );
  NOR4_X1 U21471 ( .A1(n23192), .A2(n23193), .A3(n23194), .A4(n23195), .ZN(
        n23191) );
  OAI221_X1 U21472 ( .B1(n20612), .B2(n24548), .C1(n20648), .C2(n24542), .A(
        n23198), .ZN(n23193) );
  OAI221_X1 U21473 ( .B1(n20475), .B2(n24572), .C1(n7367), .C2(n24566), .A(
        n23197), .ZN(n23194) );
  OAI221_X1 U21474 ( .B1(n20576), .B2(n24524), .C1(n866), .C2(n24518), .A(
        n23199), .ZN(n23192) );
  NOR4_X1 U21475 ( .A1(n23174), .A2(n23175), .A3(n23176), .A4(n23177), .ZN(
        n23173) );
  OAI221_X1 U21476 ( .B1(n20611), .B2(n24548), .C1(n20647), .C2(n24542), .A(
        n23180), .ZN(n23175) );
  OAI221_X1 U21477 ( .B1(n20474), .B2(n24572), .C1(n7365), .C2(n24566), .A(
        n23179), .ZN(n23176) );
  OAI221_X1 U21478 ( .B1(n20575), .B2(n24524), .C1(n865), .C2(n24518), .A(
        n23181), .ZN(n23174) );
  NOR4_X1 U21479 ( .A1(n23156), .A2(n23157), .A3(n23158), .A4(n23159), .ZN(
        n23155) );
  OAI221_X1 U21480 ( .B1(n20610), .B2(n24548), .C1(n20646), .C2(n24542), .A(
        n23162), .ZN(n23157) );
  OAI221_X1 U21481 ( .B1(n20473), .B2(n24572), .C1(n7363), .C2(n24566), .A(
        n23161), .ZN(n23158) );
  OAI221_X1 U21482 ( .B1(n20574), .B2(n24524), .C1(n864), .C2(n24518), .A(
        n23163), .ZN(n23156) );
  NOR4_X1 U21483 ( .A1(n23138), .A2(n23139), .A3(n23140), .A4(n23141), .ZN(
        n23137) );
  OAI221_X1 U21484 ( .B1(n20609), .B2(n24548), .C1(n20645), .C2(n24542), .A(
        n23144), .ZN(n23139) );
  OAI221_X1 U21485 ( .B1(n20472), .B2(n24572), .C1(n7361), .C2(n24566), .A(
        n23143), .ZN(n23140) );
  OAI221_X1 U21486 ( .B1(n20573), .B2(n24524), .C1(n863), .C2(n24518), .A(
        n23145), .ZN(n23138) );
  NOR4_X1 U21487 ( .A1(n23120), .A2(n23121), .A3(n23122), .A4(n23123), .ZN(
        n23119) );
  OAI221_X1 U21488 ( .B1(n20608), .B2(n24548), .C1(n20644), .C2(n24542), .A(
        n23126), .ZN(n23121) );
  OAI221_X1 U21489 ( .B1(n20471), .B2(n24572), .C1(n7359), .C2(n24566), .A(
        n23125), .ZN(n23122) );
  OAI221_X1 U21490 ( .B1(n20572), .B2(n24524), .C1(n862), .C2(n24518), .A(
        n23127), .ZN(n23120) );
  NOR4_X1 U21491 ( .A1(n23102), .A2(n23103), .A3(n23104), .A4(n23105), .ZN(
        n23101) );
  OAI221_X1 U21492 ( .B1(n20607), .B2(n24548), .C1(n20643), .C2(n24542), .A(
        n23108), .ZN(n23103) );
  OAI221_X1 U21493 ( .B1(n20470), .B2(n24572), .C1(n7357), .C2(n24566), .A(
        n23107), .ZN(n23104) );
  OAI221_X1 U21494 ( .B1(n20571), .B2(n24524), .C1(n861), .C2(n24518), .A(
        n23109), .ZN(n23102) );
  NOR4_X1 U21495 ( .A1(n23084), .A2(n23085), .A3(n23086), .A4(n23087), .ZN(
        n23083) );
  OAI221_X1 U21496 ( .B1(n20606), .B2(n24549), .C1(n20642), .C2(n24543), .A(
        n23090), .ZN(n23085) );
  OAI221_X1 U21497 ( .B1(n20469), .B2(n24573), .C1(n7355), .C2(n24567), .A(
        n23089), .ZN(n23086) );
  OAI221_X1 U21498 ( .B1(n20570), .B2(n24525), .C1(n860), .C2(n24519), .A(
        n23091), .ZN(n23084) );
  NOR4_X1 U21499 ( .A1(n23066), .A2(n23067), .A3(n23068), .A4(n23069), .ZN(
        n23065) );
  OAI221_X1 U21500 ( .B1(n20605), .B2(n24549), .C1(n20641), .C2(n24543), .A(
        n23072), .ZN(n23067) );
  OAI221_X1 U21501 ( .B1(n20468), .B2(n24573), .C1(n7353), .C2(n24567), .A(
        n23071), .ZN(n23068) );
  OAI221_X1 U21502 ( .B1(n20569), .B2(n24525), .C1(n859), .C2(n24519), .A(
        n23073), .ZN(n23066) );
  NOR4_X1 U21503 ( .A1(n23048), .A2(n23049), .A3(n23050), .A4(n23051), .ZN(
        n23047) );
  OAI221_X1 U21504 ( .B1(n20604), .B2(n24549), .C1(n20640), .C2(n24543), .A(
        n23054), .ZN(n23049) );
  OAI221_X1 U21505 ( .B1(n20467), .B2(n24573), .C1(n7351), .C2(n24567), .A(
        n23053), .ZN(n23050) );
  OAI221_X1 U21506 ( .B1(n20568), .B2(n24525), .C1(n858), .C2(n24519), .A(
        n23055), .ZN(n23048) );
  NOR4_X1 U21507 ( .A1(n23030), .A2(n23031), .A3(n23032), .A4(n23033), .ZN(
        n23029) );
  OAI221_X1 U21508 ( .B1(n20603), .B2(n24549), .C1(n20639), .C2(n24543), .A(
        n23036), .ZN(n23031) );
  OAI221_X1 U21509 ( .B1(n20466), .B2(n24573), .C1(n7349), .C2(n24567), .A(
        n23035), .ZN(n23032) );
  OAI221_X1 U21510 ( .B1(n20567), .B2(n24525), .C1(n857), .C2(n24519), .A(
        n23037), .ZN(n23030) );
  AOI221_X1 U21511 ( .B1(n24786), .B2(n8285), .C1(n24780), .C2(n8733), .A(
        n22536), .ZN(n22535) );
  OAI22_X1 U21512 ( .A1(n8988), .A2(n24774), .B1(n19737), .B2(n24768), .ZN(
        n22536) );
  AOI221_X1 U21513 ( .B1(n24786), .B2(n8284), .C1(n24780), .C2(n8732), .A(
        n22517), .ZN(n22516) );
  OAI22_X1 U21514 ( .A1(n8986), .A2(n24774), .B1(n19736), .B2(n24768), .ZN(
        n22517) );
  AOI221_X1 U21515 ( .B1(n24786), .B2(n8283), .C1(n24780), .C2(n8731), .A(
        n22498), .ZN(n22497) );
  OAI22_X1 U21516 ( .A1(n8984), .A2(n24774), .B1(n19735), .B2(n24768), .ZN(
        n22498) );
  AOI221_X1 U21517 ( .B1(n24786), .B2(n8282), .C1(n24780), .C2(n8730), .A(
        n22479), .ZN(n22478) );
  OAI22_X1 U21518 ( .A1(n8982), .A2(n24774), .B1(n19734), .B2(n24768), .ZN(
        n22479) );
  AOI221_X1 U21519 ( .B1(n24786), .B2(n8281), .C1(n24780), .C2(n8729), .A(
        n22460), .ZN(n22459) );
  OAI22_X1 U21520 ( .A1(n8980), .A2(n24774), .B1(n19733), .B2(n24768), .ZN(
        n22460) );
  AOI221_X1 U21521 ( .B1(n24786), .B2(n8280), .C1(n24780), .C2(n8728), .A(
        n22441), .ZN(n22440) );
  OAI22_X1 U21522 ( .A1(n8978), .A2(n24774), .B1(n19732), .B2(n24768), .ZN(
        n22441) );
  AOI221_X1 U21523 ( .B1(n24786), .B2(n8279), .C1(n24780), .C2(n8727), .A(
        n22422), .ZN(n22421) );
  OAI22_X1 U21524 ( .A1(n8976), .A2(n24774), .B1(n19731), .B2(n24768), .ZN(
        n22422) );
  AOI221_X1 U21525 ( .B1(n24786), .B2(n8278), .C1(n24780), .C2(n8726), .A(
        n22403), .ZN(n22402) );
  OAI22_X1 U21526 ( .A1(n8974), .A2(n24774), .B1(n19730), .B2(n24768), .ZN(
        n22403) );
  AOI221_X1 U21527 ( .B1(n24786), .B2(n8277), .C1(n24780), .C2(n8725), .A(
        n22384), .ZN(n22383) );
  OAI22_X1 U21528 ( .A1(n8972), .A2(n24774), .B1(n19729), .B2(n24768), .ZN(
        n22384) );
  AOI221_X1 U21529 ( .B1(n24786), .B2(n8276), .C1(n24780), .C2(n8724), .A(
        n22365), .ZN(n22364) );
  OAI22_X1 U21530 ( .A1(n8970), .A2(n24774), .B1(n19728), .B2(n24768), .ZN(
        n22365) );
  AOI221_X1 U21531 ( .B1(n24786), .B2(n8275), .C1(n24780), .C2(n8723), .A(
        n22346), .ZN(n22345) );
  OAI22_X1 U21532 ( .A1(n8968), .A2(n24774), .B1(n19727), .B2(n24768), .ZN(
        n22346) );
  AOI221_X1 U21533 ( .B1(n24786), .B2(n8274), .C1(n24780), .C2(n8722), .A(
        n22327), .ZN(n22326) );
  OAI22_X1 U21534 ( .A1(n8966), .A2(n24774), .B1(n19726), .B2(n24768), .ZN(
        n22327) );
  AOI221_X1 U21535 ( .B1(n24787), .B2(n8273), .C1(n24781), .C2(n8721), .A(
        n22308), .ZN(n22307) );
  OAI22_X1 U21536 ( .A1(n8964), .A2(n24775), .B1(n19725), .B2(n24769), .ZN(
        n22308) );
  AOI221_X1 U21537 ( .B1(n24787), .B2(n8272), .C1(n24781), .C2(n8720), .A(
        n22289), .ZN(n22288) );
  OAI22_X1 U21538 ( .A1(n8962), .A2(n24775), .B1(n19724), .B2(n24769), .ZN(
        n22289) );
  AOI221_X1 U21539 ( .B1(n24787), .B2(n8271), .C1(n24781), .C2(n8719), .A(
        n22270), .ZN(n22269) );
  OAI22_X1 U21540 ( .A1(n8960), .A2(n24775), .B1(n19723), .B2(n24769), .ZN(
        n22270) );
  AOI221_X1 U21541 ( .B1(n24787), .B2(n8270), .C1(n24781), .C2(n8718), .A(
        n22251), .ZN(n22250) );
  OAI22_X1 U21542 ( .A1(n8958), .A2(n24775), .B1(n19722), .B2(n24769), .ZN(
        n22251) );
  AOI221_X1 U21543 ( .B1(n24787), .B2(n8269), .C1(n24781), .C2(n8717), .A(
        n22232), .ZN(n22231) );
  OAI22_X1 U21544 ( .A1(n8956), .A2(n24775), .B1(n19721), .B2(n24769), .ZN(
        n22232) );
  AOI221_X1 U21545 ( .B1(n24787), .B2(n8268), .C1(n24781), .C2(n8716), .A(
        n22213), .ZN(n22212) );
  OAI22_X1 U21546 ( .A1(n8954), .A2(n24775), .B1(n19720), .B2(n24769), .ZN(
        n22213) );
  AOI221_X1 U21547 ( .B1(n24787), .B2(n8267), .C1(n24781), .C2(n8715), .A(
        n22194), .ZN(n22193) );
  OAI22_X1 U21548 ( .A1(n8952), .A2(n24775), .B1(n19719), .B2(n24769), .ZN(
        n22194) );
  AOI221_X1 U21549 ( .B1(n24787), .B2(n8266), .C1(n24781), .C2(n8714), .A(
        n22175), .ZN(n22174) );
  OAI22_X1 U21550 ( .A1(n8950), .A2(n24775), .B1(n19718), .B2(n24769), .ZN(
        n22175) );
  AOI221_X1 U21551 ( .B1(n24787), .B2(n8265), .C1(n24781), .C2(n8713), .A(
        n22156), .ZN(n22155) );
  OAI22_X1 U21552 ( .A1(n8948), .A2(n24775), .B1(n19717), .B2(n24769), .ZN(
        n22156) );
  AOI221_X1 U21553 ( .B1(n24787), .B2(n8264), .C1(n24781), .C2(n8712), .A(
        n22137), .ZN(n22136) );
  OAI22_X1 U21554 ( .A1(n8946), .A2(n24775), .B1(n19716), .B2(n24769), .ZN(
        n22137) );
  AOI221_X1 U21555 ( .B1(n24787), .B2(n8263), .C1(n24781), .C2(n8711), .A(
        n22118), .ZN(n22117) );
  OAI22_X1 U21556 ( .A1(n8944), .A2(n24775), .B1(n19715), .B2(n24769), .ZN(
        n22118) );
  AOI221_X1 U21557 ( .B1(n24787), .B2(n8262), .C1(n24781), .C2(n8710), .A(
        n22099), .ZN(n22098) );
  OAI22_X1 U21558 ( .A1(n8942), .A2(n24775), .B1(n19714), .B2(n24769), .ZN(
        n22099) );
  AOI221_X1 U21559 ( .B1(n24788), .B2(n8261), .C1(n24782), .C2(n8709), .A(
        n22080), .ZN(n22079) );
  OAI22_X1 U21560 ( .A1(n8940), .A2(n24776), .B1(n19713), .B2(n24770), .ZN(
        n22080) );
  AOI221_X1 U21561 ( .B1(n24788), .B2(n8260), .C1(n24782), .C2(n8708), .A(
        n22061), .ZN(n22060) );
  OAI22_X1 U21562 ( .A1(n8938), .A2(n24776), .B1(n19712), .B2(n24770), .ZN(
        n22061) );
  AOI221_X1 U21563 ( .B1(n24788), .B2(n8259), .C1(n24782), .C2(n8707), .A(
        n22042), .ZN(n22041) );
  OAI22_X1 U21564 ( .A1(n8936), .A2(n24776), .B1(n19711), .B2(n24770), .ZN(
        n22042) );
  AOI221_X1 U21565 ( .B1(n24788), .B2(n8258), .C1(n24782), .C2(n8706), .A(
        n22023), .ZN(n22022) );
  OAI22_X1 U21566 ( .A1(n8934), .A2(n24776), .B1(n19710), .B2(n24770), .ZN(
        n22023) );
  AOI221_X1 U21567 ( .B1(n24788), .B2(n8257), .C1(n24782), .C2(n8705), .A(
        n22004), .ZN(n22003) );
  OAI22_X1 U21568 ( .A1(n8932), .A2(n24776), .B1(n19709), .B2(n24770), .ZN(
        n22004) );
  AOI221_X1 U21569 ( .B1(n24788), .B2(n8256), .C1(n24782), .C2(n8704), .A(
        n21985), .ZN(n21984) );
  OAI22_X1 U21570 ( .A1(n8930), .A2(n24776), .B1(n19708), .B2(n24770), .ZN(
        n21985) );
  AOI221_X1 U21571 ( .B1(n24788), .B2(n8255), .C1(n24782), .C2(n8703), .A(
        n21966), .ZN(n21965) );
  OAI22_X1 U21572 ( .A1(n8928), .A2(n24776), .B1(n20186), .B2(n24770), .ZN(
        n21966) );
  AOI221_X1 U21573 ( .B1(n24788), .B2(n8254), .C1(n24782), .C2(n8702), .A(
        n21947), .ZN(n21946) );
  OAI22_X1 U21574 ( .A1(n8926), .A2(n24776), .B1(n20185), .B2(n24770), .ZN(
        n21947) );
  AOI221_X1 U21575 ( .B1(n24788), .B2(n8253), .C1(n24782), .C2(n8701), .A(
        n21928), .ZN(n21927) );
  OAI22_X1 U21576 ( .A1(n8924), .A2(n24776), .B1(n20184), .B2(n24770), .ZN(
        n21928) );
  AOI221_X1 U21577 ( .B1(n24788), .B2(n8252), .C1(n24782), .C2(n8700), .A(
        n21909), .ZN(n21908) );
  OAI22_X1 U21578 ( .A1(n8922), .A2(n24776), .B1(n20183), .B2(n24770), .ZN(
        n21909) );
  AOI221_X1 U21579 ( .B1(n24788), .B2(n8251), .C1(n24782), .C2(n8699), .A(
        n21890), .ZN(n21889) );
  OAI22_X1 U21580 ( .A1(n8920), .A2(n24776), .B1(n20182), .B2(n24770), .ZN(
        n21890) );
  AOI221_X1 U21581 ( .B1(n24788), .B2(n8250), .C1(n24782), .C2(n8698), .A(
        n21871), .ZN(n21870) );
  OAI22_X1 U21582 ( .A1(n8918), .A2(n24776), .B1(n20181), .B2(n24770), .ZN(
        n21871) );
  AOI221_X1 U21583 ( .B1(n24789), .B2(n8249), .C1(n24783), .C2(n8697), .A(
        n21852), .ZN(n21851) );
  OAI22_X1 U21584 ( .A1(n8916), .A2(n24777), .B1(n20180), .B2(n24771), .ZN(
        n21852) );
  AOI221_X1 U21585 ( .B1(n24789), .B2(n8248), .C1(n24783), .C2(n8696), .A(
        n21833), .ZN(n21832) );
  OAI22_X1 U21586 ( .A1(n8914), .A2(n24777), .B1(n20179), .B2(n24771), .ZN(
        n21833) );
  AOI221_X1 U21587 ( .B1(n24789), .B2(n8247), .C1(n24783), .C2(n8695), .A(
        n21814), .ZN(n21813) );
  OAI22_X1 U21588 ( .A1(n8912), .A2(n24777), .B1(n20178), .B2(n24771), .ZN(
        n21814) );
  AOI221_X1 U21589 ( .B1(n24789), .B2(n8246), .C1(n24783), .C2(n8694), .A(
        n21795), .ZN(n21794) );
  OAI22_X1 U21590 ( .A1(n8910), .A2(n24777), .B1(n20177), .B2(n24771), .ZN(
        n21795) );
  AOI221_X1 U21591 ( .B1(n24789), .B2(n8245), .C1(n24783), .C2(n8693), .A(
        n21776), .ZN(n21775) );
  OAI22_X1 U21592 ( .A1(n8908), .A2(n24777), .B1(n20176), .B2(n24771), .ZN(
        n21776) );
  AOI221_X1 U21593 ( .B1(n24789), .B2(n8244), .C1(n24783), .C2(n8692), .A(
        n21757), .ZN(n21756) );
  OAI22_X1 U21594 ( .A1(n8906), .A2(n24777), .B1(n20175), .B2(n24771), .ZN(
        n21757) );
  AOI221_X1 U21595 ( .B1(n24789), .B2(n8243), .C1(n24783), .C2(n8691), .A(
        n21738), .ZN(n21737) );
  OAI22_X1 U21596 ( .A1(n8904), .A2(n24777), .B1(n20174), .B2(n24771), .ZN(
        n21738) );
  AOI221_X1 U21597 ( .B1(n24789), .B2(n8242), .C1(n24783), .C2(n8690), .A(
        n21719), .ZN(n21718) );
  OAI22_X1 U21598 ( .A1(n8902), .A2(n24777), .B1(n20173), .B2(n24771), .ZN(
        n21719) );
  AOI221_X1 U21599 ( .B1(n24789), .B2(n8241), .C1(n24783), .C2(n8689), .A(
        n21700), .ZN(n21699) );
  OAI22_X1 U21600 ( .A1(n8900), .A2(n24777), .B1(n20172), .B2(n24771), .ZN(
        n21700) );
  AOI221_X1 U21601 ( .B1(n24789), .B2(n8240), .C1(n24783), .C2(n8688), .A(
        n21681), .ZN(n21680) );
  OAI22_X1 U21602 ( .A1(n8898), .A2(n24777), .B1(n20171), .B2(n24771), .ZN(
        n21681) );
  AOI221_X1 U21603 ( .B1(n24789), .B2(n8239), .C1(n24783), .C2(n8687), .A(
        n21662), .ZN(n21661) );
  OAI22_X1 U21604 ( .A1(n8896), .A2(n24777), .B1(n20170), .B2(n24771), .ZN(
        n21662) );
  AOI221_X1 U21605 ( .B1(n24789), .B2(n8238), .C1(n24783), .C2(n8686), .A(
        n21643), .ZN(n21642) );
  OAI22_X1 U21606 ( .A1(n8894), .A2(n24777), .B1(n20169), .B2(n24771), .ZN(
        n21643) );
  AOI221_X1 U21607 ( .B1(n24790), .B2(n8237), .C1(n24784), .C2(n8685), .A(
        n21624), .ZN(n21623) );
  OAI22_X1 U21608 ( .A1(n8892), .A2(n24778), .B1(n20168), .B2(n24772), .ZN(
        n21624) );
  AOI221_X1 U21609 ( .B1(n24790), .B2(n8236), .C1(n24784), .C2(n8684), .A(
        n21605), .ZN(n21604) );
  OAI22_X1 U21610 ( .A1(n8890), .A2(n24778), .B1(n20167), .B2(n24772), .ZN(
        n21605) );
  AOI221_X1 U21611 ( .B1(n24790), .B2(n8235), .C1(n24784), .C2(n8683), .A(
        n21586), .ZN(n21585) );
  OAI22_X1 U21612 ( .A1(n8888), .A2(n24778), .B1(n20166), .B2(n24772), .ZN(
        n21586) );
  AOI221_X1 U21613 ( .B1(n24790), .B2(n8234), .C1(n24784), .C2(n8682), .A(
        n21567), .ZN(n21566) );
  OAI22_X1 U21614 ( .A1(n8886), .A2(n24778), .B1(n20165), .B2(n24772), .ZN(
        n21567) );
  AOI221_X1 U21615 ( .B1(n24790), .B2(n8233), .C1(n24784), .C2(n8681), .A(
        n21548), .ZN(n21547) );
  OAI22_X1 U21616 ( .A1(n8884), .A2(n24778), .B1(n20164), .B2(n24772), .ZN(
        n21548) );
  AOI221_X1 U21617 ( .B1(n24790), .B2(n8232), .C1(n24784), .C2(n8680), .A(
        n21529), .ZN(n21528) );
  OAI22_X1 U21618 ( .A1(n8882), .A2(n24778), .B1(n20163), .B2(n24772), .ZN(
        n21529) );
  AOI221_X1 U21619 ( .B1(n24790), .B2(n8231), .C1(n24784), .C2(n8679), .A(
        n21510), .ZN(n21509) );
  OAI22_X1 U21620 ( .A1(n8880), .A2(n24778), .B1(n20162), .B2(n24772), .ZN(
        n21510) );
  AOI221_X1 U21621 ( .B1(n24790), .B2(n8230), .C1(n24784), .C2(n8678), .A(
        n21491), .ZN(n21490) );
  OAI22_X1 U21622 ( .A1(n8878), .A2(n24778), .B1(n20161), .B2(n24772), .ZN(
        n21491) );
  AOI221_X1 U21623 ( .B1(n24790), .B2(n8229), .C1(n24784), .C2(n8677), .A(
        n21472), .ZN(n21471) );
  OAI22_X1 U21624 ( .A1(n8876), .A2(n24778), .B1(n20160), .B2(n24772), .ZN(
        n21472) );
  AOI221_X1 U21625 ( .B1(n24790), .B2(n8228), .C1(n24784), .C2(n8676), .A(
        n21453), .ZN(n21452) );
  OAI22_X1 U21626 ( .A1(n8874), .A2(n24778), .B1(n20159), .B2(n24772), .ZN(
        n21453) );
  AOI221_X1 U21627 ( .B1(n24790), .B2(n8227), .C1(n24784), .C2(n8675), .A(
        n21434), .ZN(n21433) );
  OAI22_X1 U21628 ( .A1(n8872), .A2(n24778), .B1(n20158), .B2(n24772), .ZN(
        n21434) );
  AOI221_X1 U21629 ( .B1(n24790), .B2(n8226), .C1(n24784), .C2(n8674), .A(
        n21415), .ZN(n21414) );
  OAI22_X1 U21630 ( .A1(n8870), .A2(n24778), .B1(n20157), .B2(n24772), .ZN(
        n21415) );
  AOI221_X1 U21631 ( .B1(n24791), .B2(n8225), .C1(n24785), .C2(n8673), .A(
        n21396), .ZN(n21395) );
  OAI22_X1 U21632 ( .A1(n8868), .A2(n24779), .B1(n20148), .B2(n24773), .ZN(
        n21396) );
  AOI221_X1 U21633 ( .B1(n24791), .B2(n8224), .C1(n24785), .C2(n8672), .A(
        n21377), .ZN(n21376) );
  OAI22_X1 U21634 ( .A1(n8866), .A2(n24779), .B1(n20147), .B2(n24773), .ZN(
        n21377) );
  AOI221_X1 U21635 ( .B1(n24791), .B2(n8223), .C1(n24785), .C2(n8671), .A(
        n21358), .ZN(n21357) );
  OAI22_X1 U21636 ( .A1(n8864), .A2(n24779), .B1(n20146), .B2(n24773), .ZN(
        n21358) );
  AOI221_X1 U21637 ( .B1(n24791), .B2(n8222), .C1(n24785), .C2(n8670), .A(
        n21309), .ZN(n21306) );
  OAI22_X1 U21638 ( .A1(n8862), .A2(n24779), .B1(n20145), .B2(n24773), .ZN(
        n21309) );
  AOI221_X1 U21639 ( .B1(n24690), .B2(n20073), .C1(n24684), .C2(n19523), .A(
        n22552), .ZN(n22551) );
  OAI22_X1 U21640 ( .A1(n896), .A2(n24678), .B1(n21074), .B2(n24672), .ZN(
        n22552) );
  AOI221_X1 U21641 ( .B1(n24690), .B2(n20072), .C1(n24684), .C2(n19522), .A(
        n22525), .ZN(n22524) );
  OAI22_X1 U21642 ( .A1(n895), .A2(n24678), .B1(n21073), .B2(n24672), .ZN(
        n22525) );
  AOI221_X1 U21643 ( .B1(n24690), .B2(n20071), .C1(n24684), .C2(n19521), .A(
        n22506), .ZN(n22505) );
  OAI22_X1 U21644 ( .A1(n894), .A2(n24678), .B1(n21072), .B2(n24672), .ZN(
        n22506) );
  AOI221_X1 U21645 ( .B1(n24690), .B2(n20070), .C1(n24684), .C2(n19520), .A(
        n22487), .ZN(n22486) );
  OAI22_X1 U21646 ( .A1(n893), .A2(n24678), .B1(n21071), .B2(n24672), .ZN(
        n22487) );
  AOI221_X1 U21647 ( .B1(n24690), .B2(n20069), .C1(n24684), .C2(n19519), .A(
        n22468), .ZN(n22467) );
  OAI22_X1 U21648 ( .A1(n892), .A2(n24678), .B1(n21070), .B2(n24672), .ZN(
        n22468) );
  AOI221_X1 U21649 ( .B1(n24690), .B2(n20068), .C1(n24684), .C2(n19518), .A(
        n22449), .ZN(n22448) );
  OAI22_X1 U21650 ( .A1(n891), .A2(n24678), .B1(n21069), .B2(n24672), .ZN(
        n22449) );
  AOI221_X1 U21651 ( .B1(n24690), .B2(n20067), .C1(n24684), .C2(n19517), .A(
        n22430), .ZN(n22429) );
  OAI22_X1 U21652 ( .A1(n890), .A2(n24678), .B1(n21068), .B2(n24672), .ZN(
        n22430) );
  AOI221_X1 U21653 ( .B1(n24690), .B2(n20066), .C1(n24684), .C2(n19516), .A(
        n22411), .ZN(n22410) );
  OAI22_X1 U21654 ( .A1(n889), .A2(n24678), .B1(n21067), .B2(n24672), .ZN(
        n22411) );
  AOI221_X1 U21655 ( .B1(n24690), .B2(n20065), .C1(n24684), .C2(n19515), .A(
        n22392), .ZN(n22391) );
  OAI22_X1 U21656 ( .A1(n888), .A2(n24678), .B1(n21066), .B2(n24672), .ZN(
        n22392) );
  AOI221_X1 U21657 ( .B1(n24690), .B2(n20064), .C1(n24684), .C2(n19514), .A(
        n22373), .ZN(n22372) );
  OAI22_X1 U21658 ( .A1(n887), .A2(n24678), .B1(n21065), .B2(n24672), .ZN(
        n22373) );
  AOI221_X1 U21659 ( .B1(n24690), .B2(n20063), .C1(n24684), .C2(n19513), .A(
        n22354), .ZN(n22353) );
  OAI22_X1 U21660 ( .A1(n886), .A2(n24678), .B1(n21064), .B2(n24672), .ZN(
        n22354) );
  AOI221_X1 U21661 ( .B1(n24690), .B2(n20062), .C1(n24684), .C2(n19512), .A(
        n22335), .ZN(n22334) );
  OAI22_X1 U21662 ( .A1(n885), .A2(n24678), .B1(n21063), .B2(n24672), .ZN(
        n22335) );
  AOI221_X1 U21663 ( .B1(n24691), .B2(n20061), .C1(n24685), .C2(n19511), .A(
        n22316), .ZN(n22315) );
  OAI22_X1 U21664 ( .A1(n884), .A2(n24679), .B1(n21062), .B2(n24673), .ZN(
        n22316) );
  AOI221_X1 U21665 ( .B1(n24691), .B2(n20060), .C1(n24685), .C2(n19510), .A(
        n22297), .ZN(n22296) );
  OAI22_X1 U21666 ( .A1(n883), .A2(n24679), .B1(n21061), .B2(n24673), .ZN(
        n22297) );
  AOI221_X1 U21667 ( .B1(n24691), .B2(n20059), .C1(n24685), .C2(n19509), .A(
        n22278), .ZN(n22277) );
  OAI22_X1 U21668 ( .A1(n882), .A2(n24679), .B1(n21060), .B2(n24673), .ZN(
        n22278) );
  AOI221_X1 U21669 ( .B1(n24691), .B2(n20058), .C1(n24685), .C2(n19508), .A(
        n22259), .ZN(n22258) );
  OAI22_X1 U21670 ( .A1(n881), .A2(n24679), .B1(n21059), .B2(n24673), .ZN(
        n22259) );
  AOI221_X1 U21671 ( .B1(n24691), .B2(n20057), .C1(n24685), .C2(n19507), .A(
        n22240), .ZN(n22239) );
  OAI22_X1 U21672 ( .A1(n880), .A2(n24679), .B1(n21058), .B2(n24673), .ZN(
        n22240) );
  AOI221_X1 U21673 ( .B1(n24691), .B2(n20056), .C1(n24685), .C2(n19506), .A(
        n22221), .ZN(n22220) );
  OAI22_X1 U21674 ( .A1(n879), .A2(n24679), .B1(n21057), .B2(n24673), .ZN(
        n22221) );
  AOI221_X1 U21675 ( .B1(n24691), .B2(n20055), .C1(n24685), .C2(n19505), .A(
        n22202), .ZN(n22201) );
  OAI22_X1 U21676 ( .A1(n878), .A2(n24679), .B1(n21056), .B2(n24673), .ZN(
        n22202) );
  AOI221_X1 U21677 ( .B1(n24691), .B2(n20054), .C1(n24685), .C2(n19504), .A(
        n22183), .ZN(n22182) );
  OAI22_X1 U21678 ( .A1(n877), .A2(n24679), .B1(n21055), .B2(n24673), .ZN(
        n22183) );
  AOI221_X1 U21679 ( .B1(n24691), .B2(n20053), .C1(n24685), .C2(n19503), .A(
        n22164), .ZN(n22163) );
  OAI22_X1 U21680 ( .A1(n876), .A2(n24679), .B1(n21054), .B2(n24673), .ZN(
        n22164) );
  AOI221_X1 U21681 ( .B1(n24691), .B2(n20052), .C1(n24685), .C2(n19502), .A(
        n22145), .ZN(n22144) );
  OAI22_X1 U21682 ( .A1(n875), .A2(n24679), .B1(n21053), .B2(n24673), .ZN(
        n22145) );
  AOI221_X1 U21683 ( .B1(n24691), .B2(n20051), .C1(n24685), .C2(n19501), .A(
        n22126), .ZN(n22125) );
  OAI22_X1 U21684 ( .A1(n874), .A2(n24679), .B1(n21052), .B2(n24673), .ZN(
        n22126) );
  AOI221_X1 U21685 ( .B1(n24691), .B2(n20050), .C1(n24685), .C2(n19500), .A(
        n22107), .ZN(n22106) );
  OAI22_X1 U21686 ( .A1(n873), .A2(n24679), .B1(n21051), .B2(n24673), .ZN(
        n22107) );
  AOI221_X1 U21687 ( .B1(n24692), .B2(n19929), .C1(n24686), .C2(n19499), .A(
        n22088), .ZN(n22087) );
  OAI22_X1 U21688 ( .A1(n872), .A2(n24680), .B1(n20942), .B2(n24674), .ZN(
        n22088) );
  AOI221_X1 U21689 ( .B1(n24692), .B2(n19928), .C1(n24686), .C2(n19498), .A(
        n22069), .ZN(n22068) );
  OAI22_X1 U21690 ( .A1(n871), .A2(n24680), .B1(n20941), .B2(n24674), .ZN(
        n22069) );
  AOI221_X1 U21691 ( .B1(n24692), .B2(n19927), .C1(n24686), .C2(n19497), .A(
        n22050), .ZN(n22049) );
  OAI22_X1 U21692 ( .A1(n870), .A2(n24680), .B1(n20940), .B2(n24674), .ZN(
        n22050) );
  AOI221_X1 U21693 ( .B1(n24692), .B2(n19926), .C1(n24686), .C2(n19496), .A(
        n22031), .ZN(n22030) );
  OAI22_X1 U21694 ( .A1(n869), .A2(n24680), .B1(n20939), .B2(n24674), .ZN(
        n22031) );
  AOI221_X1 U21695 ( .B1(n24692), .B2(n19925), .C1(n24686), .C2(n19495), .A(
        n22012), .ZN(n22011) );
  OAI22_X1 U21696 ( .A1(n868), .A2(n24680), .B1(n20938), .B2(n24674), .ZN(
        n22012) );
  AOI221_X1 U21697 ( .B1(n24692), .B2(n19924), .C1(n24686), .C2(n19494), .A(
        n21993), .ZN(n21992) );
  OAI22_X1 U21698 ( .A1(n867), .A2(n24680), .B1(n20937), .B2(n24674), .ZN(
        n21993) );
  AOI221_X1 U21699 ( .B1(n24692), .B2(n19923), .C1(n24686), .C2(n19493), .A(
        n21974), .ZN(n21973) );
  OAI22_X1 U21700 ( .A1(n866), .A2(n24680), .B1(n20936), .B2(n24674), .ZN(
        n21974) );
  AOI221_X1 U21701 ( .B1(n24692), .B2(n19922), .C1(n24686), .C2(n19492), .A(
        n21955), .ZN(n21954) );
  OAI22_X1 U21702 ( .A1(n865), .A2(n24680), .B1(n20935), .B2(n24674), .ZN(
        n21955) );
  AOI221_X1 U21703 ( .B1(n24692), .B2(n19921), .C1(n24686), .C2(n19491), .A(
        n21936), .ZN(n21935) );
  OAI22_X1 U21704 ( .A1(n864), .A2(n24680), .B1(n20934), .B2(n24674), .ZN(
        n21936) );
  AOI221_X1 U21705 ( .B1(n24692), .B2(n19920), .C1(n24686), .C2(n19490), .A(
        n21917), .ZN(n21916) );
  OAI22_X1 U21706 ( .A1(n863), .A2(n24680), .B1(n20933), .B2(n24674), .ZN(
        n21917) );
  AOI221_X1 U21707 ( .B1(n24692), .B2(n19919), .C1(n24686), .C2(n19489), .A(
        n21898), .ZN(n21897) );
  OAI22_X1 U21708 ( .A1(n862), .A2(n24680), .B1(n20932), .B2(n24674), .ZN(
        n21898) );
  AOI221_X1 U21709 ( .B1(n24692), .B2(n19918), .C1(n24686), .C2(n19488), .A(
        n21879), .ZN(n21878) );
  OAI22_X1 U21710 ( .A1(n861), .A2(n24680), .B1(n20931), .B2(n24674), .ZN(
        n21879) );
  AOI221_X1 U21711 ( .B1(n24693), .B2(n19917), .C1(n24687), .C2(n19487), .A(
        n21860), .ZN(n21859) );
  OAI22_X1 U21712 ( .A1(n860), .A2(n24681), .B1(n20930), .B2(n24675), .ZN(
        n21860) );
  AOI221_X1 U21713 ( .B1(n24693), .B2(n19916), .C1(n24687), .C2(n19486), .A(
        n21841), .ZN(n21840) );
  OAI22_X1 U21714 ( .A1(n859), .A2(n24681), .B1(n20929), .B2(n24675), .ZN(
        n21841) );
  AOI221_X1 U21715 ( .B1(n24693), .B2(n19915), .C1(n24687), .C2(n19485), .A(
        n21822), .ZN(n21821) );
  OAI22_X1 U21716 ( .A1(n858), .A2(n24681), .B1(n20928), .B2(n24675), .ZN(
        n21822) );
  AOI221_X1 U21717 ( .B1(n24693), .B2(n19914), .C1(n24687), .C2(n19484), .A(
        n21803), .ZN(n21802) );
  OAI22_X1 U21718 ( .A1(n857), .A2(n24681), .B1(n20927), .B2(n24675), .ZN(
        n21803) );
  AOI221_X1 U21719 ( .B1(n24693), .B2(n19913), .C1(n24687), .C2(n19483), .A(
        n21784), .ZN(n21783) );
  OAI22_X1 U21720 ( .A1(n856), .A2(n24681), .B1(n20926), .B2(n24675), .ZN(
        n21784) );
  AOI221_X1 U21721 ( .B1(n24693), .B2(n19912), .C1(n24687), .C2(n19482), .A(
        n21765), .ZN(n21764) );
  OAI22_X1 U21722 ( .A1(n855), .A2(n24681), .B1(n20925), .B2(n24675), .ZN(
        n21765) );
  AOI221_X1 U21723 ( .B1(n24693), .B2(n19911), .C1(n24687), .C2(n19481), .A(
        n21746), .ZN(n21745) );
  OAI22_X1 U21724 ( .A1(n854), .A2(n24681), .B1(n20924), .B2(n24675), .ZN(
        n21746) );
  AOI221_X1 U21725 ( .B1(n24693), .B2(n19910), .C1(n24687), .C2(n19480), .A(
        n21727), .ZN(n21726) );
  OAI22_X1 U21726 ( .A1(n853), .A2(n24681), .B1(n20923), .B2(n24675), .ZN(
        n21727) );
  AOI221_X1 U21727 ( .B1(n24693), .B2(n19909), .C1(n24687), .C2(n19479), .A(
        n21708), .ZN(n21707) );
  OAI22_X1 U21728 ( .A1(n852), .A2(n24681), .B1(n20922), .B2(n24675), .ZN(
        n21708) );
  AOI221_X1 U21729 ( .B1(n24693), .B2(n19908), .C1(n24687), .C2(n19478), .A(
        n21689), .ZN(n21688) );
  OAI22_X1 U21730 ( .A1(n851), .A2(n24681), .B1(n20921), .B2(n24675), .ZN(
        n21689) );
  AOI221_X1 U21731 ( .B1(n24693), .B2(n19907), .C1(n24687), .C2(n19477), .A(
        n21670), .ZN(n21669) );
  OAI22_X1 U21732 ( .A1(n850), .A2(n24681), .B1(n20920), .B2(n24675), .ZN(
        n21670) );
  AOI221_X1 U21733 ( .B1(n24693), .B2(n19906), .C1(n24687), .C2(n19476), .A(
        n21651), .ZN(n21650) );
  OAI22_X1 U21734 ( .A1(n849), .A2(n24681), .B1(n20919), .B2(n24675), .ZN(
        n21651) );
  AOI221_X1 U21735 ( .B1(n24694), .B2(n19905), .C1(n24688), .C2(n19475), .A(
        n21632), .ZN(n21631) );
  OAI22_X1 U21736 ( .A1(n848), .A2(n24682), .B1(n20918), .B2(n24676), .ZN(
        n21632) );
  AOI221_X1 U21737 ( .B1(n24694), .B2(n19904), .C1(n24688), .C2(n19474), .A(
        n21613), .ZN(n21612) );
  OAI22_X1 U21738 ( .A1(n847), .A2(n24682), .B1(n20917), .B2(n24676), .ZN(
        n21613) );
  AOI221_X1 U21739 ( .B1(n24694), .B2(n19903), .C1(n24688), .C2(n19473), .A(
        n21594), .ZN(n21593) );
  OAI22_X1 U21740 ( .A1(n846), .A2(n24682), .B1(n20916), .B2(n24676), .ZN(
        n21594) );
  AOI221_X1 U21741 ( .B1(n24694), .B2(n19902), .C1(n24688), .C2(n19472), .A(
        n21575), .ZN(n21574) );
  OAI22_X1 U21742 ( .A1(n845), .A2(n24682), .B1(n20915), .B2(n24676), .ZN(
        n21575) );
  AOI221_X1 U21743 ( .B1(n24694), .B2(n19901), .C1(n24688), .C2(n19471), .A(
        n21556), .ZN(n21555) );
  OAI22_X1 U21744 ( .A1(n844), .A2(n24682), .B1(n20914), .B2(n24676), .ZN(
        n21556) );
  AOI221_X1 U21745 ( .B1(n24694), .B2(n19900), .C1(n24688), .C2(n19470), .A(
        n21537), .ZN(n21536) );
  OAI22_X1 U21746 ( .A1(n843), .A2(n24682), .B1(n20913), .B2(n24676), .ZN(
        n21537) );
  AOI221_X1 U21747 ( .B1(n24694), .B2(n19899), .C1(n24688), .C2(n19469), .A(
        n21518), .ZN(n21517) );
  OAI22_X1 U21748 ( .A1(n842), .A2(n24682), .B1(n20912), .B2(n24676), .ZN(
        n21518) );
  AOI221_X1 U21749 ( .B1(n24694), .B2(n19898), .C1(n24688), .C2(n19468), .A(
        n21499), .ZN(n21498) );
  OAI22_X1 U21750 ( .A1(n841), .A2(n24682), .B1(n20911), .B2(n24676), .ZN(
        n21499) );
  AOI221_X1 U21751 ( .B1(n24694), .B2(n19897), .C1(n24688), .C2(n19467), .A(
        n21480), .ZN(n21479) );
  OAI22_X1 U21752 ( .A1(n840), .A2(n24682), .B1(n20910), .B2(n24676), .ZN(
        n21480) );
  AOI221_X1 U21753 ( .B1(n24694), .B2(n19896), .C1(n24688), .C2(n19466), .A(
        n21461), .ZN(n21460) );
  OAI22_X1 U21754 ( .A1(n839), .A2(n24682), .B1(n20909), .B2(n24676), .ZN(
        n21461) );
  AOI221_X1 U21755 ( .B1(n24694), .B2(n19895), .C1(n24688), .C2(n19465), .A(
        n21442), .ZN(n21441) );
  OAI22_X1 U21756 ( .A1(n838), .A2(n24682), .B1(n20908), .B2(n24676), .ZN(
        n21442) );
  AOI221_X1 U21757 ( .B1(n24694), .B2(n19894), .C1(n24688), .C2(n19464), .A(
        n21423), .ZN(n21422) );
  OAI22_X1 U21758 ( .A1(n837), .A2(n24682), .B1(n20907), .B2(n24676), .ZN(
        n21423) );
  AOI221_X1 U21759 ( .B1(n24695), .B2(n19813), .C1(n24689), .C2(n19463), .A(
        n21404), .ZN(n21403) );
  OAI22_X1 U21760 ( .A1(n836), .A2(n24683), .B1(n20534), .B2(n24677), .ZN(
        n21404) );
  AOI221_X1 U21761 ( .B1(n24695), .B2(n19812), .C1(n24689), .C2(n19462), .A(
        n21385), .ZN(n21384) );
  OAI22_X1 U21762 ( .A1(n835), .A2(n24683), .B1(n20533), .B2(n24677), .ZN(
        n21385) );
  AOI221_X1 U21763 ( .B1(n24695), .B2(n19811), .C1(n24689), .C2(n19461), .A(
        n21366), .ZN(n21365) );
  OAI22_X1 U21764 ( .A1(n834), .A2(n24683), .B1(n20532), .B2(n24677), .ZN(
        n21366) );
  AOI221_X1 U21765 ( .B1(n24695), .B2(n19810), .C1(n24689), .C2(n19460), .A(
        n21333), .ZN(n21330) );
  OAI22_X1 U21766 ( .A1(n833), .A2(n24683), .B1(n20531), .B2(n24677), .ZN(
        n21333) );
  AOI221_X1 U21767 ( .B1(n24762), .B2(n8029), .C1(n24756), .C2(n8413), .A(
        n22541), .ZN(n22534) );
  OAI22_X1 U21768 ( .A1(n7427), .A2(n24750), .B1(n19707), .B2(n24744), .ZN(
        n22541) );
  AOI221_X1 U21769 ( .B1(n24762), .B2(n8028), .C1(n24756), .C2(n8412), .A(
        n22518), .ZN(n22515) );
  OAI22_X1 U21770 ( .A1(n7425), .A2(n24750), .B1(n19706), .B2(n24744), .ZN(
        n22518) );
  AOI221_X1 U21771 ( .B1(n24762), .B2(n8027), .C1(n24756), .C2(n8411), .A(
        n22499), .ZN(n22496) );
  OAI22_X1 U21772 ( .A1(n7423), .A2(n24750), .B1(n19705), .B2(n24744), .ZN(
        n22499) );
  AOI221_X1 U21773 ( .B1(n24762), .B2(n8026), .C1(n24756), .C2(n8410), .A(
        n22480), .ZN(n22477) );
  OAI22_X1 U21774 ( .A1(n7421), .A2(n24750), .B1(n19704), .B2(n24744), .ZN(
        n22480) );
  AOI221_X1 U21775 ( .B1(n24762), .B2(n8025), .C1(n24756), .C2(n8409), .A(
        n22461), .ZN(n22458) );
  OAI22_X1 U21776 ( .A1(n7419), .A2(n24750), .B1(n19703), .B2(n24744), .ZN(
        n22461) );
  AOI221_X1 U21777 ( .B1(n24762), .B2(n8024), .C1(n24756), .C2(n8408), .A(
        n22442), .ZN(n22439) );
  OAI22_X1 U21778 ( .A1(n7417), .A2(n24750), .B1(n19702), .B2(n24744), .ZN(
        n22442) );
  AOI221_X1 U21779 ( .B1(n24762), .B2(n8023), .C1(n24756), .C2(n8407), .A(
        n22423), .ZN(n22420) );
  OAI22_X1 U21780 ( .A1(n7415), .A2(n24750), .B1(n19701), .B2(n24744), .ZN(
        n22423) );
  AOI221_X1 U21781 ( .B1(n24762), .B2(n8022), .C1(n24756), .C2(n8406), .A(
        n22404), .ZN(n22401) );
  OAI22_X1 U21782 ( .A1(n7413), .A2(n24750), .B1(n19700), .B2(n24744), .ZN(
        n22404) );
  AOI221_X1 U21783 ( .B1(n24762), .B2(n8021), .C1(n24756), .C2(n8405), .A(
        n22385), .ZN(n22382) );
  OAI22_X1 U21784 ( .A1(n7411), .A2(n24750), .B1(n19699), .B2(n24744), .ZN(
        n22385) );
  AOI221_X1 U21785 ( .B1(n24762), .B2(n8020), .C1(n24756), .C2(n8404), .A(
        n22366), .ZN(n22363) );
  OAI22_X1 U21786 ( .A1(n7409), .A2(n24750), .B1(n19698), .B2(n24744), .ZN(
        n22366) );
  AOI221_X1 U21787 ( .B1(n24762), .B2(n8019), .C1(n24756), .C2(n8403), .A(
        n22347), .ZN(n22344) );
  OAI22_X1 U21788 ( .A1(n7407), .A2(n24750), .B1(n19697), .B2(n24744), .ZN(
        n22347) );
  AOI221_X1 U21789 ( .B1(n24762), .B2(n8018), .C1(n24756), .C2(n8402), .A(
        n22328), .ZN(n22325) );
  OAI22_X1 U21790 ( .A1(n7405), .A2(n24750), .B1(n19696), .B2(n24744), .ZN(
        n22328) );
  AOI221_X1 U21791 ( .B1(n24763), .B2(n8017), .C1(n24757), .C2(n8401), .A(
        n22309), .ZN(n22306) );
  OAI22_X1 U21792 ( .A1(n7403), .A2(n24751), .B1(n19695), .B2(n24745), .ZN(
        n22309) );
  AOI221_X1 U21793 ( .B1(n24763), .B2(n8016), .C1(n24757), .C2(n8400), .A(
        n22290), .ZN(n22287) );
  OAI22_X1 U21794 ( .A1(n7401), .A2(n24751), .B1(n19694), .B2(n24745), .ZN(
        n22290) );
  AOI221_X1 U21795 ( .B1(n24763), .B2(n8015), .C1(n24757), .C2(n8399), .A(
        n22271), .ZN(n22268) );
  OAI22_X1 U21796 ( .A1(n7399), .A2(n24751), .B1(n19693), .B2(n24745), .ZN(
        n22271) );
  AOI221_X1 U21797 ( .B1(n24763), .B2(n8014), .C1(n24757), .C2(n8398), .A(
        n22252), .ZN(n22249) );
  OAI22_X1 U21798 ( .A1(n7397), .A2(n24751), .B1(n19692), .B2(n24745), .ZN(
        n22252) );
  AOI221_X1 U21799 ( .B1(n24763), .B2(n8013), .C1(n24757), .C2(n8397), .A(
        n22233), .ZN(n22230) );
  OAI22_X1 U21800 ( .A1(n7395), .A2(n24751), .B1(n19691), .B2(n24745), .ZN(
        n22233) );
  AOI221_X1 U21801 ( .B1(n24763), .B2(n8012), .C1(n24757), .C2(n8396), .A(
        n22214), .ZN(n22211) );
  OAI22_X1 U21802 ( .A1(n7393), .A2(n24751), .B1(n19690), .B2(n24745), .ZN(
        n22214) );
  AOI221_X1 U21803 ( .B1(n24763), .B2(n8011), .C1(n24757), .C2(n8395), .A(
        n22195), .ZN(n22192) );
  OAI22_X1 U21804 ( .A1(n7391), .A2(n24751), .B1(n19689), .B2(n24745), .ZN(
        n22195) );
  AOI221_X1 U21805 ( .B1(n24763), .B2(n8010), .C1(n24757), .C2(n8394), .A(
        n22176), .ZN(n22173) );
  OAI22_X1 U21806 ( .A1(n7389), .A2(n24751), .B1(n19688), .B2(n24745), .ZN(
        n22176) );
  AOI221_X1 U21807 ( .B1(n24763), .B2(n8009), .C1(n24757), .C2(n8393), .A(
        n22157), .ZN(n22154) );
  OAI22_X1 U21808 ( .A1(n7387), .A2(n24751), .B1(n19687), .B2(n24745), .ZN(
        n22157) );
  AOI221_X1 U21809 ( .B1(n24763), .B2(n8008), .C1(n24757), .C2(n8392), .A(
        n22138), .ZN(n22135) );
  OAI22_X1 U21810 ( .A1(n7385), .A2(n24751), .B1(n19686), .B2(n24745), .ZN(
        n22138) );
  AOI221_X1 U21811 ( .B1(n24763), .B2(n8007), .C1(n24757), .C2(n8391), .A(
        n22119), .ZN(n22116) );
  OAI22_X1 U21812 ( .A1(n7383), .A2(n24751), .B1(n19685), .B2(n24745), .ZN(
        n22119) );
  AOI221_X1 U21813 ( .B1(n24763), .B2(n8006), .C1(n24757), .C2(n8390), .A(
        n22100), .ZN(n22097) );
  OAI22_X1 U21814 ( .A1(n7381), .A2(n24751), .B1(n19684), .B2(n24745), .ZN(
        n22100) );
  AOI221_X1 U21815 ( .B1(n24764), .B2(n8005), .C1(n24758), .C2(n8389), .A(
        n22081), .ZN(n22078) );
  OAI22_X1 U21816 ( .A1(n7379), .A2(n24752), .B1(n19683), .B2(n24746), .ZN(
        n22081) );
  AOI221_X1 U21817 ( .B1(n24764), .B2(n8004), .C1(n24758), .C2(n8388), .A(
        n22062), .ZN(n22059) );
  OAI22_X1 U21818 ( .A1(n7377), .A2(n24752), .B1(n19682), .B2(n24746), .ZN(
        n22062) );
  AOI221_X1 U21819 ( .B1(n24764), .B2(n8003), .C1(n24758), .C2(n8387), .A(
        n22043), .ZN(n22040) );
  OAI22_X1 U21820 ( .A1(n7375), .A2(n24752), .B1(n19681), .B2(n24746), .ZN(
        n22043) );
  AOI221_X1 U21821 ( .B1(n24764), .B2(n8002), .C1(n24758), .C2(n8386), .A(
        n22024), .ZN(n22021) );
  OAI22_X1 U21822 ( .A1(n7373), .A2(n24752), .B1(n19680), .B2(n24746), .ZN(
        n22024) );
  AOI221_X1 U21823 ( .B1(n24764), .B2(n8001), .C1(n24758), .C2(n8385), .A(
        n22005), .ZN(n22002) );
  OAI22_X1 U21824 ( .A1(n7371), .A2(n24752), .B1(n19679), .B2(n24746), .ZN(
        n22005) );
  AOI221_X1 U21825 ( .B1(n24764), .B2(n8000), .C1(n24758), .C2(n8384), .A(
        n21986), .ZN(n21983) );
  OAI22_X1 U21826 ( .A1(n7369), .A2(n24752), .B1(n19678), .B2(n24746), .ZN(
        n21986) );
  AOI221_X1 U21827 ( .B1(n24764), .B2(n7999), .C1(n24758), .C2(n8383), .A(
        n21967), .ZN(n21964) );
  OAI22_X1 U21828 ( .A1(n7367), .A2(n24752), .B1(n19677), .B2(n24746), .ZN(
        n21967) );
  AOI221_X1 U21829 ( .B1(n24764), .B2(n7998), .C1(n24758), .C2(n8382), .A(
        n21948), .ZN(n21945) );
  OAI22_X1 U21830 ( .A1(n7365), .A2(n24752), .B1(n19676), .B2(n24746), .ZN(
        n21948) );
  AOI221_X1 U21831 ( .B1(n24764), .B2(n7997), .C1(n24758), .C2(n8381), .A(
        n21929), .ZN(n21926) );
  OAI22_X1 U21832 ( .A1(n7363), .A2(n24752), .B1(n19675), .B2(n24746), .ZN(
        n21929) );
  AOI221_X1 U21833 ( .B1(n24764), .B2(n7996), .C1(n24758), .C2(n8380), .A(
        n21910), .ZN(n21907) );
  OAI22_X1 U21834 ( .A1(n7361), .A2(n24752), .B1(n19674), .B2(n24746), .ZN(
        n21910) );
  AOI221_X1 U21835 ( .B1(n24764), .B2(n7995), .C1(n24758), .C2(n8379), .A(
        n21891), .ZN(n21888) );
  OAI22_X1 U21836 ( .A1(n7359), .A2(n24752), .B1(n19673), .B2(n24746), .ZN(
        n21891) );
  AOI221_X1 U21837 ( .B1(n24764), .B2(n7994), .C1(n24758), .C2(n8378), .A(
        n21872), .ZN(n21869) );
  OAI22_X1 U21838 ( .A1(n7357), .A2(n24752), .B1(n19672), .B2(n24746), .ZN(
        n21872) );
  AOI221_X1 U21839 ( .B1(n24765), .B2(n7993), .C1(n24759), .C2(n8377), .A(
        n21853), .ZN(n21850) );
  OAI22_X1 U21840 ( .A1(n7355), .A2(n24753), .B1(n19671), .B2(n24747), .ZN(
        n21853) );
  AOI221_X1 U21841 ( .B1(n24765), .B2(n7992), .C1(n24759), .C2(n8376), .A(
        n21834), .ZN(n21831) );
  OAI22_X1 U21842 ( .A1(n7353), .A2(n24753), .B1(n19670), .B2(n24747), .ZN(
        n21834) );
  AOI221_X1 U21843 ( .B1(n24765), .B2(n7991), .C1(n24759), .C2(n8375), .A(
        n21815), .ZN(n21812) );
  OAI22_X1 U21844 ( .A1(n7351), .A2(n24753), .B1(n19669), .B2(n24747), .ZN(
        n21815) );
  AOI221_X1 U21845 ( .B1(n24765), .B2(n7990), .C1(n24759), .C2(n8374), .A(
        n21796), .ZN(n21793) );
  OAI22_X1 U21846 ( .A1(n7349), .A2(n24753), .B1(n19668), .B2(n24747), .ZN(
        n21796) );
  AOI221_X1 U21847 ( .B1(n24765), .B2(n7989), .C1(n24759), .C2(n8373), .A(
        n21777), .ZN(n21774) );
  OAI22_X1 U21848 ( .A1(n7347), .A2(n24753), .B1(n19667), .B2(n24747), .ZN(
        n21777) );
  AOI221_X1 U21849 ( .B1(n24765), .B2(n7988), .C1(n24759), .C2(n8372), .A(
        n21758), .ZN(n21755) );
  OAI22_X1 U21850 ( .A1(n7345), .A2(n24753), .B1(n19666), .B2(n24747), .ZN(
        n21758) );
  AOI221_X1 U21851 ( .B1(n24765), .B2(n7987), .C1(n24759), .C2(n8371), .A(
        n21739), .ZN(n21736) );
  OAI22_X1 U21852 ( .A1(n7343), .A2(n24753), .B1(n19665), .B2(n24747), .ZN(
        n21739) );
  AOI221_X1 U21853 ( .B1(n24765), .B2(n7986), .C1(n24759), .C2(n8370), .A(
        n21720), .ZN(n21717) );
  OAI22_X1 U21854 ( .A1(n7341), .A2(n24753), .B1(n19664), .B2(n24747), .ZN(
        n21720) );
  AOI221_X1 U21855 ( .B1(n24765), .B2(n7985), .C1(n24759), .C2(n8369), .A(
        n21701), .ZN(n21698) );
  OAI22_X1 U21856 ( .A1(n7339), .A2(n24753), .B1(n19663), .B2(n24747), .ZN(
        n21701) );
  AOI221_X1 U21857 ( .B1(n24765), .B2(n7984), .C1(n24759), .C2(n8368), .A(
        n21682), .ZN(n21679) );
  OAI22_X1 U21858 ( .A1(n7337), .A2(n24753), .B1(n19662), .B2(n24747), .ZN(
        n21682) );
  AOI221_X1 U21859 ( .B1(n24765), .B2(n7983), .C1(n24759), .C2(n8367), .A(
        n21663), .ZN(n21660) );
  OAI22_X1 U21860 ( .A1(n7335), .A2(n24753), .B1(n19661), .B2(n24747), .ZN(
        n21663) );
  AOI221_X1 U21861 ( .B1(n24765), .B2(n7982), .C1(n24759), .C2(n8366), .A(
        n21644), .ZN(n21641) );
  OAI22_X1 U21862 ( .A1(n7333), .A2(n24753), .B1(n19660), .B2(n24747), .ZN(
        n21644) );
  AOI221_X1 U21863 ( .B1(n24766), .B2(n7981), .C1(n24760), .C2(n8365), .A(
        n21625), .ZN(n21622) );
  OAI22_X1 U21864 ( .A1(n7331), .A2(n24754), .B1(n19659), .B2(n24748), .ZN(
        n21625) );
  AOI221_X1 U21865 ( .B1(n24766), .B2(n7980), .C1(n24760), .C2(n8364), .A(
        n21606), .ZN(n21603) );
  OAI22_X1 U21866 ( .A1(n7329), .A2(n24754), .B1(n19658), .B2(n24748), .ZN(
        n21606) );
  AOI221_X1 U21867 ( .B1(n24766), .B2(n7979), .C1(n24760), .C2(n8363), .A(
        n21587), .ZN(n21584) );
  OAI22_X1 U21868 ( .A1(n7327), .A2(n24754), .B1(n19657), .B2(n24748), .ZN(
        n21587) );
  AOI221_X1 U21869 ( .B1(n24766), .B2(n7978), .C1(n24760), .C2(n8362), .A(
        n21568), .ZN(n21565) );
  OAI22_X1 U21870 ( .A1(n7325), .A2(n24754), .B1(n19656), .B2(n24748), .ZN(
        n21568) );
  AOI221_X1 U21871 ( .B1(n24766), .B2(n7977), .C1(n24760), .C2(n8361), .A(
        n21549), .ZN(n21546) );
  OAI22_X1 U21872 ( .A1(n7323), .A2(n24754), .B1(n19655), .B2(n24748), .ZN(
        n21549) );
  AOI221_X1 U21873 ( .B1(n24766), .B2(n7976), .C1(n24760), .C2(n8360), .A(
        n21530), .ZN(n21527) );
  OAI22_X1 U21874 ( .A1(n7321), .A2(n24754), .B1(n19654), .B2(n24748), .ZN(
        n21530) );
  AOI221_X1 U21875 ( .B1(n24766), .B2(n7975), .C1(n24760), .C2(n8359), .A(
        n21511), .ZN(n21508) );
  OAI22_X1 U21876 ( .A1(n7319), .A2(n24754), .B1(n19653), .B2(n24748), .ZN(
        n21511) );
  AOI221_X1 U21877 ( .B1(n24766), .B2(n7974), .C1(n24760), .C2(n8358), .A(
        n21492), .ZN(n21489) );
  OAI22_X1 U21878 ( .A1(n7317), .A2(n24754), .B1(n19652), .B2(n24748), .ZN(
        n21492) );
  AOI221_X1 U21879 ( .B1(n24766), .B2(n7973), .C1(n24760), .C2(n8357), .A(
        n21473), .ZN(n21470) );
  OAI22_X1 U21880 ( .A1(n7315), .A2(n24754), .B1(n19651), .B2(n24748), .ZN(
        n21473) );
  AOI221_X1 U21881 ( .B1(n24766), .B2(n7972), .C1(n24760), .C2(n8356), .A(
        n21454), .ZN(n21451) );
  OAI22_X1 U21882 ( .A1(n7313), .A2(n24754), .B1(n19650), .B2(n24748), .ZN(
        n21454) );
  AOI221_X1 U21883 ( .B1(n24766), .B2(n7971), .C1(n24760), .C2(n8355), .A(
        n21435), .ZN(n21432) );
  OAI22_X1 U21884 ( .A1(n7311), .A2(n24754), .B1(n19649), .B2(n24748), .ZN(
        n21435) );
  AOI221_X1 U21885 ( .B1(n24766), .B2(n7970), .C1(n24760), .C2(n8354), .A(
        n21416), .ZN(n21413) );
  OAI22_X1 U21886 ( .A1(n7309), .A2(n24754), .B1(n19648), .B2(n24748), .ZN(
        n21416) );
  AOI221_X1 U21887 ( .B1(n24767), .B2(n7969), .C1(n24761), .C2(n8353), .A(
        n21397), .ZN(n21394) );
  OAI22_X1 U21888 ( .A1(n7307), .A2(n24755), .B1(n20152), .B2(n24749), .ZN(
        n21397) );
  AOI221_X1 U21889 ( .B1(n24767), .B2(n7968), .C1(n24761), .C2(n8352), .A(
        n21378), .ZN(n21375) );
  OAI22_X1 U21890 ( .A1(n7305), .A2(n24755), .B1(n20151), .B2(n24749), .ZN(
        n21378) );
  AOI221_X1 U21891 ( .B1(n24767), .B2(n7967), .C1(n24761), .C2(n8351), .A(
        n21359), .ZN(n21356) );
  OAI22_X1 U21892 ( .A1(n7303), .A2(n24755), .B1(n20150), .B2(n24749), .ZN(
        n21359) );
  AOI221_X1 U21893 ( .B1(n24767), .B2(n7966), .C1(n24761), .C2(n8350), .A(
        n21314), .ZN(n21305) );
  OAI22_X1 U21894 ( .A1(n7301), .A2(n24755), .B1(n20149), .B2(n24749), .ZN(
        n21314) );
  AOI221_X1 U21895 ( .B1(n24671), .B2(n19399), .C1(n24665), .C2(n19817), .A(
        n21405), .ZN(n21402) );
  OAI22_X1 U21896 ( .A1(n20257), .A2(n24659), .B1(n20538), .B2(n24653), .ZN(
        n21405) );
  AOI221_X1 U21897 ( .B1(n24671), .B2(n19398), .C1(n24665), .C2(n19816), .A(
        n21386), .ZN(n21383) );
  OAI22_X1 U21898 ( .A1(n20256), .A2(n24659), .B1(n20537), .B2(n24653), .ZN(
        n21386) );
  AOI221_X1 U21899 ( .B1(n24671), .B2(n19397), .C1(n24665), .C2(n19815), .A(
        n21367), .ZN(n21364) );
  OAI22_X1 U21900 ( .A1(n20255), .A2(n24659), .B1(n20536), .B2(n24653), .ZN(
        n21367) );
  AOI221_X1 U21901 ( .B1(n24671), .B2(n19396), .C1(n24665), .C2(n19814), .A(
        n21338), .ZN(n21329) );
  OAI22_X1 U21902 ( .A1(n20254), .A2(n24659), .B1(n20535), .B2(n24653), .ZN(
        n21338) );
  AOI221_X1 U21903 ( .B1(n24738), .B2(n19647), .C1(n24732), .C2(n19587), .A(
        n22544), .ZN(n22533) );
  OAI22_X1 U21904 ( .A1(n21146), .A2(n24726), .B1(n20798), .B2(n24720), .ZN(
        n22544) );
  AOI221_X1 U21905 ( .B1(n24738), .B2(n19646), .C1(n24732), .C2(n19586), .A(
        n22519), .ZN(n22514) );
  OAI22_X1 U21906 ( .A1(n21145), .A2(n24726), .B1(n20797), .B2(n24720), .ZN(
        n22519) );
  AOI221_X1 U21907 ( .B1(n24738), .B2(n19645), .C1(n24732), .C2(n19585), .A(
        n22500), .ZN(n22495) );
  OAI22_X1 U21908 ( .A1(n21144), .A2(n24726), .B1(n20796), .B2(n24720), .ZN(
        n22500) );
  AOI221_X1 U21909 ( .B1(n24738), .B2(n19644), .C1(n24732), .C2(n19584), .A(
        n22481), .ZN(n22476) );
  OAI22_X1 U21910 ( .A1(n21143), .A2(n24726), .B1(n20795), .B2(n24720), .ZN(
        n22481) );
  AOI221_X1 U21911 ( .B1(n24738), .B2(n19643), .C1(n24732), .C2(n19583), .A(
        n22462), .ZN(n22457) );
  OAI22_X1 U21912 ( .A1(n21142), .A2(n24726), .B1(n20794), .B2(n24720), .ZN(
        n22462) );
  AOI221_X1 U21913 ( .B1(n24738), .B2(n19642), .C1(n24732), .C2(n19582), .A(
        n22443), .ZN(n22438) );
  OAI22_X1 U21914 ( .A1(n21141), .A2(n24726), .B1(n20793), .B2(n24720), .ZN(
        n22443) );
  AOI221_X1 U21915 ( .B1(n24738), .B2(n19641), .C1(n24732), .C2(n19581), .A(
        n22424), .ZN(n22419) );
  OAI22_X1 U21916 ( .A1(n21140), .A2(n24726), .B1(n20792), .B2(n24720), .ZN(
        n22424) );
  AOI221_X1 U21917 ( .B1(n24738), .B2(n19640), .C1(n24732), .C2(n19580), .A(
        n22405), .ZN(n22400) );
  OAI22_X1 U21918 ( .A1(n21139), .A2(n24726), .B1(n20791), .B2(n24720), .ZN(
        n22405) );
  AOI221_X1 U21919 ( .B1(n24738), .B2(n19639), .C1(n24732), .C2(n19579), .A(
        n22386), .ZN(n22381) );
  OAI22_X1 U21920 ( .A1(n21138), .A2(n24726), .B1(n20790), .B2(n24720), .ZN(
        n22386) );
  AOI221_X1 U21921 ( .B1(n24738), .B2(n19638), .C1(n24732), .C2(n19578), .A(
        n22367), .ZN(n22362) );
  OAI22_X1 U21922 ( .A1(n21137), .A2(n24726), .B1(n20789), .B2(n24720), .ZN(
        n22367) );
  AOI221_X1 U21923 ( .B1(n24738), .B2(n19637), .C1(n24732), .C2(n19577), .A(
        n22348), .ZN(n22343) );
  OAI22_X1 U21924 ( .A1(n21136), .A2(n24726), .B1(n20788), .B2(n24720), .ZN(
        n22348) );
  AOI221_X1 U21925 ( .B1(n24738), .B2(n19636), .C1(n24732), .C2(n19576), .A(
        n22329), .ZN(n22324) );
  OAI22_X1 U21926 ( .A1(n21135), .A2(n24726), .B1(n20787), .B2(n24720), .ZN(
        n22329) );
  AOI221_X1 U21927 ( .B1(n24739), .B2(n19635), .C1(n24733), .C2(n19575), .A(
        n22310), .ZN(n22305) );
  OAI22_X1 U21928 ( .A1(n21134), .A2(n24727), .B1(n20786), .B2(n24721), .ZN(
        n22310) );
  AOI221_X1 U21929 ( .B1(n24739), .B2(n19634), .C1(n24733), .C2(n19574), .A(
        n22291), .ZN(n22286) );
  OAI22_X1 U21930 ( .A1(n21133), .A2(n24727), .B1(n20785), .B2(n24721), .ZN(
        n22291) );
  AOI221_X1 U21931 ( .B1(n24739), .B2(n19633), .C1(n24733), .C2(n19573), .A(
        n22272), .ZN(n22267) );
  OAI22_X1 U21932 ( .A1(n21132), .A2(n24727), .B1(n20784), .B2(n24721), .ZN(
        n22272) );
  AOI221_X1 U21933 ( .B1(n24739), .B2(n19632), .C1(n24733), .C2(n19572), .A(
        n22253), .ZN(n22248) );
  OAI22_X1 U21934 ( .A1(n21131), .A2(n24727), .B1(n20783), .B2(n24721), .ZN(
        n22253) );
  AOI221_X1 U21935 ( .B1(n24739), .B2(n19631), .C1(n24733), .C2(n19571), .A(
        n22234), .ZN(n22229) );
  OAI22_X1 U21936 ( .A1(n21130), .A2(n24727), .B1(n20782), .B2(n24721), .ZN(
        n22234) );
  AOI221_X1 U21937 ( .B1(n24739), .B2(n19630), .C1(n24733), .C2(n19570), .A(
        n22215), .ZN(n22210) );
  OAI22_X1 U21938 ( .A1(n21129), .A2(n24727), .B1(n20781), .B2(n24721), .ZN(
        n22215) );
  AOI221_X1 U21939 ( .B1(n24739), .B2(n19629), .C1(n24733), .C2(n19569), .A(
        n22196), .ZN(n22191) );
  OAI22_X1 U21940 ( .A1(n21128), .A2(n24727), .B1(n20780), .B2(n24721), .ZN(
        n22196) );
  AOI221_X1 U21941 ( .B1(n24739), .B2(n19628), .C1(n24733), .C2(n19568), .A(
        n22177), .ZN(n22172) );
  OAI22_X1 U21942 ( .A1(n21127), .A2(n24727), .B1(n20779), .B2(n24721), .ZN(
        n22177) );
  AOI221_X1 U21943 ( .B1(n24739), .B2(n19627), .C1(n24733), .C2(n19567), .A(
        n22158), .ZN(n22153) );
  OAI22_X1 U21944 ( .A1(n21126), .A2(n24727), .B1(n20778), .B2(n24721), .ZN(
        n22158) );
  AOI221_X1 U21945 ( .B1(n24739), .B2(n19626), .C1(n24733), .C2(n19566), .A(
        n22139), .ZN(n22134) );
  OAI22_X1 U21946 ( .A1(n21125), .A2(n24727), .B1(n20777), .B2(n24721), .ZN(
        n22139) );
  AOI221_X1 U21947 ( .B1(n24739), .B2(n19625), .C1(n24733), .C2(n19565), .A(
        n22120), .ZN(n22115) );
  OAI22_X1 U21948 ( .A1(n21124), .A2(n24727), .B1(n20776), .B2(n24721), .ZN(
        n22120) );
  AOI221_X1 U21949 ( .B1(n24739), .B2(n19624), .C1(n24733), .C2(n19564), .A(
        n22101), .ZN(n22096) );
  OAI22_X1 U21950 ( .A1(n21123), .A2(n24727), .B1(n20775), .B2(n24721), .ZN(
        n22101) );
  AOI221_X1 U21951 ( .B1(n24740), .B2(n19623), .C1(n24734), .C2(n19563), .A(
        n22082), .ZN(n22077) );
  OAI22_X1 U21952 ( .A1(n21050), .A2(n24728), .B1(n20654), .B2(n24722), .ZN(
        n22082) );
  AOI221_X1 U21953 ( .B1(n24740), .B2(n19622), .C1(n24734), .C2(n19562), .A(
        n22063), .ZN(n22058) );
  OAI22_X1 U21954 ( .A1(n21049), .A2(n24728), .B1(n20653), .B2(n24722), .ZN(
        n22063) );
  AOI221_X1 U21955 ( .B1(n24740), .B2(n19621), .C1(n24734), .C2(n19561), .A(
        n22044), .ZN(n22039) );
  OAI22_X1 U21956 ( .A1(n21048), .A2(n24728), .B1(n20652), .B2(n24722), .ZN(
        n22044) );
  AOI221_X1 U21957 ( .B1(n24740), .B2(n19620), .C1(n24734), .C2(n19560), .A(
        n22025), .ZN(n22020) );
  OAI22_X1 U21958 ( .A1(n21047), .A2(n24728), .B1(n20651), .B2(n24722), .ZN(
        n22025) );
  AOI221_X1 U21959 ( .B1(n24740), .B2(n19619), .C1(n24734), .C2(n19559), .A(
        n22006), .ZN(n22001) );
  OAI22_X1 U21960 ( .A1(n21046), .A2(n24728), .B1(n20650), .B2(n24722), .ZN(
        n22006) );
  AOI221_X1 U21961 ( .B1(n24740), .B2(n19618), .C1(n24734), .C2(n19558), .A(
        n21987), .ZN(n21982) );
  OAI22_X1 U21962 ( .A1(n21045), .A2(n24728), .B1(n20649), .B2(n24722), .ZN(
        n21987) );
  AOI221_X1 U21963 ( .B1(n24740), .B2(n19617), .C1(n24734), .C2(n19557), .A(
        n21968), .ZN(n21963) );
  OAI22_X1 U21964 ( .A1(n21044), .A2(n24728), .B1(n20648), .B2(n24722), .ZN(
        n21968) );
  AOI221_X1 U21965 ( .B1(n24740), .B2(n19616), .C1(n24734), .C2(n19556), .A(
        n21949), .ZN(n21944) );
  OAI22_X1 U21966 ( .A1(n21043), .A2(n24728), .B1(n20647), .B2(n24722), .ZN(
        n21949) );
  AOI221_X1 U21967 ( .B1(n24740), .B2(n19615), .C1(n24734), .C2(n19555), .A(
        n21930), .ZN(n21925) );
  OAI22_X1 U21968 ( .A1(n21042), .A2(n24728), .B1(n20646), .B2(n24722), .ZN(
        n21930) );
  AOI221_X1 U21969 ( .B1(n24740), .B2(n19614), .C1(n24734), .C2(n19554), .A(
        n21911), .ZN(n21906) );
  OAI22_X1 U21970 ( .A1(n21041), .A2(n24728), .B1(n20645), .B2(n24722), .ZN(
        n21911) );
  AOI221_X1 U21971 ( .B1(n24740), .B2(n19613), .C1(n24734), .C2(n19553), .A(
        n21892), .ZN(n21887) );
  OAI22_X1 U21972 ( .A1(n21040), .A2(n24728), .B1(n20644), .B2(n24722), .ZN(
        n21892) );
  AOI221_X1 U21973 ( .B1(n24740), .B2(n19612), .C1(n24734), .C2(n19552), .A(
        n21873), .ZN(n21868) );
  OAI22_X1 U21974 ( .A1(n21039), .A2(n24728), .B1(n20643), .B2(n24722), .ZN(
        n21873) );
  AOI221_X1 U21975 ( .B1(n24741), .B2(n19611), .C1(n24735), .C2(n19551), .A(
        n21854), .ZN(n21849) );
  OAI22_X1 U21976 ( .A1(n21038), .A2(n24729), .B1(n20642), .B2(n24723), .ZN(
        n21854) );
  AOI221_X1 U21977 ( .B1(n24741), .B2(n19610), .C1(n24735), .C2(n19550), .A(
        n21835), .ZN(n21830) );
  OAI22_X1 U21978 ( .A1(n21037), .A2(n24729), .B1(n20641), .B2(n24723), .ZN(
        n21835) );
  AOI221_X1 U21979 ( .B1(n24741), .B2(n19609), .C1(n24735), .C2(n19549), .A(
        n21816), .ZN(n21811) );
  OAI22_X1 U21980 ( .A1(n21036), .A2(n24729), .B1(n20640), .B2(n24723), .ZN(
        n21816) );
  AOI221_X1 U21981 ( .B1(n24741), .B2(n19608), .C1(n24735), .C2(n19548), .A(
        n21797), .ZN(n21792) );
  OAI22_X1 U21982 ( .A1(n21035), .A2(n24729), .B1(n20639), .B2(n24723), .ZN(
        n21797) );
  AOI221_X1 U21983 ( .B1(n24741), .B2(n19607), .C1(n24735), .C2(n19547), .A(
        n21778), .ZN(n21773) );
  OAI22_X1 U21984 ( .A1(n21034), .A2(n24729), .B1(n20638), .B2(n24723), .ZN(
        n21778) );
  AOI221_X1 U21985 ( .B1(n24741), .B2(n19606), .C1(n24735), .C2(n19546), .A(
        n21759), .ZN(n21754) );
  OAI22_X1 U21986 ( .A1(n21033), .A2(n24729), .B1(n20637), .B2(n24723), .ZN(
        n21759) );
  AOI221_X1 U21987 ( .B1(n24741), .B2(n19605), .C1(n24735), .C2(n19545), .A(
        n21740), .ZN(n21735) );
  OAI22_X1 U21988 ( .A1(n21032), .A2(n24729), .B1(n20636), .B2(n24723), .ZN(
        n21740) );
  AOI221_X1 U21989 ( .B1(n24741), .B2(n19604), .C1(n24735), .C2(n19544), .A(
        n21721), .ZN(n21716) );
  OAI22_X1 U21990 ( .A1(n21031), .A2(n24729), .B1(n20635), .B2(n24723), .ZN(
        n21721) );
  AOI221_X1 U21991 ( .B1(n24741), .B2(n19603), .C1(n24735), .C2(n19543), .A(
        n21702), .ZN(n21697) );
  OAI22_X1 U21992 ( .A1(n21030), .A2(n24729), .B1(n20634), .B2(n24723), .ZN(
        n21702) );
  AOI221_X1 U21993 ( .B1(n24741), .B2(n19602), .C1(n24735), .C2(n19542), .A(
        n21683), .ZN(n21678) );
  OAI22_X1 U21994 ( .A1(n21029), .A2(n24729), .B1(n20633), .B2(n24723), .ZN(
        n21683) );
  AOI221_X1 U21995 ( .B1(n24741), .B2(n19601), .C1(n24735), .C2(n19541), .A(
        n21664), .ZN(n21659) );
  OAI22_X1 U21996 ( .A1(n21028), .A2(n24729), .B1(n20632), .B2(n24723), .ZN(
        n21664) );
  AOI221_X1 U21997 ( .B1(n24741), .B2(n19600), .C1(n24735), .C2(n19540), .A(
        n21645), .ZN(n21640) );
  OAI22_X1 U21998 ( .A1(n21027), .A2(n24729), .B1(n20631), .B2(n24723), .ZN(
        n21645) );
  AOI221_X1 U21999 ( .B1(n24742), .B2(n19599), .C1(n24736), .C2(n19539), .A(
        n21626), .ZN(n21621) );
  OAI22_X1 U22000 ( .A1(n21026), .A2(n24730), .B1(n20630), .B2(n24724), .ZN(
        n21626) );
  AOI221_X1 U22001 ( .B1(n24742), .B2(n19598), .C1(n24736), .C2(n19538), .A(
        n21607), .ZN(n21602) );
  OAI22_X1 U22002 ( .A1(n21025), .A2(n24730), .B1(n20629), .B2(n24724), .ZN(
        n21607) );
  AOI221_X1 U22003 ( .B1(n24742), .B2(n19597), .C1(n24736), .C2(n19537), .A(
        n21588), .ZN(n21583) );
  OAI22_X1 U22004 ( .A1(n21024), .A2(n24730), .B1(n20628), .B2(n24724), .ZN(
        n21588) );
  AOI221_X1 U22005 ( .B1(n24742), .B2(n19596), .C1(n24736), .C2(n19536), .A(
        n21569), .ZN(n21564) );
  OAI22_X1 U22006 ( .A1(n21023), .A2(n24730), .B1(n20627), .B2(n24724), .ZN(
        n21569) );
  AOI221_X1 U22007 ( .B1(n24742), .B2(n19595), .C1(n24736), .C2(n19535), .A(
        n21550), .ZN(n21545) );
  OAI22_X1 U22008 ( .A1(n21022), .A2(n24730), .B1(n20626), .B2(n24724), .ZN(
        n21550) );
  AOI221_X1 U22009 ( .B1(n24742), .B2(n19594), .C1(n24736), .C2(n19534), .A(
        n21531), .ZN(n21526) );
  OAI22_X1 U22010 ( .A1(n21021), .A2(n24730), .B1(n20625), .B2(n24724), .ZN(
        n21531) );
  AOI221_X1 U22011 ( .B1(n24742), .B2(n19593), .C1(n24736), .C2(n19533), .A(
        n21512), .ZN(n21507) );
  OAI22_X1 U22012 ( .A1(n21020), .A2(n24730), .B1(n20624), .B2(n24724), .ZN(
        n21512) );
  AOI221_X1 U22013 ( .B1(n24742), .B2(n19592), .C1(n24736), .C2(n19532), .A(
        n21493), .ZN(n21488) );
  OAI22_X1 U22014 ( .A1(n21019), .A2(n24730), .B1(n20623), .B2(n24724), .ZN(
        n21493) );
  AOI221_X1 U22015 ( .B1(n24742), .B2(n19591), .C1(n24736), .C2(n19531), .A(
        n21474), .ZN(n21469) );
  OAI22_X1 U22016 ( .A1(n21018), .A2(n24730), .B1(n20622), .B2(n24724), .ZN(
        n21474) );
  AOI221_X1 U22017 ( .B1(n24742), .B2(n19590), .C1(n24736), .C2(n19530), .A(
        n21455), .ZN(n21450) );
  OAI22_X1 U22018 ( .A1(n21017), .A2(n24730), .B1(n20621), .B2(n24724), .ZN(
        n21455) );
  AOI221_X1 U22019 ( .B1(n24742), .B2(n19589), .C1(n24736), .C2(n19529), .A(
        n21436), .ZN(n21431) );
  OAI22_X1 U22020 ( .A1(n21016), .A2(n24730), .B1(n20620), .B2(n24724), .ZN(
        n21436) );
  AOI221_X1 U22021 ( .B1(n24742), .B2(n19588), .C1(n24736), .C2(n19528), .A(
        n21417), .ZN(n21412) );
  OAI22_X1 U22022 ( .A1(n21015), .A2(n24730), .B1(n20619), .B2(n24724), .ZN(
        n21417) );
  AOI221_X1 U22023 ( .B1(n24743), .B2(n20156), .C1(n24737), .C2(n19527), .A(
        n21398), .ZN(n21393) );
  OAI22_X1 U22024 ( .A1(n20546), .A2(n24731), .B1(n20517), .B2(n24725), .ZN(
        n21398) );
  AOI221_X1 U22025 ( .B1(n24647), .B2(n17652), .C1(n24641), .C2(n24208), .A(
        n21406), .ZN(n21401) );
  OAI22_X1 U22026 ( .A1(n20525), .A2(n24635), .B1(n20542), .B2(n24629), .ZN(
        n21406) );
  AOI221_X1 U22027 ( .B1(n24743), .B2(n20155), .C1(n24737), .C2(n19526), .A(
        n21379), .ZN(n21374) );
  OAI22_X1 U22028 ( .A1(n20545), .A2(n24731), .B1(n20516), .B2(n24725), .ZN(
        n21379) );
  AOI221_X1 U22029 ( .B1(n24647), .B2(n17655), .C1(n24641), .C2(n24209), .A(
        n21387), .ZN(n21382) );
  OAI22_X1 U22030 ( .A1(n20524), .A2(n24635), .B1(n20541), .B2(n24629), .ZN(
        n21387) );
  AOI221_X1 U22031 ( .B1(n24743), .B2(n20154), .C1(n24737), .C2(n19525), .A(
        n21360), .ZN(n21355) );
  OAI22_X1 U22032 ( .A1(n20544), .A2(n24731), .B1(n20515), .B2(n24725), .ZN(
        n21360) );
  AOI221_X1 U22033 ( .B1(n24647), .B2(n17658), .C1(n24641), .C2(n24210), .A(
        n21368), .ZN(n21363) );
  OAI22_X1 U22034 ( .A1(n20523), .A2(n24635), .B1(n20540), .B2(n24629), .ZN(
        n21368) );
  AOI221_X1 U22035 ( .B1(n24743), .B2(n20153), .C1(n24737), .C2(n19524), .A(
        n21319), .ZN(n21304) );
  OAI22_X1 U22036 ( .A1(n20543), .A2(n24731), .B1(n20514), .B2(n24725), .ZN(
        n21319) );
  AOI221_X1 U22037 ( .B1(n24647), .B2(n17661), .C1(n24641), .C2(n24211), .A(
        n21343), .ZN(n21328) );
  OAI22_X1 U22038 ( .A1(n20522), .A2(n24635), .B1(n20539), .B2(n24629), .ZN(
        n21343) );
  AOI221_X1 U22039 ( .B1(n24714), .B2(n20025), .C1(n24708), .C2(n20049), .A(
        n22547), .ZN(n22532) );
  OAI22_X1 U22040 ( .A1(n20505), .A2(n24702), .B1(n20822), .B2(n24696), .ZN(
        n22547) );
  AOI221_X1 U22041 ( .B1(n24618), .B2(n17540), .C1(n24612), .C2(n7709), .A(
        n22559), .ZN(n22548) );
  OAI22_X1 U22042 ( .A1(n20445), .A2(n24606), .B1(n20397), .B2(n24600), .ZN(
        n22559) );
  AOI221_X1 U22043 ( .B1(n24714), .B2(n20024), .C1(n24708), .C2(n20048), .A(
        n22520), .ZN(n22513) );
  OAI22_X1 U22044 ( .A1(n20504), .A2(n24702), .B1(n20821), .B2(n24696), .ZN(
        n22520) );
  AOI221_X1 U22045 ( .B1(n24618), .B2(n17543), .C1(n24612), .C2(n7708), .A(
        n22528), .ZN(n22521) );
  OAI22_X1 U22046 ( .A1(n20444), .A2(n24606), .B1(n20396), .B2(n24600), .ZN(
        n22528) );
  AOI221_X1 U22047 ( .B1(n24714), .B2(n20023), .C1(n24708), .C2(n20047), .A(
        n22501), .ZN(n22494) );
  OAI22_X1 U22048 ( .A1(n20503), .A2(n24702), .B1(n20820), .B2(n24696), .ZN(
        n22501) );
  AOI221_X1 U22049 ( .B1(n24618), .B2(n17546), .C1(n24612), .C2(n7707), .A(
        n22509), .ZN(n22502) );
  OAI22_X1 U22050 ( .A1(n20443), .A2(n24606), .B1(n20395), .B2(n24600), .ZN(
        n22509) );
  AOI221_X1 U22051 ( .B1(n24714), .B2(n20022), .C1(n24708), .C2(n20046), .A(
        n22482), .ZN(n22475) );
  OAI22_X1 U22052 ( .A1(n20502), .A2(n24702), .B1(n20819), .B2(n24696), .ZN(
        n22482) );
  AOI221_X1 U22053 ( .B1(n24618), .B2(n17549), .C1(n24612), .C2(n7706), .A(
        n22490), .ZN(n22483) );
  OAI22_X1 U22054 ( .A1(n20442), .A2(n24606), .B1(n20394), .B2(n24600), .ZN(
        n22490) );
  AOI221_X1 U22055 ( .B1(n24714), .B2(n20021), .C1(n24708), .C2(n20045), .A(
        n22463), .ZN(n22456) );
  OAI22_X1 U22056 ( .A1(n20501), .A2(n24702), .B1(n20818), .B2(n24696), .ZN(
        n22463) );
  AOI221_X1 U22057 ( .B1(n24618), .B2(n17552), .C1(n24612), .C2(n7705), .A(
        n22471), .ZN(n22464) );
  OAI22_X1 U22058 ( .A1(n20441), .A2(n24606), .B1(n20393), .B2(n24600), .ZN(
        n22471) );
  AOI221_X1 U22059 ( .B1(n24714), .B2(n20020), .C1(n24708), .C2(n20044), .A(
        n22444), .ZN(n22437) );
  OAI22_X1 U22060 ( .A1(n20500), .A2(n24702), .B1(n20817), .B2(n24696), .ZN(
        n22444) );
  AOI221_X1 U22061 ( .B1(n24618), .B2(n17555), .C1(n24612), .C2(n7704), .A(
        n22452), .ZN(n22445) );
  OAI22_X1 U22062 ( .A1(n20440), .A2(n24606), .B1(n20392), .B2(n24600), .ZN(
        n22452) );
  AOI221_X1 U22063 ( .B1(n24714), .B2(n20019), .C1(n24708), .C2(n20043), .A(
        n22425), .ZN(n22418) );
  OAI22_X1 U22064 ( .A1(n20499), .A2(n24702), .B1(n20816), .B2(n24696), .ZN(
        n22425) );
  AOI221_X1 U22065 ( .B1(n24618), .B2(n17558), .C1(n24612), .C2(n7703), .A(
        n22433), .ZN(n22426) );
  OAI22_X1 U22066 ( .A1(n20439), .A2(n24606), .B1(n20391), .B2(n24600), .ZN(
        n22433) );
  AOI221_X1 U22067 ( .B1(n24714), .B2(n20018), .C1(n24708), .C2(n20042), .A(
        n22406), .ZN(n22399) );
  OAI22_X1 U22068 ( .A1(n20498), .A2(n24702), .B1(n20815), .B2(n24696), .ZN(
        n22406) );
  AOI221_X1 U22069 ( .B1(n24618), .B2(n17561), .C1(n24612), .C2(n7702), .A(
        n22414), .ZN(n22407) );
  OAI22_X1 U22070 ( .A1(n20438), .A2(n24606), .B1(n20390), .B2(n24600), .ZN(
        n22414) );
  AOI221_X1 U22071 ( .B1(n24714), .B2(n20017), .C1(n24708), .C2(n20041), .A(
        n22387), .ZN(n22380) );
  OAI22_X1 U22072 ( .A1(n20497), .A2(n24702), .B1(n20814), .B2(n24696), .ZN(
        n22387) );
  AOI221_X1 U22073 ( .B1(n24618), .B2(n17564), .C1(n24612), .C2(n7701), .A(
        n22395), .ZN(n22388) );
  OAI22_X1 U22074 ( .A1(n20437), .A2(n24606), .B1(n20389), .B2(n24600), .ZN(
        n22395) );
  AOI221_X1 U22075 ( .B1(n24714), .B2(n20016), .C1(n24708), .C2(n20040), .A(
        n22368), .ZN(n22361) );
  OAI22_X1 U22076 ( .A1(n20496), .A2(n24702), .B1(n20813), .B2(n24696), .ZN(
        n22368) );
  AOI221_X1 U22077 ( .B1(n24618), .B2(n17567), .C1(n24612), .C2(n7700), .A(
        n22376), .ZN(n22369) );
  OAI22_X1 U22078 ( .A1(n20436), .A2(n24606), .B1(n20388), .B2(n24600), .ZN(
        n22376) );
  AOI221_X1 U22079 ( .B1(n24714), .B2(n20015), .C1(n24708), .C2(n20039), .A(
        n22349), .ZN(n22342) );
  OAI22_X1 U22080 ( .A1(n20495), .A2(n24702), .B1(n20812), .B2(n24696), .ZN(
        n22349) );
  AOI221_X1 U22081 ( .B1(n24618), .B2(n17570), .C1(n24612), .C2(n7699), .A(
        n22357), .ZN(n22350) );
  OAI22_X1 U22082 ( .A1(n20435), .A2(n24606), .B1(n20387), .B2(n24600), .ZN(
        n22357) );
  AOI221_X1 U22083 ( .B1(n24714), .B2(n20014), .C1(n24708), .C2(n20038), .A(
        n22330), .ZN(n22323) );
  OAI22_X1 U22084 ( .A1(n20494), .A2(n24702), .B1(n20811), .B2(n24696), .ZN(
        n22330) );
  AOI221_X1 U22085 ( .B1(n24618), .B2(n17573), .C1(n24612), .C2(n7698), .A(
        n22338), .ZN(n22331) );
  OAI22_X1 U22086 ( .A1(n20434), .A2(n24606), .B1(n20386), .B2(n24600), .ZN(
        n22338) );
  AOI221_X1 U22087 ( .B1(n24715), .B2(n20013), .C1(n24709), .C2(n20037), .A(
        n22311), .ZN(n22304) );
  OAI22_X1 U22088 ( .A1(n20493), .A2(n24703), .B1(n20810), .B2(n24697), .ZN(
        n22311) );
  AOI221_X1 U22089 ( .B1(n24619), .B2(n17576), .C1(n24613), .C2(n7697), .A(
        n22319), .ZN(n22312) );
  OAI22_X1 U22090 ( .A1(n20433), .A2(n24607), .B1(n20385), .B2(n24601), .ZN(
        n22319) );
  AOI221_X1 U22091 ( .B1(n24715), .B2(n20012), .C1(n24709), .C2(n20036), .A(
        n22292), .ZN(n22285) );
  OAI22_X1 U22092 ( .A1(n20492), .A2(n24703), .B1(n20809), .B2(n24697), .ZN(
        n22292) );
  AOI221_X1 U22093 ( .B1(n24619), .B2(n17579), .C1(n24613), .C2(n7696), .A(
        n22300), .ZN(n22293) );
  OAI22_X1 U22094 ( .A1(n20432), .A2(n24607), .B1(n20384), .B2(n24601), .ZN(
        n22300) );
  AOI221_X1 U22095 ( .B1(n24715), .B2(n20011), .C1(n24709), .C2(n20035), .A(
        n22273), .ZN(n22266) );
  OAI22_X1 U22096 ( .A1(n20491), .A2(n24703), .B1(n20808), .B2(n24697), .ZN(
        n22273) );
  AOI221_X1 U22097 ( .B1(n24619), .B2(n17582), .C1(n24613), .C2(n7695), .A(
        n22281), .ZN(n22274) );
  OAI22_X1 U22098 ( .A1(n20431), .A2(n24607), .B1(n20383), .B2(n24601), .ZN(
        n22281) );
  AOI221_X1 U22099 ( .B1(n24715), .B2(n20010), .C1(n24709), .C2(n20034), .A(
        n22254), .ZN(n22247) );
  OAI22_X1 U22100 ( .A1(n20490), .A2(n24703), .B1(n20807), .B2(n24697), .ZN(
        n22254) );
  AOI221_X1 U22101 ( .B1(n24619), .B2(n17585), .C1(n24613), .C2(n7694), .A(
        n22262), .ZN(n22255) );
  OAI22_X1 U22102 ( .A1(n20430), .A2(n24607), .B1(n20382), .B2(n24601), .ZN(
        n22262) );
  AOI221_X1 U22103 ( .B1(n24715), .B2(n20009), .C1(n24709), .C2(n20033), .A(
        n22235), .ZN(n22228) );
  OAI22_X1 U22104 ( .A1(n20489), .A2(n24703), .B1(n20806), .B2(n24697), .ZN(
        n22235) );
  AOI221_X1 U22105 ( .B1(n24619), .B2(n17588), .C1(n24613), .C2(n7693), .A(
        n22243), .ZN(n22236) );
  OAI22_X1 U22106 ( .A1(n20429), .A2(n24607), .B1(n20381), .B2(n24601), .ZN(
        n22243) );
  AOI221_X1 U22107 ( .B1(n24715), .B2(n20008), .C1(n24709), .C2(n20032), .A(
        n22216), .ZN(n22209) );
  OAI22_X1 U22108 ( .A1(n20488), .A2(n24703), .B1(n20805), .B2(n24697), .ZN(
        n22216) );
  AOI221_X1 U22109 ( .B1(n24619), .B2(n17591), .C1(n24613), .C2(n7692), .A(
        n22224), .ZN(n22217) );
  OAI22_X1 U22110 ( .A1(n20428), .A2(n24607), .B1(n20380), .B2(n24601), .ZN(
        n22224) );
  AOI221_X1 U22111 ( .B1(n24715), .B2(n20007), .C1(n24709), .C2(n20031), .A(
        n22197), .ZN(n22190) );
  OAI22_X1 U22112 ( .A1(n20487), .A2(n24703), .B1(n20804), .B2(n24697), .ZN(
        n22197) );
  AOI221_X1 U22113 ( .B1(n24619), .B2(n17594), .C1(n24613), .C2(n7691), .A(
        n22205), .ZN(n22198) );
  OAI22_X1 U22114 ( .A1(n20427), .A2(n24607), .B1(n20379), .B2(n24601), .ZN(
        n22205) );
  AOI221_X1 U22115 ( .B1(n24715), .B2(n20006), .C1(n24709), .C2(n20030), .A(
        n22178), .ZN(n22171) );
  OAI22_X1 U22116 ( .A1(n20486), .A2(n24703), .B1(n20803), .B2(n24697), .ZN(
        n22178) );
  AOI221_X1 U22117 ( .B1(n24619), .B2(n17597), .C1(n24613), .C2(n7690), .A(
        n22186), .ZN(n22179) );
  OAI22_X1 U22118 ( .A1(n20426), .A2(n24607), .B1(n20378), .B2(n24601), .ZN(
        n22186) );
  AOI221_X1 U22119 ( .B1(n24715), .B2(n20005), .C1(n24709), .C2(n20029), .A(
        n22159), .ZN(n22152) );
  OAI22_X1 U22120 ( .A1(n20485), .A2(n24703), .B1(n20802), .B2(n24697), .ZN(
        n22159) );
  AOI221_X1 U22121 ( .B1(n24619), .B2(n17600), .C1(n24613), .C2(n7689), .A(
        n22167), .ZN(n22160) );
  OAI22_X1 U22122 ( .A1(n20425), .A2(n24607), .B1(n20377), .B2(n24601), .ZN(
        n22167) );
  AOI221_X1 U22123 ( .B1(n24715), .B2(n20004), .C1(n24709), .C2(n20028), .A(
        n22140), .ZN(n22133) );
  OAI22_X1 U22124 ( .A1(n20484), .A2(n24703), .B1(n20801), .B2(n24697), .ZN(
        n22140) );
  AOI221_X1 U22125 ( .B1(n24619), .B2(n17603), .C1(n24613), .C2(n7688), .A(
        n22148), .ZN(n22141) );
  OAI22_X1 U22126 ( .A1(n20424), .A2(n24607), .B1(n20376), .B2(n24601), .ZN(
        n22148) );
  AOI221_X1 U22127 ( .B1(n24715), .B2(n20003), .C1(n24709), .C2(n20027), .A(
        n22121), .ZN(n22114) );
  OAI22_X1 U22128 ( .A1(n20483), .A2(n24703), .B1(n20800), .B2(n24697), .ZN(
        n22121) );
  AOI221_X1 U22129 ( .B1(n24619), .B2(n17606), .C1(n24613), .C2(n7687), .A(
        n22129), .ZN(n22122) );
  OAI22_X1 U22130 ( .A1(n20423), .A2(n24607), .B1(n20375), .B2(n24601), .ZN(
        n22129) );
  AOI221_X1 U22131 ( .B1(n24715), .B2(n20002), .C1(n24709), .C2(n20026), .A(
        n22102), .ZN(n22095) );
  OAI22_X1 U22132 ( .A1(n20482), .A2(n24703), .B1(n20799), .B2(n24697), .ZN(
        n22102) );
  AOI221_X1 U22133 ( .B1(n24619), .B2(n17609), .C1(n24613), .C2(n7686), .A(
        n22110), .ZN(n22103) );
  OAI22_X1 U22134 ( .A1(n20422), .A2(n24607), .B1(n20374), .B2(n24601), .ZN(
        n22110) );
  AOI221_X1 U22135 ( .B1(n24716), .B2(n19857), .C1(n24710), .C2(n19893), .A(
        n22083), .ZN(n22076) );
  OAI22_X1 U22136 ( .A1(n20481), .A2(n24704), .B1(n20690), .B2(n24698), .ZN(
        n22083) );
  AOI221_X1 U22137 ( .B1(n24620), .B2(n17612), .C1(n24614), .C2(n7685), .A(
        n22091), .ZN(n22084) );
  OAI22_X1 U22138 ( .A1(n20373), .A2(n24608), .B1(n20301), .B2(n24602), .ZN(
        n22091) );
  AOI221_X1 U22139 ( .B1(n24716), .B2(n19856), .C1(n24710), .C2(n19892), .A(
        n22064), .ZN(n22057) );
  OAI22_X1 U22140 ( .A1(n20480), .A2(n24704), .B1(n20689), .B2(n24698), .ZN(
        n22064) );
  AOI221_X1 U22141 ( .B1(n24620), .B2(n17615), .C1(n24614), .C2(n7684), .A(
        n22072), .ZN(n22065) );
  OAI22_X1 U22142 ( .A1(n20372), .A2(n24608), .B1(n20300), .B2(n24602), .ZN(
        n22072) );
  AOI221_X1 U22143 ( .B1(n24716), .B2(n19855), .C1(n24710), .C2(n19891), .A(
        n22045), .ZN(n22038) );
  OAI22_X1 U22144 ( .A1(n20479), .A2(n24704), .B1(n20688), .B2(n24698), .ZN(
        n22045) );
  AOI221_X1 U22145 ( .B1(n24620), .B2(n17618), .C1(n24614), .C2(n7683), .A(
        n22053), .ZN(n22046) );
  OAI22_X1 U22146 ( .A1(n20371), .A2(n24608), .B1(n20299), .B2(n24602), .ZN(
        n22053) );
  AOI221_X1 U22147 ( .B1(n24716), .B2(n19854), .C1(n24710), .C2(n19890), .A(
        n22026), .ZN(n22019) );
  OAI22_X1 U22148 ( .A1(n20478), .A2(n24704), .B1(n20687), .B2(n24698), .ZN(
        n22026) );
  AOI221_X1 U22149 ( .B1(n24620), .B2(n17621), .C1(n24614), .C2(n7682), .A(
        n22034), .ZN(n22027) );
  OAI22_X1 U22150 ( .A1(n20370), .A2(n24608), .B1(n20298), .B2(n24602), .ZN(
        n22034) );
  AOI221_X1 U22151 ( .B1(n24716), .B2(n19853), .C1(n24710), .C2(n19889), .A(
        n22007), .ZN(n22000) );
  OAI22_X1 U22152 ( .A1(n20477), .A2(n24704), .B1(n20686), .B2(n24698), .ZN(
        n22007) );
  AOI221_X1 U22153 ( .B1(n24620), .B2(n17624), .C1(n24614), .C2(n7681), .A(
        n22015), .ZN(n22008) );
  OAI22_X1 U22154 ( .A1(n20369), .A2(n24608), .B1(n20297), .B2(n24602), .ZN(
        n22015) );
  AOI221_X1 U22155 ( .B1(n24716), .B2(n19852), .C1(n24710), .C2(n19888), .A(
        n21988), .ZN(n21981) );
  OAI22_X1 U22156 ( .A1(n20476), .A2(n24704), .B1(n20685), .B2(n24698), .ZN(
        n21988) );
  AOI221_X1 U22157 ( .B1(n24620), .B2(n17471), .C1(n24614), .C2(n20144), .A(
        n21996), .ZN(n21989) );
  OAI22_X1 U22158 ( .A1(n20368), .A2(n24608), .B1(n20296), .B2(n24602), .ZN(
        n21996) );
  AOI221_X1 U22159 ( .B1(n24716), .B2(n19851), .C1(n24710), .C2(n19887), .A(
        n21969), .ZN(n21962) );
  OAI22_X1 U22160 ( .A1(n20475), .A2(n24704), .B1(n20684), .B2(n24698), .ZN(
        n21969) );
  AOI221_X1 U22161 ( .B1(n24620), .B2(n17474), .C1(n24614), .C2(n20143), .A(
        n21977), .ZN(n21970) );
  OAI22_X1 U22162 ( .A1(n20367), .A2(n24608), .B1(n20295), .B2(n24602), .ZN(
        n21977) );
  AOI221_X1 U22163 ( .B1(n24716), .B2(n19850), .C1(n24710), .C2(n19886), .A(
        n21950), .ZN(n21943) );
  OAI22_X1 U22164 ( .A1(n20474), .A2(n24704), .B1(n20683), .B2(n24698), .ZN(
        n21950) );
  AOI221_X1 U22165 ( .B1(n24620), .B2(n17477), .C1(n24614), .C2(n20142), .A(
        n21958), .ZN(n21951) );
  OAI22_X1 U22166 ( .A1(n20366), .A2(n24608), .B1(n20294), .B2(n24602), .ZN(
        n21958) );
  AOI221_X1 U22167 ( .B1(n24716), .B2(n19849), .C1(n24710), .C2(n19885), .A(
        n21931), .ZN(n21924) );
  OAI22_X1 U22168 ( .A1(n20473), .A2(n24704), .B1(n20682), .B2(n24698), .ZN(
        n21931) );
  AOI221_X1 U22169 ( .B1(n24620), .B2(n17480), .C1(n24614), .C2(n20141), .A(
        n21939), .ZN(n21932) );
  OAI22_X1 U22170 ( .A1(n20365), .A2(n24608), .B1(n20293), .B2(n24602), .ZN(
        n21939) );
  AOI221_X1 U22171 ( .B1(n24716), .B2(n19848), .C1(n24710), .C2(n19884), .A(
        n21912), .ZN(n21905) );
  OAI22_X1 U22172 ( .A1(n20472), .A2(n24704), .B1(n20681), .B2(n24698), .ZN(
        n21912) );
  AOI221_X1 U22173 ( .B1(n24620), .B2(n17483), .C1(n24614), .C2(n20140), .A(
        n21920), .ZN(n21913) );
  OAI22_X1 U22174 ( .A1(n20364), .A2(n24608), .B1(n20292), .B2(n24602), .ZN(
        n21920) );
  AOI221_X1 U22175 ( .B1(n24716), .B2(n19847), .C1(n24710), .C2(n19883), .A(
        n21893), .ZN(n21886) );
  OAI22_X1 U22176 ( .A1(n20471), .A2(n24704), .B1(n20680), .B2(n24698), .ZN(
        n21893) );
  AOI221_X1 U22177 ( .B1(n24620), .B2(n17486), .C1(n24614), .C2(n20139), .A(
        n21901), .ZN(n21894) );
  OAI22_X1 U22178 ( .A1(n20363), .A2(n24608), .B1(n20291), .B2(n24602), .ZN(
        n21901) );
  AOI221_X1 U22179 ( .B1(n24716), .B2(n19846), .C1(n24710), .C2(n19882), .A(
        n21874), .ZN(n21867) );
  OAI22_X1 U22180 ( .A1(n20470), .A2(n24704), .B1(n20679), .B2(n24698), .ZN(
        n21874) );
  AOI221_X1 U22181 ( .B1(n24620), .B2(n17489), .C1(n24614), .C2(n20133), .A(
        n21882), .ZN(n21875) );
  OAI22_X1 U22182 ( .A1(n20362), .A2(n24608), .B1(n20290), .B2(n24602), .ZN(
        n21882) );
  AOI221_X1 U22183 ( .B1(n24717), .B2(n19845), .C1(n24711), .C2(n19881), .A(
        n21855), .ZN(n21848) );
  OAI22_X1 U22184 ( .A1(n20469), .A2(n24705), .B1(n20678), .B2(n24699), .ZN(
        n21855) );
  AOI221_X1 U22185 ( .B1(n24621), .B2(n17492), .C1(n24615), .C2(n20138), .A(
        n21863), .ZN(n21856) );
  OAI22_X1 U22186 ( .A1(n20361), .A2(n24609), .B1(n20289), .B2(n24603), .ZN(
        n21863) );
  AOI221_X1 U22187 ( .B1(n24717), .B2(n19844), .C1(n24711), .C2(n19880), .A(
        n21836), .ZN(n21829) );
  OAI22_X1 U22188 ( .A1(n20468), .A2(n24705), .B1(n20677), .B2(n24699), .ZN(
        n21836) );
  AOI221_X1 U22189 ( .B1(n24621), .B2(n17495), .C1(n24615), .C2(n20137), .A(
        n21844), .ZN(n21837) );
  OAI22_X1 U22190 ( .A1(n20360), .A2(n24609), .B1(n20288), .B2(n24603), .ZN(
        n21844) );
  AOI221_X1 U22191 ( .B1(n24717), .B2(n19843), .C1(n24711), .C2(n19879), .A(
        n21817), .ZN(n21810) );
  OAI22_X1 U22192 ( .A1(n20467), .A2(n24705), .B1(n20676), .B2(n24699), .ZN(
        n21817) );
  AOI221_X1 U22193 ( .B1(n24621), .B2(n17498), .C1(n24615), .C2(n20136), .A(
        n21825), .ZN(n21818) );
  OAI22_X1 U22194 ( .A1(n20359), .A2(n24609), .B1(n20287), .B2(n24603), .ZN(
        n21825) );
  AOI221_X1 U22195 ( .B1(n24717), .B2(n19842), .C1(n24711), .C2(n19878), .A(
        n21798), .ZN(n21791) );
  OAI22_X1 U22196 ( .A1(n20466), .A2(n24705), .B1(n20675), .B2(n24699), .ZN(
        n21798) );
  AOI221_X1 U22197 ( .B1(n24621), .B2(n17501), .C1(n24615), .C2(n20132), .A(
        n21806), .ZN(n21799) );
  OAI22_X1 U22198 ( .A1(n20358), .A2(n24609), .B1(n20286), .B2(n24603), .ZN(
        n21806) );
  AOI221_X1 U22199 ( .B1(n24717), .B2(n19841), .C1(n24711), .C2(n19877), .A(
        n21779), .ZN(n21772) );
  OAI22_X1 U22200 ( .A1(n20465), .A2(n24705), .B1(n20674), .B2(n24699), .ZN(
        n21779) );
  AOI221_X1 U22201 ( .B1(n24621), .B2(n17504), .C1(n24615), .C2(n20135), .A(
        n21787), .ZN(n21780) );
  OAI22_X1 U22202 ( .A1(n20357), .A2(n24609), .B1(n20285), .B2(n24603), .ZN(
        n21787) );
  AOI221_X1 U22203 ( .B1(n24717), .B2(n19840), .C1(n24711), .C2(n19876), .A(
        n21760), .ZN(n21753) );
  OAI22_X1 U22204 ( .A1(n20464), .A2(n24705), .B1(n20673), .B2(n24699), .ZN(
        n21760) );
  AOI221_X1 U22205 ( .B1(n24621), .B2(n17507), .C1(n24615), .C2(n20131), .A(
        n21768), .ZN(n21761) );
  OAI22_X1 U22206 ( .A1(n20356), .A2(n24609), .B1(n20284), .B2(n24603), .ZN(
        n21768) );
  AOI221_X1 U22207 ( .B1(n24717), .B2(n19839), .C1(n24711), .C2(n19875), .A(
        n21741), .ZN(n21734) );
  OAI22_X1 U22208 ( .A1(n20463), .A2(n24705), .B1(n20672), .B2(n24699), .ZN(
        n21741) );
  AOI221_X1 U22209 ( .B1(n24621), .B2(n17510), .C1(n24615), .C2(n20134), .A(
        n21749), .ZN(n21742) );
  OAI22_X1 U22210 ( .A1(n20355), .A2(n24609), .B1(n20283), .B2(n24603), .ZN(
        n21749) );
  AOI221_X1 U22211 ( .B1(n24717), .B2(n19838), .C1(n24711), .C2(n19874), .A(
        n21722), .ZN(n21715) );
  OAI22_X1 U22212 ( .A1(n20462), .A2(n24705), .B1(n20671), .B2(n24699), .ZN(
        n21722) );
  AOI221_X1 U22213 ( .B1(n24621), .B2(n17513), .C1(n24615), .C2(n20130), .A(
        n21730), .ZN(n21723) );
  OAI22_X1 U22214 ( .A1(n20354), .A2(n24609), .B1(n20282), .B2(n24603), .ZN(
        n21730) );
  AOI221_X1 U22215 ( .B1(n24717), .B2(n19837), .C1(n24711), .C2(n19873), .A(
        n21703), .ZN(n21696) );
  OAI22_X1 U22216 ( .A1(n20461), .A2(n24705), .B1(n20670), .B2(n24699), .ZN(
        n21703) );
  AOI221_X1 U22217 ( .B1(n24621), .B2(n17516), .C1(n24615), .C2(n20129), .A(
        n21711), .ZN(n21704) );
  OAI22_X1 U22218 ( .A1(n20353), .A2(n24609), .B1(n20281), .B2(n24603), .ZN(
        n21711) );
  AOI221_X1 U22219 ( .B1(n24717), .B2(n19836), .C1(n24711), .C2(n19872), .A(
        n21684), .ZN(n21677) );
  OAI22_X1 U22220 ( .A1(n20460), .A2(n24705), .B1(n20669), .B2(n24699), .ZN(
        n21684) );
  AOI221_X1 U22221 ( .B1(n24621), .B2(n17519), .C1(n24615), .C2(n20128), .A(
        n21692), .ZN(n21685) );
  OAI22_X1 U22222 ( .A1(n20352), .A2(n24609), .B1(n20280), .B2(n24603), .ZN(
        n21692) );
  AOI221_X1 U22223 ( .B1(n24717), .B2(n19835), .C1(n24711), .C2(n19871), .A(
        n21665), .ZN(n21658) );
  OAI22_X1 U22224 ( .A1(n20459), .A2(n24705), .B1(n20668), .B2(n24699), .ZN(
        n21665) );
  AOI221_X1 U22225 ( .B1(n24621), .B2(n17522), .C1(n24615), .C2(n20127), .A(
        n21673), .ZN(n21666) );
  OAI22_X1 U22226 ( .A1(n20351), .A2(n24609), .B1(n20279), .B2(n24603), .ZN(
        n21673) );
  AOI221_X1 U22227 ( .B1(n24717), .B2(n19834), .C1(n24711), .C2(n19870), .A(
        n21646), .ZN(n21639) );
  OAI22_X1 U22228 ( .A1(n20458), .A2(n24705), .B1(n20667), .B2(n24699), .ZN(
        n21646) );
  AOI221_X1 U22229 ( .B1(n24621), .B2(n17525), .C1(n24615), .C2(n20126), .A(
        n21654), .ZN(n21647) );
  OAI22_X1 U22230 ( .A1(n20350), .A2(n24609), .B1(n20278), .B2(n24603), .ZN(
        n21654) );
  AOI221_X1 U22231 ( .B1(n24718), .B2(n19833), .C1(n24712), .C2(n19869), .A(
        n21627), .ZN(n21620) );
  OAI22_X1 U22232 ( .A1(n20457), .A2(n24706), .B1(n20666), .B2(n24700), .ZN(
        n21627) );
  AOI221_X1 U22233 ( .B1(n24622), .B2(n17528), .C1(n24616), .C2(n20125), .A(
        n21635), .ZN(n21628) );
  OAI22_X1 U22234 ( .A1(n20349), .A2(n24610), .B1(n20277), .B2(n24604), .ZN(
        n21635) );
  AOI221_X1 U22235 ( .B1(n24718), .B2(n19832), .C1(n24712), .C2(n19868), .A(
        n21608), .ZN(n21601) );
  OAI22_X1 U22236 ( .A1(n20456), .A2(n24706), .B1(n20665), .B2(n24700), .ZN(
        n21608) );
  AOI221_X1 U22237 ( .B1(n24622), .B2(n17531), .C1(n24616), .C2(n20124), .A(
        n21616), .ZN(n21609) );
  OAI22_X1 U22238 ( .A1(n20348), .A2(n24610), .B1(n20276), .B2(n24604), .ZN(
        n21616) );
  AOI221_X1 U22239 ( .B1(n24718), .B2(n19831), .C1(n24712), .C2(n19867), .A(
        n21589), .ZN(n21582) );
  OAI22_X1 U22240 ( .A1(n20455), .A2(n24706), .B1(n20664), .B2(n24700), .ZN(
        n21589) );
  AOI221_X1 U22241 ( .B1(n24622), .B2(n17534), .C1(n24616), .C2(n20123), .A(
        n21597), .ZN(n21590) );
  OAI22_X1 U22242 ( .A1(n20347), .A2(n24610), .B1(n20275), .B2(n24604), .ZN(
        n21597) );
  AOI221_X1 U22243 ( .B1(n24718), .B2(n19830), .C1(n24712), .C2(n19866), .A(
        n21570), .ZN(n21563) );
  OAI22_X1 U22244 ( .A1(n20454), .A2(n24706), .B1(n20663), .B2(n24700), .ZN(
        n21570) );
  AOI221_X1 U22245 ( .B1(n24622), .B2(n17537), .C1(n24616), .C2(n20122), .A(
        n21578), .ZN(n21571) );
  OAI22_X1 U22246 ( .A1(n20346), .A2(n24610), .B1(n20274), .B2(n24604), .ZN(
        n21578) );
  AOI221_X1 U22247 ( .B1(n24718), .B2(n19829), .C1(n24712), .C2(n19865), .A(
        n21551), .ZN(n21544) );
  OAI22_X1 U22248 ( .A1(n20453), .A2(n24706), .B1(n20662), .B2(n24700), .ZN(
        n21551) );
  AOI221_X1 U22249 ( .B1(n24622), .B2(n17627), .C1(n24616), .C2(n7657), .A(
        n21559), .ZN(n21552) );
  OAI22_X1 U22250 ( .A1(n20345), .A2(n24610), .B1(n20273), .B2(n24604), .ZN(
        n21559) );
  AOI221_X1 U22251 ( .B1(n24718), .B2(n19828), .C1(n24712), .C2(n19864), .A(
        n21532), .ZN(n21525) );
  OAI22_X1 U22252 ( .A1(n20452), .A2(n24706), .B1(n20661), .B2(n24700), .ZN(
        n21532) );
  AOI221_X1 U22253 ( .B1(n24622), .B2(n17630), .C1(n24616), .C2(n7656), .A(
        n21540), .ZN(n21533) );
  OAI22_X1 U22254 ( .A1(n20344), .A2(n24610), .B1(n20272), .B2(n24604), .ZN(
        n21540) );
  AOI221_X1 U22255 ( .B1(n24718), .B2(n19827), .C1(n24712), .C2(n19863), .A(
        n21513), .ZN(n21506) );
  OAI22_X1 U22256 ( .A1(n20451), .A2(n24706), .B1(n20660), .B2(n24700), .ZN(
        n21513) );
  AOI221_X1 U22257 ( .B1(n24622), .B2(n17633), .C1(n24616), .C2(n7655), .A(
        n21521), .ZN(n21514) );
  OAI22_X1 U22258 ( .A1(n20343), .A2(n24610), .B1(n20271), .B2(n24604), .ZN(
        n21521) );
  AOI221_X1 U22259 ( .B1(n24718), .B2(n19826), .C1(n24712), .C2(n19862), .A(
        n21494), .ZN(n21487) );
  OAI22_X1 U22260 ( .A1(n20450), .A2(n24706), .B1(n20659), .B2(n24700), .ZN(
        n21494) );
  AOI221_X1 U22261 ( .B1(n24622), .B2(n17636), .C1(n24616), .C2(n7654), .A(
        n21502), .ZN(n21495) );
  OAI22_X1 U22262 ( .A1(n20342), .A2(n24610), .B1(n20270), .B2(n24604), .ZN(
        n21502) );
  AOI221_X1 U22263 ( .B1(n24718), .B2(n19825), .C1(n24712), .C2(n19861), .A(
        n21475), .ZN(n21468) );
  OAI22_X1 U22264 ( .A1(n20449), .A2(n24706), .B1(n20658), .B2(n24700), .ZN(
        n21475) );
  AOI221_X1 U22265 ( .B1(n24622), .B2(n17639), .C1(n24616), .C2(n7653), .A(
        n21483), .ZN(n21476) );
  OAI22_X1 U22266 ( .A1(n20341), .A2(n24610), .B1(n20269), .B2(n24604), .ZN(
        n21483) );
  AOI221_X1 U22267 ( .B1(n24718), .B2(n19824), .C1(n24712), .C2(n19860), .A(
        n21456), .ZN(n21449) );
  OAI22_X1 U22268 ( .A1(n20448), .A2(n24706), .B1(n20657), .B2(n24700), .ZN(
        n21456) );
  AOI221_X1 U22269 ( .B1(n24622), .B2(n17642), .C1(n24616), .C2(n7652), .A(
        n21464), .ZN(n21457) );
  OAI22_X1 U22270 ( .A1(n20340), .A2(n24610), .B1(n20268), .B2(n24604), .ZN(
        n21464) );
  AOI221_X1 U22271 ( .B1(n24718), .B2(n19823), .C1(n24712), .C2(n19859), .A(
        n21437), .ZN(n21430) );
  OAI22_X1 U22272 ( .A1(n20447), .A2(n24706), .B1(n20656), .B2(n24700), .ZN(
        n21437) );
  AOI221_X1 U22273 ( .B1(n24622), .B2(n17645), .C1(n24616), .C2(n7651), .A(
        n21445), .ZN(n21438) );
  OAI22_X1 U22274 ( .A1(n20339), .A2(n24610), .B1(n20267), .B2(n24604), .ZN(
        n21445) );
  AOI221_X1 U22275 ( .B1(n24718), .B2(n19822), .C1(n24712), .C2(n19858), .A(
        n21418), .ZN(n21411) );
  OAI22_X1 U22276 ( .A1(n20446), .A2(n24706), .B1(n20655), .B2(n24700), .ZN(
        n21418) );
  AOI221_X1 U22277 ( .B1(n24622), .B2(n17648), .C1(n24616), .C2(n7650), .A(
        n21426), .ZN(n21419) );
  OAI22_X1 U22278 ( .A1(n20338), .A2(n24610), .B1(n20266), .B2(n24604), .ZN(
        n21426) );
  AOI221_X1 U22279 ( .B1(n24719), .B2(n19805), .C1(n24713), .C2(n19809), .A(
        n21399), .ZN(n21392) );
  OAI22_X1 U22280 ( .A1(n20265), .A2(n24707), .B1(n20521), .B2(n24701), .ZN(
        n21399) );
  AOI221_X1 U22281 ( .B1(n24623), .B2(n17651), .C1(n24617), .C2(n7649), .A(
        n21407), .ZN(n21400) );
  OAI22_X1 U22282 ( .A1(n20261), .A2(n24611), .B1(n20253), .B2(n24605), .ZN(
        n21407) );
  AOI221_X1 U22283 ( .B1(n24719), .B2(n19804), .C1(n24713), .C2(n19808), .A(
        n21380), .ZN(n21373) );
  OAI22_X1 U22284 ( .A1(n20264), .A2(n24707), .B1(n20520), .B2(n24701), .ZN(
        n21380) );
  AOI221_X1 U22285 ( .B1(n24623), .B2(n17654), .C1(n24617), .C2(n7648), .A(
        n21388), .ZN(n21381) );
  OAI22_X1 U22286 ( .A1(n20260), .A2(n24611), .B1(n20252), .B2(n24605), .ZN(
        n21388) );
  AOI221_X1 U22287 ( .B1(n24719), .B2(n19803), .C1(n24713), .C2(n19807), .A(
        n21361), .ZN(n21354) );
  OAI22_X1 U22288 ( .A1(n20263), .A2(n24707), .B1(n20519), .B2(n24701), .ZN(
        n21361) );
  AOI221_X1 U22289 ( .B1(n24623), .B2(n17657), .C1(n24617), .C2(n7647), .A(
        n21369), .ZN(n21362) );
  OAI22_X1 U22290 ( .A1(n20259), .A2(n24611), .B1(n20251), .B2(n24605), .ZN(
        n21369) );
  AOI221_X1 U22291 ( .B1(n24719), .B2(n19802), .C1(n24713), .C2(n19806), .A(
        n21324), .ZN(n21303) );
  OAI22_X1 U22292 ( .A1(n20262), .A2(n24707), .B1(n20518), .B2(n24701), .ZN(
        n21324) );
  AOI221_X1 U22293 ( .B1(n24623), .B2(n17660), .C1(n24617), .C2(n7646), .A(
        n21348), .ZN(n21327) );
  OAI22_X1 U22294 ( .A1(n20258), .A2(n24611), .B1(n20250), .B2(n24605), .ZN(
        n21348) );
  OAI221_X1 U22295 ( .B1(n7346), .B2(n24597), .C1(n7474), .C2(n24591), .A(
        n23016), .ZN(n23015) );
  AOI22_X1 U22296 ( .A1(n24585), .A2(n7989), .B1(n24579), .B2(n19547), .ZN(
        n23016) );
  OAI221_X1 U22297 ( .B1(n7344), .B2(n24597), .C1(n7472), .C2(n24591), .A(
        n22998), .ZN(n22997) );
  AOI22_X1 U22298 ( .A1(n24585), .A2(n7988), .B1(n24579), .B2(n19546), .ZN(
        n22998) );
  OAI221_X1 U22299 ( .B1(n7342), .B2(n24597), .C1(n7470), .C2(n24591), .A(
        n22980), .ZN(n22979) );
  AOI22_X1 U22300 ( .A1(n24585), .A2(n7987), .B1(n24579), .B2(n19545), .ZN(
        n22980) );
  OAI221_X1 U22301 ( .B1(n7340), .B2(n24597), .C1(n7468), .C2(n24591), .A(
        n22962), .ZN(n22961) );
  AOI22_X1 U22302 ( .A1(n24585), .A2(n7986), .B1(n24579), .B2(n19544), .ZN(
        n22962) );
  OAI221_X1 U22303 ( .B1(n7338), .B2(n24597), .C1(n7466), .C2(n24591), .A(
        n22944), .ZN(n22943) );
  AOI22_X1 U22304 ( .A1(n24585), .A2(n7985), .B1(n24579), .B2(n19543), .ZN(
        n22944) );
  OAI221_X1 U22305 ( .B1(n7336), .B2(n24597), .C1(n7464), .C2(n24591), .A(
        n22926), .ZN(n22925) );
  AOI22_X1 U22306 ( .A1(n24585), .A2(n7984), .B1(n24579), .B2(n19542), .ZN(
        n22926) );
  OAI221_X1 U22307 ( .B1(n7334), .B2(n24597), .C1(n7462), .C2(n24591), .A(
        n22908), .ZN(n22907) );
  AOI22_X1 U22308 ( .A1(n24585), .A2(n7983), .B1(n24579), .B2(n19541), .ZN(
        n22908) );
  OAI221_X1 U22309 ( .B1(n7332), .B2(n24597), .C1(n7460), .C2(n24591), .A(
        n22890), .ZN(n22889) );
  AOI22_X1 U22310 ( .A1(n24585), .A2(n7982), .B1(n24579), .B2(n19540), .ZN(
        n22890) );
  OAI221_X1 U22311 ( .B1(n7330), .B2(n24598), .C1(n7458), .C2(n24592), .A(
        n22872), .ZN(n22871) );
  AOI22_X1 U22312 ( .A1(n24586), .A2(n7981), .B1(n24580), .B2(n19539), .ZN(
        n22872) );
  OAI221_X1 U22313 ( .B1(n7328), .B2(n24598), .C1(n7456), .C2(n24592), .A(
        n22854), .ZN(n22853) );
  AOI22_X1 U22314 ( .A1(n24586), .A2(n7980), .B1(n24580), .B2(n19538), .ZN(
        n22854) );
  OAI221_X1 U22315 ( .B1(n7326), .B2(n24598), .C1(n7454), .C2(n24592), .A(
        n22836), .ZN(n22835) );
  AOI22_X1 U22316 ( .A1(n24586), .A2(n7979), .B1(n24580), .B2(n19537), .ZN(
        n22836) );
  OAI221_X1 U22317 ( .B1(n7324), .B2(n24598), .C1(n7452), .C2(n24592), .A(
        n22818), .ZN(n22817) );
  AOI22_X1 U22318 ( .A1(n24586), .A2(n7978), .B1(n24580), .B2(n19536), .ZN(
        n22818) );
  OAI221_X1 U22319 ( .B1(n7322), .B2(n24598), .C1(n7450), .C2(n24592), .A(
        n22800), .ZN(n22799) );
  AOI22_X1 U22320 ( .A1(n24586), .A2(n7977), .B1(n24580), .B2(n19535), .ZN(
        n22800) );
  OAI221_X1 U22321 ( .B1(n7320), .B2(n24598), .C1(n7448), .C2(n24592), .A(
        n22782), .ZN(n22781) );
  AOI22_X1 U22322 ( .A1(n24586), .A2(n7976), .B1(n24580), .B2(n19534), .ZN(
        n22782) );
  OAI221_X1 U22323 ( .B1(n7318), .B2(n24598), .C1(n7446), .C2(n24592), .A(
        n22764), .ZN(n22763) );
  AOI22_X1 U22324 ( .A1(n24586), .A2(n7975), .B1(n24580), .B2(n19533), .ZN(
        n22764) );
  OAI221_X1 U22325 ( .B1(n7316), .B2(n24598), .C1(n7444), .C2(n24592), .A(
        n22746), .ZN(n22745) );
  AOI22_X1 U22326 ( .A1(n24586), .A2(n7974), .B1(n24580), .B2(n19532), .ZN(
        n22746) );
  OAI221_X1 U22327 ( .B1(n7314), .B2(n24598), .C1(n7442), .C2(n24592), .A(
        n22728), .ZN(n22727) );
  AOI22_X1 U22328 ( .A1(n24586), .A2(n7973), .B1(n24580), .B2(n19531), .ZN(
        n22728) );
  OAI221_X1 U22329 ( .B1(n7312), .B2(n24598), .C1(n7440), .C2(n24592), .A(
        n22710), .ZN(n22709) );
  AOI22_X1 U22330 ( .A1(n24586), .A2(n7972), .B1(n24580), .B2(n19530), .ZN(
        n22710) );
  OAI221_X1 U22331 ( .B1(n7310), .B2(n24598), .C1(n7438), .C2(n24592), .A(
        n22692), .ZN(n22691) );
  AOI22_X1 U22332 ( .A1(n24586), .A2(n7971), .B1(n24580), .B2(n19529), .ZN(
        n22692) );
  OAI221_X1 U22333 ( .B1(n7308), .B2(n24598), .C1(n7436), .C2(n24592), .A(
        n22674), .ZN(n22673) );
  AOI22_X1 U22334 ( .A1(n24586), .A2(n7970), .B1(n24580), .B2(n19528), .ZN(
        n22674) );
  OAI221_X1 U22335 ( .B1(n7402), .B2(n24595), .C1(n7530), .C2(n24589), .A(
        n23520), .ZN(n23519) );
  AOI22_X1 U22336 ( .A1(n24583), .A2(n8017), .B1(n24577), .B2(n19575), .ZN(
        n23520) );
  OAI221_X1 U22337 ( .B1(n7400), .B2(n24595), .C1(n7528), .C2(n24589), .A(
        n23502), .ZN(n23501) );
  AOI22_X1 U22338 ( .A1(n24583), .A2(n8016), .B1(n24577), .B2(n19574), .ZN(
        n23502) );
  OAI221_X1 U22339 ( .B1(n7398), .B2(n24595), .C1(n7526), .C2(n24589), .A(
        n23484), .ZN(n23483) );
  AOI22_X1 U22340 ( .A1(n24583), .A2(n8015), .B1(n24577), .B2(n19573), .ZN(
        n23484) );
  OAI221_X1 U22341 ( .B1(n7396), .B2(n24595), .C1(n7524), .C2(n24589), .A(
        n23466), .ZN(n23465) );
  AOI22_X1 U22342 ( .A1(n24583), .A2(n8014), .B1(n24577), .B2(n19572), .ZN(
        n23466) );
  OAI221_X1 U22343 ( .B1(n7394), .B2(n24595), .C1(n7522), .C2(n24589), .A(
        n23448), .ZN(n23447) );
  AOI22_X1 U22344 ( .A1(n24583), .A2(n8013), .B1(n24577), .B2(n19571), .ZN(
        n23448) );
  OAI221_X1 U22345 ( .B1(n7392), .B2(n24595), .C1(n7520), .C2(n24589), .A(
        n23430), .ZN(n23429) );
  AOI22_X1 U22346 ( .A1(n24583), .A2(n8012), .B1(n24577), .B2(n19570), .ZN(
        n23430) );
  OAI221_X1 U22347 ( .B1(n7390), .B2(n24595), .C1(n7518), .C2(n24589), .A(
        n23412), .ZN(n23411) );
  AOI22_X1 U22348 ( .A1(n24583), .A2(n8011), .B1(n24577), .B2(n19569), .ZN(
        n23412) );
  OAI221_X1 U22349 ( .B1(n7388), .B2(n24595), .C1(n7516), .C2(n24589), .A(
        n23394), .ZN(n23393) );
  AOI22_X1 U22350 ( .A1(n24583), .A2(n8010), .B1(n24577), .B2(n19568), .ZN(
        n23394) );
  OAI221_X1 U22351 ( .B1(n7386), .B2(n24595), .C1(n7514), .C2(n24589), .A(
        n23376), .ZN(n23375) );
  AOI22_X1 U22352 ( .A1(n24583), .A2(n8009), .B1(n24577), .B2(n19567), .ZN(
        n23376) );
  OAI221_X1 U22353 ( .B1(n7384), .B2(n24595), .C1(n7512), .C2(n24589), .A(
        n23358), .ZN(n23357) );
  AOI22_X1 U22354 ( .A1(n24583), .A2(n8008), .B1(n24577), .B2(n19566), .ZN(
        n23358) );
  OAI221_X1 U22355 ( .B1(n7382), .B2(n24595), .C1(n7510), .C2(n24589), .A(
        n23340), .ZN(n23339) );
  AOI22_X1 U22356 ( .A1(n24583), .A2(n8007), .B1(n24577), .B2(n19565), .ZN(
        n23340) );
  OAI221_X1 U22357 ( .B1(n7380), .B2(n24595), .C1(n7508), .C2(n24589), .A(
        n23322), .ZN(n23321) );
  AOI22_X1 U22358 ( .A1(n24583), .A2(n8006), .B1(n24577), .B2(n19564), .ZN(
        n23322) );
  OAI221_X1 U22359 ( .B1(n7378), .B2(n24596), .C1(n7506), .C2(n24590), .A(
        n23304), .ZN(n23303) );
  AOI22_X1 U22360 ( .A1(n24584), .A2(n8005), .B1(n24578), .B2(n19563), .ZN(
        n23304) );
  OAI221_X1 U22361 ( .B1(n7376), .B2(n24596), .C1(n7504), .C2(n24590), .A(
        n23286), .ZN(n23285) );
  AOI22_X1 U22362 ( .A1(n24584), .A2(n8004), .B1(n24578), .B2(n19562), .ZN(
        n23286) );
  OAI221_X1 U22363 ( .B1(n7374), .B2(n24596), .C1(n7502), .C2(n24590), .A(
        n23268), .ZN(n23267) );
  AOI22_X1 U22364 ( .A1(n24584), .A2(n8003), .B1(n24578), .B2(n19561), .ZN(
        n23268) );
  OAI221_X1 U22365 ( .B1(n7372), .B2(n24596), .C1(n7500), .C2(n24590), .A(
        n23250), .ZN(n23249) );
  AOI22_X1 U22366 ( .A1(n24584), .A2(n8002), .B1(n24578), .B2(n19560), .ZN(
        n23250) );
  OAI221_X1 U22367 ( .B1(n7370), .B2(n24596), .C1(n7498), .C2(n24590), .A(
        n23232), .ZN(n23231) );
  AOI22_X1 U22368 ( .A1(n24584), .A2(n8001), .B1(n24578), .B2(n19559), .ZN(
        n23232) );
  OAI221_X1 U22369 ( .B1(n7368), .B2(n24596), .C1(n7496), .C2(n24590), .A(
        n23214), .ZN(n23213) );
  AOI22_X1 U22370 ( .A1(n24584), .A2(n8000), .B1(n24578), .B2(n19558), .ZN(
        n23214) );
  OAI221_X1 U22371 ( .B1(n7366), .B2(n24596), .C1(n7494), .C2(n24590), .A(
        n23196), .ZN(n23195) );
  AOI22_X1 U22372 ( .A1(n24584), .A2(n7999), .B1(n24578), .B2(n19557), .ZN(
        n23196) );
  OAI221_X1 U22373 ( .B1(n7364), .B2(n24596), .C1(n7492), .C2(n24590), .A(
        n23178), .ZN(n23177) );
  AOI22_X1 U22374 ( .A1(n24584), .A2(n7998), .B1(n24578), .B2(n19556), .ZN(
        n23178) );
  OAI221_X1 U22375 ( .B1(n7362), .B2(n24596), .C1(n7490), .C2(n24590), .A(
        n23160), .ZN(n23159) );
  AOI22_X1 U22376 ( .A1(n24584), .A2(n7997), .B1(n24578), .B2(n19555), .ZN(
        n23160) );
  OAI221_X1 U22377 ( .B1(n7360), .B2(n24596), .C1(n7488), .C2(n24590), .A(
        n23142), .ZN(n23141) );
  AOI22_X1 U22378 ( .A1(n24584), .A2(n7996), .B1(n24578), .B2(n19554), .ZN(
        n23142) );
  OAI221_X1 U22379 ( .B1(n7358), .B2(n24596), .C1(n7486), .C2(n24590), .A(
        n23124), .ZN(n23123) );
  AOI22_X1 U22380 ( .A1(n24584), .A2(n7995), .B1(n24578), .B2(n19553), .ZN(
        n23124) );
  OAI221_X1 U22381 ( .B1(n7356), .B2(n24596), .C1(n7484), .C2(n24590), .A(
        n23106), .ZN(n23105) );
  AOI22_X1 U22382 ( .A1(n24584), .A2(n7994), .B1(n24578), .B2(n19552), .ZN(
        n23106) );
  OAI221_X1 U22383 ( .B1(n7354), .B2(n24597), .C1(n7482), .C2(n24591), .A(
        n23088), .ZN(n23087) );
  AOI22_X1 U22384 ( .A1(n24585), .A2(n7993), .B1(n24579), .B2(n19551), .ZN(
        n23088) );
  OAI221_X1 U22385 ( .B1(n7352), .B2(n24597), .C1(n7480), .C2(n24591), .A(
        n23070), .ZN(n23069) );
  AOI22_X1 U22386 ( .A1(n24585), .A2(n7992), .B1(n24579), .B2(n19550), .ZN(
        n23070) );
  OAI221_X1 U22387 ( .B1(n7350), .B2(n24597), .C1(n7478), .C2(n24591), .A(
        n23052), .ZN(n23051) );
  AOI22_X1 U22388 ( .A1(n24585), .A2(n7991), .B1(n24579), .B2(n19549), .ZN(
        n23052) );
  OAI221_X1 U22389 ( .B1(n7348), .B2(n24597), .C1(n7476), .C2(n24591), .A(
        n23034), .ZN(n23033) );
  AOI22_X1 U22390 ( .A1(n24585), .A2(n7990), .B1(n24579), .B2(n19548), .ZN(
        n23034) );
  OAI221_X1 U22391 ( .B1(n7306), .B2(n24599), .C1(n7434), .C2(n24593), .A(
        n22656), .ZN(n22655) );
  AOI22_X1 U22392 ( .A1(n24587), .A2(n7969), .B1(n24581), .B2(n19527), .ZN(
        n22656) );
  OAI221_X1 U22393 ( .B1(n7304), .B2(n24599), .C1(n7432), .C2(n24593), .A(
        n22638), .ZN(n22637) );
  AOI22_X1 U22394 ( .A1(n24587), .A2(n7968), .B1(n24581), .B2(n19526), .ZN(
        n22638) );
  OAI221_X1 U22395 ( .B1(n7302), .B2(n24599), .C1(n7430), .C2(n24593), .A(
        n22620), .ZN(n22619) );
  AOI22_X1 U22396 ( .A1(n24587), .A2(n7967), .B1(n24581), .B2(n19525), .ZN(
        n22620) );
  OAI221_X1 U22397 ( .B1(n7300), .B2(n24599), .C1(n7428), .C2(n24593), .A(
        n22570), .ZN(n22567) );
  AOI22_X1 U22398 ( .A1(n24587), .A2(n7966), .B1(n24581), .B2(n19524), .ZN(
        n22570) );
  OAI221_X1 U22399 ( .B1(n7426), .B2(n24594), .C1(n7554), .C2(n24588), .A(
        n23736), .ZN(n23735) );
  AOI22_X1 U22400 ( .A1(n24582), .A2(n8029), .B1(n24576), .B2(n19587), .ZN(
        n23736) );
  OAI221_X1 U22401 ( .B1(n7424), .B2(n24594), .C1(n7552), .C2(n24588), .A(
        n23718), .ZN(n23717) );
  AOI22_X1 U22402 ( .A1(n24582), .A2(n8028), .B1(n24576), .B2(n19586), .ZN(
        n23718) );
  OAI221_X1 U22403 ( .B1(n7422), .B2(n24594), .C1(n7550), .C2(n24588), .A(
        n23700), .ZN(n23699) );
  AOI22_X1 U22404 ( .A1(n24582), .A2(n8027), .B1(n24576), .B2(n19585), .ZN(
        n23700) );
  OAI221_X1 U22405 ( .B1(n7420), .B2(n24594), .C1(n7548), .C2(n24588), .A(
        n23682), .ZN(n23681) );
  AOI22_X1 U22406 ( .A1(n24582), .A2(n8026), .B1(n24576), .B2(n19584), .ZN(
        n23682) );
  OAI221_X1 U22407 ( .B1(n7418), .B2(n24594), .C1(n7546), .C2(n24588), .A(
        n23664), .ZN(n23663) );
  AOI22_X1 U22408 ( .A1(n24582), .A2(n8025), .B1(n24576), .B2(n19583), .ZN(
        n23664) );
  OAI221_X1 U22409 ( .B1(n7416), .B2(n24594), .C1(n7544), .C2(n24588), .A(
        n23646), .ZN(n23645) );
  AOI22_X1 U22410 ( .A1(n24582), .A2(n8024), .B1(n24576), .B2(n19582), .ZN(
        n23646) );
  OAI221_X1 U22411 ( .B1(n7414), .B2(n24594), .C1(n7542), .C2(n24588), .A(
        n23628), .ZN(n23627) );
  AOI22_X1 U22412 ( .A1(n24582), .A2(n8023), .B1(n24576), .B2(n19581), .ZN(
        n23628) );
  OAI221_X1 U22413 ( .B1(n7412), .B2(n24594), .C1(n7540), .C2(n24588), .A(
        n23610), .ZN(n23609) );
  AOI22_X1 U22414 ( .A1(n24582), .A2(n8022), .B1(n24576), .B2(n19580), .ZN(
        n23610) );
  OAI221_X1 U22415 ( .B1(n7410), .B2(n24594), .C1(n7538), .C2(n24588), .A(
        n23592), .ZN(n23591) );
  AOI22_X1 U22416 ( .A1(n24582), .A2(n8021), .B1(n24576), .B2(n19579), .ZN(
        n23592) );
  OAI221_X1 U22417 ( .B1(n7408), .B2(n24594), .C1(n7536), .C2(n24588), .A(
        n23574), .ZN(n23573) );
  AOI22_X1 U22418 ( .A1(n24582), .A2(n8020), .B1(n24576), .B2(n19578), .ZN(
        n23574) );
  OAI221_X1 U22419 ( .B1(n7406), .B2(n24594), .C1(n7534), .C2(n24588), .A(
        n23556), .ZN(n23555) );
  AOI22_X1 U22420 ( .A1(n24582), .A2(n8019), .B1(n24576), .B2(n19577), .ZN(
        n23556) );
  OAI221_X1 U22421 ( .B1(n7404), .B2(n24594), .C1(n7532), .C2(n24588), .A(
        n23538), .ZN(n23537) );
  AOI22_X1 U22422 ( .A1(n24582), .A2(n8018), .B1(n24576), .B2(n19576), .ZN(
        n23538) );
  OAI22_X1 U22423 ( .A1(n20152), .A2(n24407), .B1(n8869), .B2(n24401), .ZN(
        n22665) );
  OAI22_X1 U22424 ( .A1(n9124), .A2(n24431), .B1(n9125), .B2(n24425), .ZN(
        n22664) );
  OAI22_X1 U22425 ( .A1(n20151), .A2(n24407), .B1(n8867), .B2(n24401), .ZN(
        n22647) );
  OAI22_X1 U22426 ( .A1(n9122), .A2(n24431), .B1(n9123), .B2(n24425), .ZN(
        n22646) );
  OAI22_X1 U22427 ( .A1(n20150), .A2(n24407), .B1(n8865), .B2(n24401), .ZN(
        n22629) );
  OAI22_X1 U22428 ( .A1(n9120), .A2(n24431), .B1(n9121), .B2(n24425), .ZN(
        n22628) );
  OAI22_X1 U22429 ( .A1(n20149), .A2(n24407), .B1(n8863), .B2(n24401), .ZN(
        n22609) );
  OAI22_X1 U22430 ( .A1(n9118), .A2(n24431), .B1(n9119), .B2(n24425), .ZN(
        n22604) );
  OAI22_X1 U22431 ( .A1(n19667), .A2(n24405), .B1(n8909), .B2(n24399), .ZN(
        n23025) );
  OAI22_X1 U22432 ( .A1(n9164), .A2(n24429), .B1(n9165), .B2(n24423), .ZN(
        n23024) );
  OAI22_X1 U22433 ( .A1(n19666), .A2(n24405), .B1(n8907), .B2(n24399), .ZN(
        n23007) );
  OAI22_X1 U22434 ( .A1(n9162), .A2(n24429), .B1(n9163), .B2(n24423), .ZN(
        n23006) );
  OAI22_X1 U22435 ( .A1(n19665), .A2(n24405), .B1(n8905), .B2(n24399), .ZN(
        n22989) );
  OAI22_X1 U22436 ( .A1(n9160), .A2(n24429), .B1(n9161), .B2(n24423), .ZN(
        n22988) );
  OAI22_X1 U22437 ( .A1(n19664), .A2(n24405), .B1(n8903), .B2(n24399), .ZN(
        n22971) );
  OAI22_X1 U22438 ( .A1(n9158), .A2(n24429), .B1(n9159), .B2(n24423), .ZN(
        n22970) );
  OAI22_X1 U22439 ( .A1(n19663), .A2(n24405), .B1(n8901), .B2(n24399), .ZN(
        n22953) );
  OAI22_X1 U22440 ( .A1(n9156), .A2(n24429), .B1(n9157), .B2(n24423), .ZN(
        n22952) );
  OAI22_X1 U22441 ( .A1(n19662), .A2(n24405), .B1(n8899), .B2(n24399), .ZN(
        n22935) );
  OAI22_X1 U22442 ( .A1(n9154), .A2(n24429), .B1(n9155), .B2(n24423), .ZN(
        n22934) );
  OAI22_X1 U22443 ( .A1(n19661), .A2(n24405), .B1(n8897), .B2(n24399), .ZN(
        n22917) );
  OAI22_X1 U22444 ( .A1(n9152), .A2(n24429), .B1(n9153), .B2(n24423), .ZN(
        n22916) );
  OAI22_X1 U22445 ( .A1(n19660), .A2(n24405), .B1(n8895), .B2(n24399), .ZN(
        n22899) );
  OAI22_X1 U22446 ( .A1(n9150), .A2(n24429), .B1(n9151), .B2(n24423), .ZN(
        n22898) );
  OAI22_X1 U22447 ( .A1(n19659), .A2(n24406), .B1(n8893), .B2(n24400), .ZN(
        n22881) );
  OAI22_X1 U22448 ( .A1(n9148), .A2(n24430), .B1(n9149), .B2(n24424), .ZN(
        n22880) );
  OAI22_X1 U22449 ( .A1(n19658), .A2(n24406), .B1(n8891), .B2(n24400), .ZN(
        n22863) );
  OAI22_X1 U22450 ( .A1(n9146), .A2(n24430), .B1(n9147), .B2(n24424), .ZN(
        n22862) );
  OAI22_X1 U22451 ( .A1(n19657), .A2(n24406), .B1(n8889), .B2(n24400), .ZN(
        n22845) );
  OAI22_X1 U22452 ( .A1(n9144), .A2(n24430), .B1(n9145), .B2(n24424), .ZN(
        n22844) );
  OAI22_X1 U22453 ( .A1(n19656), .A2(n24406), .B1(n8887), .B2(n24400), .ZN(
        n22827) );
  OAI22_X1 U22454 ( .A1(n9142), .A2(n24430), .B1(n9143), .B2(n24424), .ZN(
        n22826) );
  OAI22_X1 U22455 ( .A1(n19655), .A2(n24406), .B1(n8885), .B2(n24400), .ZN(
        n22809) );
  OAI22_X1 U22456 ( .A1(n9140), .A2(n24430), .B1(n9141), .B2(n24424), .ZN(
        n22808) );
  OAI22_X1 U22457 ( .A1(n19654), .A2(n24406), .B1(n8883), .B2(n24400), .ZN(
        n22791) );
  OAI22_X1 U22458 ( .A1(n9138), .A2(n24430), .B1(n9139), .B2(n24424), .ZN(
        n22790) );
  OAI22_X1 U22459 ( .A1(n19653), .A2(n24406), .B1(n8881), .B2(n24400), .ZN(
        n22773) );
  OAI22_X1 U22460 ( .A1(n9136), .A2(n24430), .B1(n9137), .B2(n24424), .ZN(
        n22772) );
  OAI22_X1 U22461 ( .A1(n19652), .A2(n24406), .B1(n8879), .B2(n24400), .ZN(
        n22755) );
  OAI22_X1 U22462 ( .A1(n9134), .A2(n24430), .B1(n9135), .B2(n24424), .ZN(
        n22754) );
  OAI22_X1 U22463 ( .A1(n19651), .A2(n24406), .B1(n8877), .B2(n24400), .ZN(
        n22737) );
  OAI22_X1 U22464 ( .A1(n9132), .A2(n24430), .B1(n9133), .B2(n24424), .ZN(
        n22736) );
  OAI22_X1 U22465 ( .A1(n19650), .A2(n24406), .B1(n8875), .B2(n24400), .ZN(
        n22719) );
  OAI22_X1 U22466 ( .A1(n9130), .A2(n24430), .B1(n9131), .B2(n24424), .ZN(
        n22718) );
  OAI22_X1 U22467 ( .A1(n19649), .A2(n24406), .B1(n8873), .B2(n24400), .ZN(
        n22701) );
  OAI22_X1 U22468 ( .A1(n9128), .A2(n24430), .B1(n9129), .B2(n24424), .ZN(
        n22700) );
  OAI22_X1 U22469 ( .A1(n19648), .A2(n24406), .B1(n8871), .B2(n24400), .ZN(
        n22683) );
  OAI22_X1 U22470 ( .A1(n9126), .A2(n24430), .B1(n9127), .B2(n24424), .ZN(
        n22682) );
  OAI22_X1 U22471 ( .A1(n19707), .A2(n24402), .B1(n8989), .B2(n24396), .ZN(
        n23763) );
  OAI22_X1 U22472 ( .A1(n9244), .A2(n24426), .B1(n9245), .B2(n24420), .ZN(
        n23762) );
  OAI22_X1 U22473 ( .A1(n19706), .A2(n24402), .B1(n8987), .B2(n24396), .ZN(
        n23727) );
  OAI22_X1 U22474 ( .A1(n9242), .A2(n24426), .B1(n9243), .B2(n24420), .ZN(
        n23726) );
  OAI22_X1 U22475 ( .A1(n19705), .A2(n24402), .B1(n8985), .B2(n24396), .ZN(
        n23709) );
  OAI22_X1 U22476 ( .A1(n9240), .A2(n24426), .B1(n9241), .B2(n24420), .ZN(
        n23708) );
  OAI22_X1 U22477 ( .A1(n19704), .A2(n24402), .B1(n8983), .B2(n24396), .ZN(
        n23691) );
  OAI22_X1 U22478 ( .A1(n9238), .A2(n24426), .B1(n9239), .B2(n24420), .ZN(
        n23690) );
  OAI22_X1 U22479 ( .A1(n19703), .A2(n24402), .B1(n8981), .B2(n24396), .ZN(
        n23673) );
  OAI22_X1 U22480 ( .A1(n9236), .A2(n24426), .B1(n9237), .B2(n24420), .ZN(
        n23672) );
  OAI22_X1 U22481 ( .A1(n19702), .A2(n24402), .B1(n8979), .B2(n24396), .ZN(
        n23655) );
  OAI22_X1 U22482 ( .A1(n9234), .A2(n24426), .B1(n9235), .B2(n24420), .ZN(
        n23654) );
  OAI22_X1 U22483 ( .A1(n19701), .A2(n24402), .B1(n8977), .B2(n24396), .ZN(
        n23637) );
  OAI22_X1 U22484 ( .A1(n9232), .A2(n24426), .B1(n9233), .B2(n24420), .ZN(
        n23636) );
  OAI22_X1 U22485 ( .A1(n19700), .A2(n24402), .B1(n8975), .B2(n24396), .ZN(
        n23619) );
  OAI22_X1 U22486 ( .A1(n9230), .A2(n24426), .B1(n9231), .B2(n24420), .ZN(
        n23618) );
  OAI22_X1 U22487 ( .A1(n19699), .A2(n24402), .B1(n8973), .B2(n24396), .ZN(
        n23601) );
  OAI22_X1 U22488 ( .A1(n9228), .A2(n24426), .B1(n9229), .B2(n24420), .ZN(
        n23600) );
  OAI22_X1 U22489 ( .A1(n19698), .A2(n24402), .B1(n8971), .B2(n24396), .ZN(
        n23583) );
  OAI22_X1 U22490 ( .A1(n9226), .A2(n24426), .B1(n9227), .B2(n24420), .ZN(
        n23582) );
  OAI22_X1 U22491 ( .A1(n19697), .A2(n24402), .B1(n8969), .B2(n24396), .ZN(
        n23565) );
  OAI22_X1 U22492 ( .A1(n9224), .A2(n24426), .B1(n9225), .B2(n24420), .ZN(
        n23564) );
  OAI22_X1 U22493 ( .A1(n19696), .A2(n24402), .B1(n8967), .B2(n24396), .ZN(
        n23547) );
  OAI22_X1 U22494 ( .A1(n9222), .A2(n24426), .B1(n9223), .B2(n24420), .ZN(
        n23546) );
  OAI22_X1 U22495 ( .A1(n19695), .A2(n24403), .B1(n8965), .B2(n24397), .ZN(
        n23529) );
  OAI22_X1 U22496 ( .A1(n9220), .A2(n24427), .B1(n9221), .B2(n24421), .ZN(
        n23528) );
  OAI22_X1 U22497 ( .A1(n19694), .A2(n24403), .B1(n8963), .B2(n24397), .ZN(
        n23511) );
  OAI22_X1 U22498 ( .A1(n9218), .A2(n24427), .B1(n9219), .B2(n24421), .ZN(
        n23510) );
  OAI22_X1 U22499 ( .A1(n19693), .A2(n24403), .B1(n8961), .B2(n24397), .ZN(
        n23493) );
  OAI22_X1 U22500 ( .A1(n9216), .A2(n24427), .B1(n9217), .B2(n24421), .ZN(
        n23492) );
  OAI22_X1 U22501 ( .A1(n19692), .A2(n24403), .B1(n8959), .B2(n24397), .ZN(
        n23475) );
  OAI22_X1 U22502 ( .A1(n9214), .A2(n24427), .B1(n9215), .B2(n24421), .ZN(
        n23474) );
  OAI22_X1 U22503 ( .A1(n19691), .A2(n24403), .B1(n8957), .B2(n24397), .ZN(
        n23457) );
  OAI22_X1 U22504 ( .A1(n9212), .A2(n24427), .B1(n9213), .B2(n24421), .ZN(
        n23456) );
  OAI22_X1 U22505 ( .A1(n19690), .A2(n24403), .B1(n8955), .B2(n24397), .ZN(
        n23439) );
  OAI22_X1 U22506 ( .A1(n9210), .A2(n24427), .B1(n9211), .B2(n24421), .ZN(
        n23438) );
  OAI22_X1 U22507 ( .A1(n19689), .A2(n24403), .B1(n8953), .B2(n24397), .ZN(
        n23421) );
  OAI22_X1 U22508 ( .A1(n9208), .A2(n24427), .B1(n9209), .B2(n24421), .ZN(
        n23420) );
  OAI22_X1 U22509 ( .A1(n19688), .A2(n24403), .B1(n8951), .B2(n24397), .ZN(
        n23403) );
  OAI22_X1 U22510 ( .A1(n9206), .A2(n24427), .B1(n9207), .B2(n24421), .ZN(
        n23402) );
  OAI22_X1 U22511 ( .A1(n19687), .A2(n24403), .B1(n8949), .B2(n24397), .ZN(
        n23385) );
  OAI22_X1 U22512 ( .A1(n9204), .A2(n24427), .B1(n9205), .B2(n24421), .ZN(
        n23384) );
  OAI22_X1 U22513 ( .A1(n19686), .A2(n24403), .B1(n8947), .B2(n24397), .ZN(
        n23367) );
  OAI22_X1 U22514 ( .A1(n9202), .A2(n24427), .B1(n9203), .B2(n24421), .ZN(
        n23366) );
  OAI22_X1 U22515 ( .A1(n19685), .A2(n24403), .B1(n8945), .B2(n24397), .ZN(
        n23349) );
  OAI22_X1 U22516 ( .A1(n9200), .A2(n24427), .B1(n9201), .B2(n24421), .ZN(
        n23348) );
  OAI22_X1 U22517 ( .A1(n19684), .A2(n24403), .B1(n8943), .B2(n24397), .ZN(
        n23331) );
  OAI22_X1 U22518 ( .A1(n9198), .A2(n24427), .B1(n9199), .B2(n24421), .ZN(
        n23330) );
  OAI22_X1 U22519 ( .A1(n19683), .A2(n24404), .B1(n8941), .B2(n24398), .ZN(
        n23313) );
  OAI22_X1 U22520 ( .A1(n9196), .A2(n24428), .B1(n9197), .B2(n24422), .ZN(
        n23312) );
  OAI22_X1 U22521 ( .A1(n19682), .A2(n24404), .B1(n8939), .B2(n24398), .ZN(
        n23295) );
  OAI22_X1 U22522 ( .A1(n9194), .A2(n24428), .B1(n9195), .B2(n24422), .ZN(
        n23294) );
  OAI22_X1 U22523 ( .A1(n19681), .A2(n24404), .B1(n8937), .B2(n24398), .ZN(
        n23277) );
  OAI22_X1 U22524 ( .A1(n9192), .A2(n24428), .B1(n9193), .B2(n24422), .ZN(
        n23276) );
  OAI22_X1 U22525 ( .A1(n19680), .A2(n24404), .B1(n8935), .B2(n24398), .ZN(
        n23259) );
  OAI22_X1 U22526 ( .A1(n9190), .A2(n24428), .B1(n9191), .B2(n24422), .ZN(
        n23258) );
  OAI22_X1 U22527 ( .A1(n19679), .A2(n24404), .B1(n8933), .B2(n24398), .ZN(
        n23241) );
  OAI22_X1 U22528 ( .A1(n9188), .A2(n24428), .B1(n9189), .B2(n24422), .ZN(
        n23240) );
  OAI22_X1 U22529 ( .A1(n19678), .A2(n24404), .B1(n8931), .B2(n24398), .ZN(
        n23223) );
  OAI22_X1 U22530 ( .A1(n9186), .A2(n24428), .B1(n9187), .B2(n24422), .ZN(
        n23222) );
  OAI22_X1 U22531 ( .A1(n19677), .A2(n24404), .B1(n8929), .B2(n24398), .ZN(
        n23205) );
  OAI22_X1 U22532 ( .A1(n9184), .A2(n24428), .B1(n9185), .B2(n24422), .ZN(
        n23204) );
  OAI22_X1 U22533 ( .A1(n19676), .A2(n24404), .B1(n8927), .B2(n24398), .ZN(
        n23187) );
  OAI22_X1 U22534 ( .A1(n9182), .A2(n24428), .B1(n9183), .B2(n24422), .ZN(
        n23186) );
  OAI22_X1 U22535 ( .A1(n19675), .A2(n24404), .B1(n8925), .B2(n24398), .ZN(
        n23169) );
  OAI22_X1 U22536 ( .A1(n9180), .A2(n24428), .B1(n9181), .B2(n24422), .ZN(
        n23168) );
  OAI22_X1 U22537 ( .A1(n19674), .A2(n24404), .B1(n8923), .B2(n24398), .ZN(
        n23151) );
  OAI22_X1 U22538 ( .A1(n9178), .A2(n24428), .B1(n9179), .B2(n24422), .ZN(
        n23150) );
  OAI22_X1 U22539 ( .A1(n19673), .A2(n24404), .B1(n8921), .B2(n24398), .ZN(
        n23133) );
  OAI22_X1 U22540 ( .A1(n9176), .A2(n24428), .B1(n9177), .B2(n24422), .ZN(
        n23132) );
  OAI22_X1 U22541 ( .A1(n19672), .A2(n24404), .B1(n8919), .B2(n24398), .ZN(
        n23115) );
  OAI22_X1 U22542 ( .A1(n9174), .A2(n24428), .B1(n9175), .B2(n24422), .ZN(
        n23114) );
  OAI22_X1 U22543 ( .A1(n19671), .A2(n24405), .B1(n8917), .B2(n24399), .ZN(
        n23097) );
  OAI22_X1 U22544 ( .A1(n9172), .A2(n24429), .B1(n9173), .B2(n24423), .ZN(
        n23096) );
  OAI22_X1 U22545 ( .A1(n19670), .A2(n24405), .B1(n8915), .B2(n24399), .ZN(
        n23079) );
  OAI22_X1 U22546 ( .A1(n9170), .A2(n24429), .B1(n9171), .B2(n24423), .ZN(
        n23078) );
  OAI22_X1 U22547 ( .A1(n19669), .A2(n24405), .B1(n8913), .B2(n24399), .ZN(
        n23061) );
  OAI22_X1 U22548 ( .A1(n9168), .A2(n24429), .B1(n9169), .B2(n24423), .ZN(
        n23060) );
  OAI22_X1 U22549 ( .A1(n19668), .A2(n24405), .B1(n8911), .B2(n24399), .ZN(
        n23043) );
  OAI22_X1 U22550 ( .A1(n9166), .A2(n24429), .B1(n9167), .B2(n24423), .ZN(
        n23042) );
  OAI22_X1 U22551 ( .A1(n88), .A2(n24495), .B1(n20710), .B2(n24489), .ZN(
        n23023) );
  OAI22_X1 U22552 ( .A1(n87), .A2(n24495), .B1(n20709), .B2(n24489), .ZN(
        n23005) );
  OAI22_X1 U22553 ( .A1(n86), .A2(n24495), .B1(n20708), .B2(n24489), .ZN(
        n22987) );
  OAI22_X1 U22554 ( .A1(n85), .A2(n24495), .B1(n20707), .B2(n24489), .ZN(
        n22969) );
  OAI22_X1 U22555 ( .A1(n84), .A2(n24495), .B1(n20706), .B2(n24489), .ZN(
        n22951) );
  OAI22_X1 U22556 ( .A1(n83), .A2(n24495), .B1(n20705), .B2(n24489), .ZN(
        n22933) );
  OAI22_X1 U22557 ( .A1(n82), .A2(n24495), .B1(n20704), .B2(n24489), .ZN(
        n22915) );
  OAI22_X1 U22558 ( .A1(n81), .A2(n24495), .B1(n20703), .B2(n24489), .ZN(
        n22897) );
  OAI22_X1 U22559 ( .A1(n80), .A2(n24496), .B1(n20702), .B2(n24490), .ZN(
        n22879) );
  OAI22_X1 U22560 ( .A1(n79), .A2(n24496), .B1(n20701), .B2(n24490), .ZN(
        n22861) );
  OAI22_X1 U22561 ( .A1(n78), .A2(n24496), .B1(n20700), .B2(n24490), .ZN(
        n22843) );
  OAI22_X1 U22562 ( .A1(n77), .A2(n24496), .B1(n20699), .B2(n24490), .ZN(
        n22825) );
  OAI22_X1 U22563 ( .A1(n99), .A2(n24494), .B1(n20721), .B2(n24488), .ZN(
        n23221) );
  OAI22_X1 U22564 ( .A1(n98), .A2(n24494), .B1(n20720), .B2(n24488), .ZN(
        n23203) );
  OAI22_X1 U22565 ( .A1(n97), .A2(n24494), .B1(n20719), .B2(n24488), .ZN(
        n23185) );
  OAI22_X1 U22566 ( .A1(n96), .A2(n24494), .B1(n20718), .B2(n24488), .ZN(
        n23167) );
  OAI22_X1 U22567 ( .A1(n95), .A2(n24494), .B1(n20717), .B2(n24488), .ZN(
        n23149) );
  OAI22_X1 U22568 ( .A1(n94), .A2(n24494), .B1(n20716), .B2(n24488), .ZN(
        n23131) );
  OAI22_X1 U22569 ( .A1(n93), .A2(n24494), .B1(n20715), .B2(n24488), .ZN(
        n23113) );
  OAI22_X1 U22570 ( .A1(n92), .A2(n24495), .B1(n20714), .B2(n24489), .ZN(
        n23095) );
  OAI22_X1 U22571 ( .A1(n91), .A2(n24495), .B1(n20713), .B2(n24489), .ZN(
        n23077) );
  OAI22_X1 U22572 ( .A1(n90), .A2(n24495), .B1(n20712), .B2(n24489), .ZN(
        n23059) );
  OAI22_X1 U22573 ( .A1(n89), .A2(n24495), .B1(n20711), .B2(n24489), .ZN(
        n23041) );
  AOI221_X1 U22574 ( .B1(n24666), .B2(n24272), .C1(n24660), .C2(n24148), .A(
        n22555), .ZN(n22550) );
  OAI22_X1 U22575 ( .A1(n20421), .A2(n24654), .B1(n21098), .B2(n24648), .ZN(
        n22555) );
  AOI221_X1 U22576 ( .B1(n24642), .B2(n17541), .C1(n24636), .C2(n24212), .A(
        n22556), .ZN(n22549) );
  OAI22_X1 U22577 ( .A1(n20846), .A2(n24630), .B1(n21122), .B2(n24624), .ZN(
        n22556) );
  AOI221_X1 U22578 ( .B1(n24666), .B2(n24273), .C1(n24660), .C2(n24149), .A(
        n22526), .ZN(n22523) );
  OAI22_X1 U22579 ( .A1(n20420), .A2(n24654), .B1(n21097), .B2(n24648), .ZN(
        n22526) );
  AOI221_X1 U22580 ( .B1(n24642), .B2(n17544), .C1(n24636), .C2(n24213), .A(
        n22527), .ZN(n22522) );
  OAI22_X1 U22581 ( .A1(n20845), .A2(n24630), .B1(n21121), .B2(n24624), .ZN(
        n22527) );
  AOI221_X1 U22582 ( .B1(n24666), .B2(n24274), .C1(n24660), .C2(n24150), .A(
        n22507), .ZN(n22504) );
  OAI22_X1 U22583 ( .A1(n20419), .A2(n24654), .B1(n21096), .B2(n24648), .ZN(
        n22507) );
  AOI221_X1 U22584 ( .B1(n24642), .B2(n17547), .C1(n24636), .C2(n24214), .A(
        n22508), .ZN(n22503) );
  OAI22_X1 U22585 ( .A1(n20844), .A2(n24630), .B1(n21120), .B2(n24624), .ZN(
        n22508) );
  AOI221_X1 U22586 ( .B1(n24666), .B2(n24275), .C1(n24660), .C2(n24151), .A(
        n22488), .ZN(n22485) );
  OAI22_X1 U22587 ( .A1(n20418), .A2(n24654), .B1(n21095), .B2(n24648), .ZN(
        n22488) );
  AOI221_X1 U22588 ( .B1(n24642), .B2(n17550), .C1(n24636), .C2(n24215), .A(
        n22489), .ZN(n22484) );
  OAI22_X1 U22589 ( .A1(n20843), .A2(n24630), .B1(n21119), .B2(n24624), .ZN(
        n22489) );
  AOI221_X1 U22590 ( .B1(n24666), .B2(n24276), .C1(n24660), .C2(n24152), .A(
        n22469), .ZN(n22466) );
  OAI22_X1 U22591 ( .A1(n20417), .A2(n24654), .B1(n21094), .B2(n24648), .ZN(
        n22469) );
  AOI221_X1 U22592 ( .B1(n24642), .B2(n17553), .C1(n24636), .C2(n24216), .A(
        n22470), .ZN(n22465) );
  OAI22_X1 U22593 ( .A1(n20842), .A2(n24630), .B1(n21118), .B2(n24624), .ZN(
        n22470) );
  AOI221_X1 U22594 ( .B1(n24666), .B2(n24277), .C1(n24660), .C2(n24153), .A(
        n22450), .ZN(n22447) );
  OAI22_X1 U22595 ( .A1(n20416), .A2(n24654), .B1(n21093), .B2(n24648), .ZN(
        n22450) );
  AOI221_X1 U22596 ( .B1(n24642), .B2(n17556), .C1(n24636), .C2(n24217), .A(
        n22451), .ZN(n22446) );
  OAI22_X1 U22597 ( .A1(n20841), .A2(n24630), .B1(n21117), .B2(n24624), .ZN(
        n22451) );
  AOI221_X1 U22598 ( .B1(n24666), .B2(n24278), .C1(n24660), .C2(n24154), .A(
        n22431), .ZN(n22428) );
  OAI22_X1 U22599 ( .A1(n20415), .A2(n24654), .B1(n21092), .B2(n24648), .ZN(
        n22431) );
  AOI221_X1 U22600 ( .B1(n24642), .B2(n17559), .C1(n24636), .C2(n24218), .A(
        n22432), .ZN(n22427) );
  OAI22_X1 U22601 ( .A1(n20840), .A2(n24630), .B1(n21116), .B2(n24624), .ZN(
        n22432) );
  AOI221_X1 U22602 ( .B1(n24666), .B2(n24279), .C1(n24660), .C2(n24155), .A(
        n22412), .ZN(n22409) );
  OAI22_X1 U22603 ( .A1(n20414), .A2(n24654), .B1(n21091), .B2(n24648), .ZN(
        n22412) );
  AOI221_X1 U22604 ( .B1(n24642), .B2(n17562), .C1(n24636), .C2(n24219), .A(
        n22413), .ZN(n22408) );
  OAI22_X1 U22605 ( .A1(n20839), .A2(n24630), .B1(n21115), .B2(n24624), .ZN(
        n22413) );
  AOI221_X1 U22606 ( .B1(n24666), .B2(n24280), .C1(n24660), .C2(n24156), .A(
        n22393), .ZN(n22390) );
  OAI22_X1 U22607 ( .A1(n20413), .A2(n24654), .B1(n21090), .B2(n24648), .ZN(
        n22393) );
  AOI221_X1 U22608 ( .B1(n24642), .B2(n17565), .C1(n24636), .C2(n24220), .A(
        n22394), .ZN(n22389) );
  OAI22_X1 U22609 ( .A1(n20838), .A2(n24630), .B1(n21114), .B2(n24624), .ZN(
        n22394) );
  AOI221_X1 U22610 ( .B1(n24666), .B2(n24281), .C1(n24660), .C2(n24157), .A(
        n22374), .ZN(n22371) );
  OAI22_X1 U22611 ( .A1(n20412), .A2(n24654), .B1(n21089), .B2(n24648), .ZN(
        n22374) );
  AOI221_X1 U22612 ( .B1(n24642), .B2(n17568), .C1(n24636), .C2(n24221), .A(
        n22375), .ZN(n22370) );
  OAI22_X1 U22613 ( .A1(n20837), .A2(n24630), .B1(n21113), .B2(n24624), .ZN(
        n22375) );
  AOI221_X1 U22614 ( .B1(n24666), .B2(n24282), .C1(n24660), .C2(n24158), .A(
        n22355), .ZN(n22352) );
  OAI22_X1 U22615 ( .A1(n20411), .A2(n24654), .B1(n21088), .B2(n24648), .ZN(
        n22355) );
  AOI221_X1 U22616 ( .B1(n24642), .B2(n17571), .C1(n24636), .C2(n24222), .A(
        n22356), .ZN(n22351) );
  OAI22_X1 U22617 ( .A1(n20836), .A2(n24630), .B1(n21112), .B2(n24624), .ZN(
        n22356) );
  AOI221_X1 U22618 ( .B1(n24666), .B2(n24283), .C1(n24660), .C2(n24159), .A(
        n22336), .ZN(n22333) );
  OAI22_X1 U22619 ( .A1(n20410), .A2(n24654), .B1(n21087), .B2(n24648), .ZN(
        n22336) );
  AOI221_X1 U22620 ( .B1(n24642), .B2(n17574), .C1(n24636), .C2(n24223), .A(
        n22337), .ZN(n22332) );
  OAI22_X1 U22621 ( .A1(n20835), .A2(n24630), .B1(n21111), .B2(n24624), .ZN(
        n22337) );
  AOI221_X1 U22622 ( .B1(n24667), .B2(n24284), .C1(n24661), .C2(n24160), .A(
        n22317), .ZN(n22314) );
  OAI22_X1 U22623 ( .A1(n20409), .A2(n24655), .B1(n21086), .B2(n24649), .ZN(
        n22317) );
  AOI221_X1 U22624 ( .B1(n24643), .B2(n17577), .C1(n24637), .C2(n24224), .A(
        n22318), .ZN(n22313) );
  OAI22_X1 U22625 ( .A1(n20834), .A2(n24631), .B1(n21110), .B2(n24625), .ZN(
        n22318) );
  AOI221_X1 U22626 ( .B1(n24667), .B2(n24285), .C1(n24661), .C2(n24161), .A(
        n22298), .ZN(n22295) );
  OAI22_X1 U22627 ( .A1(n20408), .A2(n24655), .B1(n21085), .B2(n24649), .ZN(
        n22298) );
  AOI221_X1 U22628 ( .B1(n24643), .B2(n17580), .C1(n24637), .C2(n24225), .A(
        n22299), .ZN(n22294) );
  OAI22_X1 U22629 ( .A1(n20833), .A2(n24631), .B1(n21109), .B2(n24625), .ZN(
        n22299) );
  AOI221_X1 U22630 ( .B1(n24667), .B2(n24286), .C1(n24661), .C2(n24162), .A(
        n22279), .ZN(n22276) );
  OAI22_X1 U22631 ( .A1(n20407), .A2(n24655), .B1(n21084), .B2(n24649), .ZN(
        n22279) );
  AOI221_X1 U22632 ( .B1(n24643), .B2(n17583), .C1(n24637), .C2(n24226), .A(
        n22280), .ZN(n22275) );
  OAI22_X1 U22633 ( .A1(n20832), .A2(n24631), .B1(n21108), .B2(n24625), .ZN(
        n22280) );
  AOI221_X1 U22634 ( .B1(n24667), .B2(n24287), .C1(n24661), .C2(n24163), .A(
        n22260), .ZN(n22257) );
  OAI22_X1 U22635 ( .A1(n20406), .A2(n24655), .B1(n21083), .B2(n24649), .ZN(
        n22260) );
  AOI221_X1 U22636 ( .B1(n24643), .B2(n17586), .C1(n24637), .C2(n24227), .A(
        n22261), .ZN(n22256) );
  OAI22_X1 U22637 ( .A1(n20831), .A2(n24631), .B1(n21107), .B2(n24625), .ZN(
        n22261) );
  AOI221_X1 U22638 ( .B1(n24667), .B2(n24288), .C1(n24661), .C2(n24164), .A(
        n22241), .ZN(n22238) );
  OAI22_X1 U22639 ( .A1(n20405), .A2(n24655), .B1(n21082), .B2(n24649), .ZN(
        n22241) );
  AOI221_X1 U22640 ( .B1(n24643), .B2(n17589), .C1(n24637), .C2(n24228), .A(
        n22242), .ZN(n22237) );
  OAI22_X1 U22641 ( .A1(n20830), .A2(n24631), .B1(n21106), .B2(n24625), .ZN(
        n22242) );
  AOI221_X1 U22642 ( .B1(n24667), .B2(n24289), .C1(n24661), .C2(n24165), .A(
        n22222), .ZN(n22219) );
  OAI22_X1 U22643 ( .A1(n20404), .A2(n24655), .B1(n21081), .B2(n24649), .ZN(
        n22222) );
  AOI221_X1 U22644 ( .B1(n24643), .B2(n17592), .C1(n24637), .C2(n24229), .A(
        n22223), .ZN(n22218) );
  OAI22_X1 U22645 ( .A1(n20829), .A2(n24631), .B1(n21105), .B2(n24625), .ZN(
        n22223) );
  AOI221_X1 U22646 ( .B1(n24667), .B2(n24290), .C1(n24661), .C2(n24166), .A(
        n22203), .ZN(n22200) );
  OAI22_X1 U22647 ( .A1(n20403), .A2(n24655), .B1(n21080), .B2(n24649), .ZN(
        n22203) );
  AOI221_X1 U22648 ( .B1(n24643), .B2(n17595), .C1(n24637), .C2(n24230), .A(
        n22204), .ZN(n22199) );
  OAI22_X1 U22649 ( .A1(n20828), .A2(n24631), .B1(n21104), .B2(n24625), .ZN(
        n22204) );
  AOI221_X1 U22650 ( .B1(n24667), .B2(n24291), .C1(n24661), .C2(n24167), .A(
        n22184), .ZN(n22181) );
  OAI22_X1 U22651 ( .A1(n20402), .A2(n24655), .B1(n21079), .B2(n24649), .ZN(
        n22184) );
  AOI221_X1 U22652 ( .B1(n24643), .B2(n17598), .C1(n24637), .C2(n24231), .A(
        n22185), .ZN(n22180) );
  OAI22_X1 U22653 ( .A1(n20827), .A2(n24631), .B1(n21103), .B2(n24625), .ZN(
        n22185) );
  AOI221_X1 U22654 ( .B1(n24667), .B2(n24292), .C1(n24661), .C2(n24168), .A(
        n22165), .ZN(n22162) );
  OAI22_X1 U22655 ( .A1(n20401), .A2(n24655), .B1(n21078), .B2(n24649), .ZN(
        n22165) );
  AOI221_X1 U22656 ( .B1(n24643), .B2(n17601), .C1(n24637), .C2(n24232), .A(
        n22166), .ZN(n22161) );
  OAI22_X1 U22657 ( .A1(n20826), .A2(n24631), .B1(n21102), .B2(n24625), .ZN(
        n22166) );
  AOI221_X1 U22658 ( .B1(n24667), .B2(n24293), .C1(n24661), .C2(n24169), .A(
        n22146), .ZN(n22143) );
  OAI22_X1 U22659 ( .A1(n20400), .A2(n24655), .B1(n21077), .B2(n24649), .ZN(
        n22146) );
  AOI221_X1 U22660 ( .B1(n24643), .B2(n17604), .C1(n24637), .C2(n24233), .A(
        n22147), .ZN(n22142) );
  OAI22_X1 U22661 ( .A1(n20825), .A2(n24631), .B1(n21101), .B2(n24625), .ZN(
        n22147) );
  AOI221_X1 U22662 ( .B1(n24667), .B2(n24294), .C1(n24661), .C2(n24170), .A(
        n22127), .ZN(n22124) );
  OAI22_X1 U22663 ( .A1(n20399), .A2(n24655), .B1(n21076), .B2(n24649), .ZN(
        n22127) );
  AOI221_X1 U22664 ( .B1(n24643), .B2(n17607), .C1(n24637), .C2(n24234), .A(
        n22128), .ZN(n22123) );
  OAI22_X1 U22665 ( .A1(n20824), .A2(n24631), .B1(n21100), .B2(n24625), .ZN(
        n22128) );
  AOI221_X1 U22666 ( .B1(n24667), .B2(n24295), .C1(n24661), .C2(n24171), .A(
        n22108), .ZN(n22105) );
  OAI22_X1 U22667 ( .A1(n20398), .A2(n24655), .B1(n21075), .B2(n24649), .ZN(
        n22108) );
  AOI221_X1 U22668 ( .B1(n24643), .B2(n17610), .C1(n24637), .C2(n24235), .A(
        n22109), .ZN(n22104) );
  OAI22_X1 U22669 ( .A1(n20823), .A2(n24631), .B1(n21099), .B2(n24625), .ZN(
        n22109) );
  AOI221_X1 U22670 ( .B1(n24668), .B2(n24296), .C1(n24662), .C2(n24172), .A(
        n22089), .ZN(n22086) );
  OAI22_X1 U22671 ( .A1(n20337), .A2(n24656), .B1(n20978), .B2(n24650), .ZN(
        n22089) );
  AOI221_X1 U22672 ( .B1(n24644), .B2(n17613), .C1(n24638), .C2(n24236), .A(
        n22090), .ZN(n22085) );
  OAI22_X1 U22673 ( .A1(n20726), .A2(n24632), .B1(n21014), .B2(n24626), .ZN(
        n22090) );
  AOI221_X1 U22674 ( .B1(n24668), .B2(n24297), .C1(n24662), .C2(n24173), .A(
        n22070), .ZN(n22067) );
  OAI22_X1 U22675 ( .A1(n20336), .A2(n24656), .B1(n20977), .B2(n24650), .ZN(
        n22070) );
  AOI221_X1 U22676 ( .B1(n24644), .B2(n17616), .C1(n24638), .C2(n24237), .A(
        n22071), .ZN(n22066) );
  OAI22_X1 U22677 ( .A1(n20725), .A2(n24632), .B1(n21013), .B2(n24626), .ZN(
        n22071) );
  AOI221_X1 U22678 ( .B1(n24668), .B2(n24298), .C1(n24662), .C2(n24174), .A(
        n22051), .ZN(n22048) );
  OAI22_X1 U22679 ( .A1(n20335), .A2(n24656), .B1(n20976), .B2(n24650), .ZN(
        n22051) );
  AOI221_X1 U22680 ( .B1(n24644), .B2(n17619), .C1(n24638), .C2(n24238), .A(
        n22052), .ZN(n22047) );
  OAI22_X1 U22681 ( .A1(n20724), .A2(n24632), .B1(n21012), .B2(n24626), .ZN(
        n22052) );
  AOI221_X1 U22682 ( .B1(n24668), .B2(n24299), .C1(n24662), .C2(n24175), .A(
        n22032), .ZN(n22029) );
  OAI22_X1 U22683 ( .A1(n20334), .A2(n24656), .B1(n20975), .B2(n24650), .ZN(
        n22032) );
  AOI221_X1 U22684 ( .B1(n24644), .B2(n17622), .C1(n24638), .C2(n24239), .A(
        n22033), .ZN(n22028) );
  OAI22_X1 U22685 ( .A1(n20723), .A2(n24632), .B1(n21011), .B2(n24626), .ZN(
        n22033) );
  AOI221_X1 U22686 ( .B1(n24668), .B2(n24300), .C1(n24662), .C2(n24176), .A(
        n22013), .ZN(n22010) );
  OAI22_X1 U22687 ( .A1(n20333), .A2(n24656), .B1(n20974), .B2(n24650), .ZN(
        n22013) );
  AOI221_X1 U22688 ( .B1(n24644), .B2(n17625), .C1(n24638), .C2(n24240), .A(
        n22014), .ZN(n22009) );
  OAI22_X1 U22689 ( .A1(n20722), .A2(n24632), .B1(n21010), .B2(n24626), .ZN(
        n22014) );
  AOI221_X1 U22690 ( .B1(n24668), .B2(n24301), .C1(n24662), .C2(n24177), .A(
        n21994), .ZN(n21991) );
  OAI22_X1 U22691 ( .A1(n20332), .A2(n24656), .B1(n20973), .B2(n24650), .ZN(
        n21994) );
  AOI221_X1 U22692 ( .B1(n24644), .B2(n17472), .C1(n24638), .C2(n24241), .A(
        n21995), .ZN(n21990) );
  OAI22_X1 U22693 ( .A1(n20721), .A2(n24632), .B1(n21009), .B2(n24626), .ZN(
        n21995) );
  AOI221_X1 U22694 ( .B1(n24668), .B2(n24302), .C1(n24662), .C2(n24178), .A(
        n21975), .ZN(n21972) );
  OAI22_X1 U22695 ( .A1(n20331), .A2(n24656), .B1(n20972), .B2(n24650), .ZN(
        n21975) );
  AOI221_X1 U22696 ( .B1(n24644), .B2(n17475), .C1(n24638), .C2(n24242), .A(
        n21976), .ZN(n21971) );
  OAI22_X1 U22697 ( .A1(n20720), .A2(n24632), .B1(n21008), .B2(n24626), .ZN(
        n21976) );
  AOI221_X1 U22698 ( .B1(n24668), .B2(n24303), .C1(n24662), .C2(n24179), .A(
        n21956), .ZN(n21953) );
  OAI22_X1 U22699 ( .A1(n20330), .A2(n24656), .B1(n20971), .B2(n24650), .ZN(
        n21956) );
  AOI221_X1 U22700 ( .B1(n24644), .B2(n17478), .C1(n24638), .C2(n24243), .A(
        n21957), .ZN(n21952) );
  OAI22_X1 U22701 ( .A1(n20719), .A2(n24632), .B1(n21007), .B2(n24626), .ZN(
        n21957) );
  AOI221_X1 U22702 ( .B1(n24668), .B2(n24304), .C1(n24662), .C2(n24180), .A(
        n21937), .ZN(n21934) );
  OAI22_X1 U22703 ( .A1(n20329), .A2(n24656), .B1(n20970), .B2(n24650), .ZN(
        n21937) );
  AOI221_X1 U22704 ( .B1(n24644), .B2(n17481), .C1(n24638), .C2(n24244), .A(
        n21938), .ZN(n21933) );
  OAI22_X1 U22705 ( .A1(n20718), .A2(n24632), .B1(n21006), .B2(n24626), .ZN(
        n21938) );
  AOI221_X1 U22706 ( .B1(n24668), .B2(n24305), .C1(n24662), .C2(n24181), .A(
        n21918), .ZN(n21915) );
  OAI22_X1 U22707 ( .A1(n20328), .A2(n24656), .B1(n20969), .B2(n24650), .ZN(
        n21918) );
  AOI221_X1 U22708 ( .B1(n24644), .B2(n17484), .C1(n24638), .C2(n24245), .A(
        n21919), .ZN(n21914) );
  OAI22_X1 U22709 ( .A1(n20717), .A2(n24632), .B1(n21005), .B2(n24626), .ZN(
        n21919) );
  AOI221_X1 U22710 ( .B1(n24668), .B2(n24306), .C1(n24662), .C2(n24182), .A(
        n21899), .ZN(n21896) );
  OAI22_X1 U22711 ( .A1(n20327), .A2(n24656), .B1(n20968), .B2(n24650), .ZN(
        n21899) );
  AOI221_X1 U22712 ( .B1(n24644), .B2(n17487), .C1(n24638), .C2(n24246), .A(
        n21900), .ZN(n21895) );
  OAI22_X1 U22713 ( .A1(n20716), .A2(n24632), .B1(n21004), .B2(n24626), .ZN(
        n21900) );
  AOI221_X1 U22714 ( .B1(n24668), .B2(n24307), .C1(n24662), .C2(n24183), .A(
        n21880), .ZN(n21877) );
  OAI22_X1 U22715 ( .A1(n20326), .A2(n24656), .B1(n20967), .B2(n24650), .ZN(
        n21880) );
  AOI221_X1 U22716 ( .B1(n24644), .B2(n17490), .C1(n24638), .C2(n24247), .A(
        n21881), .ZN(n21876) );
  OAI22_X1 U22717 ( .A1(n20715), .A2(n24632), .B1(n21003), .B2(n24626), .ZN(
        n21881) );
  AOI221_X1 U22718 ( .B1(n24669), .B2(n24308), .C1(n24663), .C2(n24184), .A(
        n21861), .ZN(n21858) );
  OAI22_X1 U22719 ( .A1(n20325), .A2(n24657), .B1(n20966), .B2(n24651), .ZN(
        n21861) );
  AOI221_X1 U22720 ( .B1(n24645), .B2(n17493), .C1(n24639), .C2(n24248), .A(
        n21862), .ZN(n21857) );
  OAI22_X1 U22721 ( .A1(n20714), .A2(n24633), .B1(n21002), .B2(n24627), .ZN(
        n21862) );
  AOI221_X1 U22722 ( .B1(n24669), .B2(n24309), .C1(n24663), .C2(n24185), .A(
        n21842), .ZN(n21839) );
  OAI22_X1 U22723 ( .A1(n20324), .A2(n24657), .B1(n20965), .B2(n24651), .ZN(
        n21842) );
  AOI221_X1 U22724 ( .B1(n24645), .B2(n17496), .C1(n24639), .C2(n24249), .A(
        n21843), .ZN(n21838) );
  OAI22_X1 U22725 ( .A1(n20713), .A2(n24633), .B1(n21001), .B2(n24627), .ZN(
        n21843) );
  AOI221_X1 U22726 ( .B1(n24669), .B2(n24310), .C1(n24663), .C2(n24186), .A(
        n21823), .ZN(n21820) );
  OAI22_X1 U22727 ( .A1(n20323), .A2(n24657), .B1(n20964), .B2(n24651), .ZN(
        n21823) );
  AOI221_X1 U22728 ( .B1(n24645), .B2(n17499), .C1(n24639), .C2(n24250), .A(
        n21824), .ZN(n21819) );
  OAI22_X1 U22729 ( .A1(n20712), .A2(n24633), .B1(n21000), .B2(n24627), .ZN(
        n21824) );
  AOI221_X1 U22730 ( .B1(n24669), .B2(n24311), .C1(n24663), .C2(n24187), .A(
        n21804), .ZN(n21801) );
  OAI22_X1 U22731 ( .A1(n20322), .A2(n24657), .B1(n20963), .B2(n24651), .ZN(
        n21804) );
  AOI221_X1 U22732 ( .B1(n24645), .B2(n17502), .C1(n24639), .C2(n24251), .A(
        n21805), .ZN(n21800) );
  OAI22_X1 U22733 ( .A1(n20711), .A2(n24633), .B1(n20999), .B2(n24627), .ZN(
        n21805) );
  AOI221_X1 U22734 ( .B1(n24669), .B2(n24312), .C1(n24663), .C2(n24188), .A(
        n21785), .ZN(n21782) );
  OAI22_X1 U22735 ( .A1(n20321), .A2(n24657), .B1(n20962), .B2(n24651), .ZN(
        n21785) );
  AOI221_X1 U22736 ( .B1(n24645), .B2(n17505), .C1(n24639), .C2(n24252), .A(
        n21786), .ZN(n21781) );
  OAI22_X1 U22737 ( .A1(n20710), .A2(n24633), .B1(n20998), .B2(n24627), .ZN(
        n21786) );
  AOI221_X1 U22738 ( .B1(n24669), .B2(n24313), .C1(n24663), .C2(n24189), .A(
        n21766), .ZN(n21763) );
  OAI22_X1 U22739 ( .A1(n20320), .A2(n24657), .B1(n20961), .B2(n24651), .ZN(
        n21766) );
  AOI221_X1 U22740 ( .B1(n24645), .B2(n17508), .C1(n24639), .C2(n24253), .A(
        n21767), .ZN(n21762) );
  OAI22_X1 U22741 ( .A1(n20709), .A2(n24633), .B1(n20997), .B2(n24627), .ZN(
        n21767) );
  AOI221_X1 U22742 ( .B1(n24669), .B2(n24314), .C1(n24663), .C2(n24190), .A(
        n21747), .ZN(n21744) );
  OAI22_X1 U22743 ( .A1(n20319), .A2(n24657), .B1(n20960), .B2(n24651), .ZN(
        n21747) );
  AOI221_X1 U22744 ( .B1(n24645), .B2(n17511), .C1(n24639), .C2(n24254), .A(
        n21748), .ZN(n21743) );
  OAI22_X1 U22745 ( .A1(n20708), .A2(n24633), .B1(n20996), .B2(n24627), .ZN(
        n21748) );
  AOI221_X1 U22746 ( .B1(n24669), .B2(n24315), .C1(n24663), .C2(n24191), .A(
        n21728), .ZN(n21725) );
  OAI22_X1 U22747 ( .A1(n20318), .A2(n24657), .B1(n20959), .B2(n24651), .ZN(
        n21728) );
  AOI221_X1 U22748 ( .B1(n24645), .B2(n17514), .C1(n24639), .C2(n24255), .A(
        n21729), .ZN(n21724) );
  OAI22_X1 U22749 ( .A1(n20707), .A2(n24633), .B1(n20995), .B2(n24627), .ZN(
        n21729) );
  AOI221_X1 U22750 ( .B1(n24669), .B2(n24316), .C1(n24663), .C2(n24192), .A(
        n21709), .ZN(n21706) );
  OAI22_X1 U22751 ( .A1(n20317), .A2(n24657), .B1(n20958), .B2(n24651), .ZN(
        n21709) );
  AOI221_X1 U22752 ( .B1(n24645), .B2(n17517), .C1(n24639), .C2(n24256), .A(
        n21710), .ZN(n21705) );
  OAI22_X1 U22753 ( .A1(n20706), .A2(n24633), .B1(n20994), .B2(n24627), .ZN(
        n21710) );
  AOI221_X1 U22754 ( .B1(n24669), .B2(n24317), .C1(n24663), .C2(n24193), .A(
        n21690), .ZN(n21687) );
  OAI22_X1 U22755 ( .A1(n20316), .A2(n24657), .B1(n20957), .B2(n24651), .ZN(
        n21690) );
  AOI221_X1 U22756 ( .B1(n24645), .B2(n17520), .C1(n24639), .C2(n24257), .A(
        n21691), .ZN(n21686) );
  OAI22_X1 U22757 ( .A1(n20705), .A2(n24633), .B1(n20993), .B2(n24627), .ZN(
        n21691) );
  AOI221_X1 U22758 ( .B1(n24669), .B2(n24318), .C1(n24663), .C2(n24194), .A(
        n21671), .ZN(n21668) );
  OAI22_X1 U22759 ( .A1(n20315), .A2(n24657), .B1(n20956), .B2(n24651), .ZN(
        n21671) );
  AOI221_X1 U22760 ( .B1(n24645), .B2(n17523), .C1(n24639), .C2(n24258), .A(
        n21672), .ZN(n21667) );
  OAI22_X1 U22761 ( .A1(n20704), .A2(n24633), .B1(n20992), .B2(n24627), .ZN(
        n21672) );
  AOI221_X1 U22762 ( .B1(n24669), .B2(n24319), .C1(n24663), .C2(n24195), .A(
        n21652), .ZN(n21649) );
  OAI22_X1 U22763 ( .A1(n20314), .A2(n24657), .B1(n20955), .B2(n24651), .ZN(
        n21652) );
  AOI221_X1 U22764 ( .B1(n24645), .B2(n17526), .C1(n24639), .C2(n24259), .A(
        n21653), .ZN(n21648) );
  OAI22_X1 U22765 ( .A1(n20703), .A2(n24633), .B1(n20991), .B2(n24627), .ZN(
        n21653) );
  AOI221_X1 U22766 ( .B1(n24670), .B2(n24320), .C1(n24664), .C2(n24196), .A(
        n21633), .ZN(n21630) );
  OAI22_X1 U22767 ( .A1(n20313), .A2(n24658), .B1(n20954), .B2(n24652), .ZN(
        n21633) );
  AOI221_X1 U22768 ( .B1(n24646), .B2(n17529), .C1(n24640), .C2(n24260), .A(
        n21634), .ZN(n21629) );
  OAI22_X1 U22769 ( .A1(n20702), .A2(n24634), .B1(n20990), .B2(n24628), .ZN(
        n21634) );
  AOI221_X1 U22770 ( .B1(n24670), .B2(n24321), .C1(n24664), .C2(n24197), .A(
        n21614), .ZN(n21611) );
  OAI22_X1 U22771 ( .A1(n20312), .A2(n24658), .B1(n20953), .B2(n24652), .ZN(
        n21614) );
  AOI221_X1 U22772 ( .B1(n24646), .B2(n17532), .C1(n24640), .C2(n24261), .A(
        n21615), .ZN(n21610) );
  OAI22_X1 U22773 ( .A1(n20701), .A2(n24634), .B1(n20989), .B2(n24628), .ZN(
        n21615) );
  AOI221_X1 U22774 ( .B1(n24670), .B2(n24322), .C1(n24664), .C2(n24198), .A(
        n21595), .ZN(n21592) );
  OAI22_X1 U22775 ( .A1(n20311), .A2(n24658), .B1(n20952), .B2(n24652), .ZN(
        n21595) );
  AOI221_X1 U22776 ( .B1(n24646), .B2(n17535), .C1(n24640), .C2(n24262), .A(
        n21596), .ZN(n21591) );
  OAI22_X1 U22777 ( .A1(n20700), .A2(n24634), .B1(n20988), .B2(n24628), .ZN(
        n21596) );
  AOI221_X1 U22778 ( .B1(n24670), .B2(n24323), .C1(n24664), .C2(n24199), .A(
        n21576), .ZN(n21573) );
  OAI22_X1 U22779 ( .A1(n20310), .A2(n24658), .B1(n20951), .B2(n24652), .ZN(
        n21576) );
  AOI221_X1 U22780 ( .B1(n24646), .B2(n17538), .C1(n24640), .C2(n24263), .A(
        n21577), .ZN(n21572) );
  OAI22_X1 U22781 ( .A1(n20699), .A2(n24634), .B1(n20987), .B2(n24628), .ZN(
        n21577) );
  AOI221_X1 U22782 ( .B1(n24670), .B2(n24324), .C1(n24664), .C2(n24200), .A(
        n21557), .ZN(n21554) );
  OAI22_X1 U22783 ( .A1(n20309), .A2(n24658), .B1(n20950), .B2(n24652), .ZN(
        n21557) );
  AOI221_X1 U22784 ( .B1(n24646), .B2(n17628), .C1(n24640), .C2(n24264), .A(
        n21558), .ZN(n21553) );
  OAI22_X1 U22785 ( .A1(n20698), .A2(n24634), .B1(n20986), .B2(n24628), .ZN(
        n21558) );
  AOI221_X1 U22786 ( .B1(n24670), .B2(n24325), .C1(n24664), .C2(n24201), .A(
        n21538), .ZN(n21535) );
  OAI22_X1 U22787 ( .A1(n20308), .A2(n24658), .B1(n20949), .B2(n24652), .ZN(
        n21538) );
  AOI221_X1 U22788 ( .B1(n24646), .B2(n17631), .C1(n24640), .C2(n24265), .A(
        n21539), .ZN(n21534) );
  OAI22_X1 U22789 ( .A1(n20697), .A2(n24634), .B1(n20985), .B2(n24628), .ZN(
        n21539) );
  AOI221_X1 U22790 ( .B1(n24670), .B2(n24326), .C1(n24664), .C2(n24202), .A(
        n21519), .ZN(n21516) );
  OAI22_X1 U22791 ( .A1(n20307), .A2(n24658), .B1(n20948), .B2(n24652), .ZN(
        n21519) );
  AOI221_X1 U22792 ( .B1(n24646), .B2(n17634), .C1(n24640), .C2(n24266), .A(
        n21520), .ZN(n21515) );
  OAI22_X1 U22793 ( .A1(n20696), .A2(n24634), .B1(n20984), .B2(n24628), .ZN(
        n21520) );
  AOI221_X1 U22794 ( .B1(n24670), .B2(n24327), .C1(n24664), .C2(n24203), .A(
        n21500), .ZN(n21497) );
  OAI22_X1 U22795 ( .A1(n20306), .A2(n24658), .B1(n20947), .B2(n24652), .ZN(
        n21500) );
  AOI221_X1 U22796 ( .B1(n24646), .B2(n17637), .C1(n24640), .C2(n24267), .A(
        n21501), .ZN(n21496) );
  OAI22_X1 U22797 ( .A1(n20695), .A2(n24634), .B1(n20983), .B2(n24628), .ZN(
        n21501) );
  AOI221_X1 U22798 ( .B1(n24670), .B2(n24328), .C1(n24664), .C2(n24204), .A(
        n21481), .ZN(n21478) );
  OAI22_X1 U22799 ( .A1(n20305), .A2(n24658), .B1(n20946), .B2(n24652), .ZN(
        n21481) );
  AOI221_X1 U22800 ( .B1(n24646), .B2(n17640), .C1(n24640), .C2(n24268), .A(
        n21482), .ZN(n21477) );
  OAI22_X1 U22801 ( .A1(n20694), .A2(n24634), .B1(n20982), .B2(n24628), .ZN(
        n21482) );
  AOI221_X1 U22802 ( .B1(n24670), .B2(n24329), .C1(n24664), .C2(n24205), .A(
        n21462), .ZN(n21459) );
  OAI22_X1 U22803 ( .A1(n20304), .A2(n24658), .B1(n20945), .B2(n24652), .ZN(
        n21462) );
  AOI221_X1 U22804 ( .B1(n24646), .B2(n17643), .C1(n24640), .C2(n24269), .A(
        n21463), .ZN(n21458) );
  OAI22_X1 U22805 ( .A1(n20693), .A2(n24634), .B1(n20981), .B2(n24628), .ZN(
        n21463) );
  AOI221_X1 U22806 ( .B1(n24670), .B2(n24330), .C1(n24664), .C2(n24206), .A(
        n21443), .ZN(n21440) );
  OAI22_X1 U22807 ( .A1(n20303), .A2(n24658), .B1(n20944), .B2(n24652), .ZN(
        n21443) );
  AOI221_X1 U22808 ( .B1(n24646), .B2(n17646), .C1(n24640), .C2(n24270), .A(
        n21444), .ZN(n21439) );
  OAI22_X1 U22809 ( .A1(n20692), .A2(n24634), .B1(n20980), .B2(n24628), .ZN(
        n21444) );
  AOI221_X1 U22810 ( .B1(n24670), .B2(n24331), .C1(n24664), .C2(n24207), .A(
        n21424), .ZN(n21421) );
  OAI22_X1 U22811 ( .A1(n20302), .A2(n24658), .B1(n20943), .B2(n24652), .ZN(
        n21424) );
  AOI221_X1 U22812 ( .B1(n24646), .B2(n17649), .C1(n24640), .C2(n24271), .A(
        n21425), .ZN(n21420) );
  OAI22_X1 U22813 ( .A1(n20691), .A2(n24634), .B1(n20979), .B2(n24628), .ZN(
        n21425) );
  OAI22_X1 U22814 ( .A1(n24824), .A2(n20213), .B1(n24818), .B2(n25467), .ZN(
        n5100) );
  OAI22_X1 U22815 ( .A1(n24824), .A2(n20212), .B1(n24818), .B2(n25470), .ZN(
        n5101) );
  OAI22_X1 U22816 ( .A1(n24824), .A2(n20211), .B1(n24818), .B2(n25473), .ZN(
        n5102) );
  OAI22_X1 U22817 ( .A1(n24824), .A2(n20210), .B1(n24818), .B2(n25476), .ZN(
        n5103) );
  OAI22_X1 U22818 ( .A1(n24823), .A2(n20209), .B1(n24818), .B2(n25479), .ZN(
        n5104) );
  OAI22_X1 U22819 ( .A1(n24823), .A2(n20208), .B1(n24818), .B2(n25482), .ZN(
        n5105) );
  OAI22_X1 U22820 ( .A1(n24823), .A2(n20207), .B1(n24818), .B2(n25485), .ZN(
        n5106) );
  OAI22_X1 U22821 ( .A1(n24823), .A2(n20206), .B1(n24818), .B2(n25488), .ZN(
        n5107) );
  OAI22_X1 U22822 ( .A1(n24823), .A2(n20205), .B1(n24818), .B2(n25491), .ZN(
        n5108) );
  OAI22_X1 U22823 ( .A1(n24822), .A2(n20204), .B1(n24818), .B2(n25494), .ZN(
        n5109) );
  OAI22_X1 U22824 ( .A1(n24822), .A2(n20203), .B1(n24818), .B2(n25497), .ZN(
        n5110) );
  OAI22_X1 U22825 ( .A1(n24822), .A2(n20202), .B1(n24818), .B2(n25500), .ZN(
        n5111) );
  OAI22_X1 U22826 ( .A1(n24822), .A2(n20201), .B1(n24817), .B2(n25503), .ZN(
        n5112) );
  OAI22_X1 U22827 ( .A1(n24822), .A2(n20200), .B1(n24817), .B2(n25506), .ZN(
        n5113) );
  OAI22_X1 U22828 ( .A1(n24821), .A2(n20199), .B1(n24817), .B2(n25509), .ZN(
        n5114) );
  OAI22_X1 U22829 ( .A1(n24821), .A2(n20198), .B1(n24817), .B2(n25512), .ZN(
        n5115) );
  OAI22_X1 U22830 ( .A1(n24821), .A2(n20197), .B1(n24817), .B2(n25515), .ZN(
        n5116) );
  OAI22_X1 U22831 ( .A1(n24821), .A2(n20196), .B1(n24817), .B2(n25518), .ZN(
        n5117) );
  OAI22_X1 U22832 ( .A1(n24821), .A2(n20195), .B1(n24817), .B2(n25521), .ZN(
        n5118) );
  OAI22_X1 U22833 ( .A1(n24820), .A2(n20194), .B1(n24817), .B2(n25524), .ZN(
        n5119) );
  OAI22_X1 U22834 ( .A1(n24820), .A2(n20193), .B1(n24817), .B2(n25527), .ZN(
        n5120) );
  OAI22_X1 U22835 ( .A1(n24820), .A2(n20192), .B1(n24817), .B2(n25530), .ZN(
        n5121) );
  OAI22_X1 U22836 ( .A1(n24820), .A2(n20191), .B1(n24817), .B2(n25533), .ZN(
        n5122) );
  OAI22_X1 U22837 ( .A1(n24820), .A2(n20190), .B1(n24817), .B2(n25553), .ZN(
        n5123) );
  AOI22_X1 U22838 ( .A1(n24561), .A2(n8053), .B1(n24555), .B2(n8245), .ZN(
        n23017) );
  AOI22_X1 U22839 ( .A1(n24537), .A2(n8309), .B1(n24531), .B2(n23936), .ZN(
        n23018) );
  AOI22_X1 U22840 ( .A1(n24561), .A2(n8052), .B1(n24555), .B2(n8244), .ZN(
        n22999) );
  AOI22_X1 U22841 ( .A1(n24537), .A2(n8308), .B1(n24531), .B2(n23938), .ZN(
        n23000) );
  AOI22_X1 U22842 ( .A1(n24561), .A2(n8051), .B1(n24555), .B2(n8243), .ZN(
        n22981) );
  AOI22_X1 U22843 ( .A1(n24537), .A2(n8307), .B1(n24531), .B2(n23940), .ZN(
        n22982) );
  AOI22_X1 U22844 ( .A1(n24561), .A2(n8050), .B1(n24555), .B2(n8242), .ZN(
        n22963) );
  AOI22_X1 U22845 ( .A1(n24537), .A2(n8306), .B1(n24531), .B2(n23942), .ZN(
        n22964) );
  AOI22_X1 U22846 ( .A1(n24561), .A2(n8049), .B1(n24555), .B2(n8241), .ZN(
        n22945) );
  AOI22_X1 U22847 ( .A1(n24537), .A2(n8305), .B1(n24531), .B2(n23944), .ZN(
        n22946) );
  AOI22_X1 U22848 ( .A1(n24561), .A2(n8048), .B1(n24555), .B2(n8240), .ZN(
        n22927) );
  AOI22_X1 U22849 ( .A1(n24537), .A2(n8304), .B1(n24531), .B2(n23946), .ZN(
        n22928) );
  AOI22_X1 U22850 ( .A1(n24561), .A2(n8047), .B1(n24555), .B2(n8239), .ZN(
        n22909) );
  AOI22_X1 U22851 ( .A1(n24537), .A2(n8303), .B1(n24531), .B2(n23948), .ZN(
        n22910) );
  AOI22_X1 U22852 ( .A1(n24561), .A2(n8046), .B1(n24555), .B2(n8238), .ZN(
        n22891) );
  AOI22_X1 U22853 ( .A1(n24537), .A2(n8302), .B1(n24531), .B2(n23950), .ZN(
        n22892) );
  AOI22_X1 U22854 ( .A1(n24562), .A2(n8045), .B1(n24556), .B2(n8237), .ZN(
        n22873) );
  AOI22_X1 U22855 ( .A1(n24538), .A2(n8301), .B1(n24532), .B2(n23952), .ZN(
        n22874) );
  AOI22_X1 U22856 ( .A1(n24562), .A2(n8044), .B1(n24556), .B2(n8236), .ZN(
        n22855) );
  AOI22_X1 U22857 ( .A1(n24538), .A2(n8300), .B1(n24532), .B2(n23953), .ZN(
        n22856) );
  AOI22_X1 U22858 ( .A1(n24562), .A2(n8043), .B1(n24556), .B2(n8235), .ZN(
        n22837) );
  AOI22_X1 U22859 ( .A1(n24538), .A2(n8299), .B1(n24532), .B2(n23954), .ZN(
        n22838) );
  AOI22_X1 U22860 ( .A1(n24562), .A2(n8042), .B1(n24556), .B2(n8234), .ZN(
        n22819) );
  AOI22_X1 U22861 ( .A1(n24538), .A2(n8298), .B1(n24532), .B2(n23955), .ZN(
        n22820) );
  AOI22_X1 U22862 ( .A1(n24562), .A2(n8041), .B1(n24556), .B2(n8233), .ZN(
        n22801) );
  AOI22_X1 U22863 ( .A1(n24538), .A2(n8297), .B1(n24532), .B2(n23956), .ZN(
        n22802) );
  AOI22_X1 U22864 ( .A1(n24562), .A2(n8040), .B1(n24556), .B2(n8232), .ZN(
        n22783) );
  AOI22_X1 U22865 ( .A1(n24538), .A2(n8296), .B1(n24532), .B2(n23957), .ZN(
        n22784) );
  AOI22_X1 U22866 ( .A1(n24562), .A2(n8039), .B1(n24556), .B2(n8231), .ZN(
        n22765) );
  AOI22_X1 U22867 ( .A1(n24538), .A2(n8295), .B1(n24532), .B2(n23958), .ZN(
        n22766) );
  AOI22_X1 U22868 ( .A1(n24562), .A2(n8038), .B1(n24556), .B2(n8230), .ZN(
        n22747) );
  AOI22_X1 U22869 ( .A1(n24538), .A2(n8294), .B1(n24532), .B2(n23959), .ZN(
        n22748) );
  AOI22_X1 U22870 ( .A1(n24562), .A2(n8037), .B1(n24556), .B2(n8229), .ZN(
        n22729) );
  AOI22_X1 U22871 ( .A1(n24538), .A2(n8293), .B1(n24532), .B2(n23960), .ZN(
        n22730) );
  AOI22_X1 U22872 ( .A1(n24562), .A2(n8036), .B1(n24556), .B2(n8228), .ZN(
        n22711) );
  AOI22_X1 U22873 ( .A1(n24538), .A2(n8292), .B1(n24532), .B2(n23961), .ZN(
        n22712) );
  AOI22_X1 U22874 ( .A1(n24562), .A2(n8035), .B1(n24556), .B2(n8227), .ZN(
        n22693) );
  AOI22_X1 U22875 ( .A1(n24538), .A2(n8291), .B1(n24532), .B2(n23962), .ZN(
        n22694) );
  AOI22_X1 U22876 ( .A1(n24562), .A2(n8034), .B1(n24556), .B2(n8226), .ZN(
        n22675) );
  AOI22_X1 U22877 ( .A1(n24538), .A2(n8290), .B1(n24532), .B2(n23963), .ZN(
        n22676) );
  AOI22_X1 U22878 ( .A1(n24563), .A2(n8033), .B1(n24557), .B2(n8225), .ZN(
        n22657) );
  AOI22_X1 U22879 ( .A1(n24539), .A2(n8289), .B1(n24533), .B2(n23964), .ZN(
        n22658) );
  AOI22_X1 U22880 ( .A1(n24563), .A2(n8032), .B1(n24557), .B2(n8224), .ZN(
        n22639) );
  AOI22_X1 U22881 ( .A1(n24539), .A2(n8288), .B1(n24533), .B2(n23965), .ZN(
        n22640) );
  AOI22_X1 U22882 ( .A1(n24563), .A2(n8031), .B1(n24557), .B2(n8223), .ZN(
        n22621) );
  AOI22_X1 U22883 ( .A1(n24539), .A2(n8287), .B1(n24533), .B2(n23966), .ZN(
        n22622) );
  AOI22_X1 U22884 ( .A1(n24563), .A2(n8030), .B1(n24557), .B2(n8222), .ZN(
        n22575) );
  AOI22_X1 U22885 ( .A1(n24539), .A2(n8286), .B1(n24533), .B2(n23967), .ZN(
        n22580) );
  AOI22_X1 U22886 ( .A1(n24558), .A2(n8093), .B1(n24552), .B2(n8285), .ZN(
        n23743) );
  AOI22_X1 U22887 ( .A1(n24534), .A2(n8349), .B1(n24528), .B2(n23856), .ZN(
        n23746) );
  AOI22_X1 U22888 ( .A1(n24558), .A2(n8092), .B1(n24552), .B2(n8284), .ZN(
        n23719) );
  AOI22_X1 U22889 ( .A1(n24534), .A2(n8348), .B1(n24528), .B2(n23858), .ZN(
        n23720) );
  AOI22_X1 U22890 ( .A1(n24558), .A2(n8091), .B1(n24552), .B2(n8283), .ZN(
        n23701) );
  AOI22_X1 U22891 ( .A1(n24534), .A2(n8347), .B1(n24528), .B2(n23860), .ZN(
        n23702) );
  AOI22_X1 U22892 ( .A1(n24558), .A2(n8090), .B1(n24552), .B2(n8282), .ZN(
        n23683) );
  AOI22_X1 U22893 ( .A1(n24534), .A2(n8346), .B1(n24528), .B2(n23862), .ZN(
        n23684) );
  AOI22_X1 U22894 ( .A1(n24558), .A2(n8089), .B1(n24552), .B2(n8281), .ZN(
        n23665) );
  AOI22_X1 U22895 ( .A1(n24534), .A2(n8345), .B1(n24528), .B2(n23864), .ZN(
        n23666) );
  AOI22_X1 U22896 ( .A1(n24558), .A2(n8088), .B1(n24552), .B2(n8280), .ZN(
        n23647) );
  AOI22_X1 U22897 ( .A1(n24534), .A2(n8344), .B1(n24528), .B2(n23866), .ZN(
        n23648) );
  AOI22_X1 U22898 ( .A1(n24558), .A2(n8087), .B1(n24552), .B2(n8279), .ZN(
        n23629) );
  AOI22_X1 U22899 ( .A1(n24534), .A2(n8343), .B1(n24528), .B2(n23868), .ZN(
        n23630) );
  AOI22_X1 U22900 ( .A1(n24558), .A2(n8086), .B1(n24552), .B2(n8278), .ZN(
        n23611) );
  AOI22_X1 U22901 ( .A1(n24534), .A2(n8342), .B1(n24528), .B2(n23870), .ZN(
        n23612) );
  AOI22_X1 U22902 ( .A1(n24558), .A2(n8085), .B1(n24552), .B2(n8277), .ZN(
        n23593) );
  AOI22_X1 U22903 ( .A1(n24534), .A2(n8341), .B1(n24528), .B2(n23872), .ZN(
        n23594) );
  AOI22_X1 U22904 ( .A1(n24558), .A2(n8084), .B1(n24552), .B2(n8276), .ZN(
        n23575) );
  AOI22_X1 U22905 ( .A1(n24534), .A2(n8340), .B1(n24528), .B2(n23874), .ZN(
        n23576) );
  AOI22_X1 U22906 ( .A1(n24558), .A2(n8083), .B1(n24552), .B2(n8275), .ZN(
        n23557) );
  AOI22_X1 U22907 ( .A1(n24534), .A2(n8339), .B1(n24528), .B2(n23876), .ZN(
        n23558) );
  AOI22_X1 U22908 ( .A1(n24558), .A2(n8082), .B1(n24552), .B2(n8274), .ZN(
        n23539) );
  AOI22_X1 U22909 ( .A1(n24534), .A2(n8338), .B1(n24528), .B2(n23878), .ZN(
        n23540) );
  AOI22_X1 U22910 ( .A1(n24559), .A2(n8081), .B1(n24553), .B2(n8273), .ZN(
        n23521) );
  AOI22_X1 U22911 ( .A1(n24535), .A2(n8337), .B1(n24529), .B2(n23880), .ZN(
        n23522) );
  AOI22_X1 U22912 ( .A1(n24559), .A2(n8080), .B1(n24553), .B2(n8272), .ZN(
        n23503) );
  AOI22_X1 U22913 ( .A1(n24535), .A2(n8336), .B1(n24529), .B2(n23882), .ZN(
        n23504) );
  AOI22_X1 U22914 ( .A1(n24559), .A2(n8079), .B1(n24553), .B2(n8271), .ZN(
        n23485) );
  AOI22_X1 U22915 ( .A1(n24535), .A2(n8335), .B1(n24529), .B2(n23884), .ZN(
        n23486) );
  AOI22_X1 U22916 ( .A1(n24559), .A2(n8078), .B1(n24553), .B2(n8270), .ZN(
        n23467) );
  AOI22_X1 U22917 ( .A1(n24535), .A2(n8334), .B1(n24529), .B2(n23886), .ZN(
        n23468) );
  AOI22_X1 U22918 ( .A1(n24559), .A2(n8077), .B1(n24553), .B2(n8269), .ZN(
        n23449) );
  AOI22_X1 U22919 ( .A1(n24535), .A2(n8333), .B1(n24529), .B2(n23888), .ZN(
        n23450) );
  AOI22_X1 U22920 ( .A1(n24559), .A2(n8076), .B1(n24553), .B2(n8268), .ZN(
        n23431) );
  AOI22_X1 U22921 ( .A1(n24535), .A2(n8332), .B1(n24529), .B2(n23890), .ZN(
        n23432) );
  AOI22_X1 U22922 ( .A1(n24559), .A2(n8075), .B1(n24553), .B2(n8267), .ZN(
        n23413) );
  AOI22_X1 U22923 ( .A1(n24535), .A2(n8331), .B1(n24529), .B2(n23892), .ZN(
        n23414) );
  AOI22_X1 U22924 ( .A1(n24559), .A2(n8074), .B1(n24553), .B2(n8266), .ZN(
        n23395) );
  AOI22_X1 U22925 ( .A1(n24535), .A2(n8330), .B1(n24529), .B2(n23894), .ZN(
        n23396) );
  AOI22_X1 U22926 ( .A1(n24559), .A2(n8073), .B1(n24553), .B2(n8265), .ZN(
        n23377) );
  AOI22_X1 U22927 ( .A1(n24535), .A2(n8329), .B1(n24529), .B2(n23896), .ZN(
        n23378) );
  AOI22_X1 U22928 ( .A1(n24559), .A2(n8072), .B1(n24553), .B2(n8264), .ZN(
        n23359) );
  AOI22_X1 U22929 ( .A1(n24535), .A2(n8328), .B1(n24529), .B2(n23898), .ZN(
        n23360) );
  AOI22_X1 U22930 ( .A1(n24559), .A2(n8071), .B1(n24553), .B2(n8263), .ZN(
        n23341) );
  AOI22_X1 U22931 ( .A1(n24535), .A2(n8327), .B1(n24529), .B2(n23900), .ZN(
        n23342) );
  AOI22_X1 U22932 ( .A1(n24559), .A2(n8070), .B1(n24553), .B2(n8262), .ZN(
        n23323) );
  AOI22_X1 U22933 ( .A1(n24535), .A2(n8326), .B1(n24529), .B2(n23902), .ZN(
        n23324) );
  AOI22_X1 U22934 ( .A1(n24560), .A2(n8069), .B1(n24554), .B2(n8261), .ZN(
        n23305) );
  AOI22_X1 U22935 ( .A1(n24536), .A2(n8325), .B1(n24530), .B2(n23904), .ZN(
        n23306) );
  AOI22_X1 U22936 ( .A1(n24560), .A2(n8068), .B1(n24554), .B2(n8260), .ZN(
        n23287) );
  AOI22_X1 U22937 ( .A1(n24536), .A2(n8324), .B1(n24530), .B2(n23906), .ZN(
        n23288) );
  AOI22_X1 U22938 ( .A1(n24560), .A2(n8067), .B1(n24554), .B2(n8259), .ZN(
        n23269) );
  AOI22_X1 U22939 ( .A1(n24536), .A2(n8323), .B1(n24530), .B2(n23908), .ZN(
        n23270) );
  AOI22_X1 U22940 ( .A1(n24560), .A2(n8066), .B1(n24554), .B2(n8258), .ZN(
        n23251) );
  AOI22_X1 U22941 ( .A1(n24536), .A2(n8322), .B1(n24530), .B2(n23910), .ZN(
        n23252) );
  AOI22_X1 U22942 ( .A1(n24560), .A2(n8065), .B1(n24554), .B2(n8257), .ZN(
        n23233) );
  AOI22_X1 U22943 ( .A1(n24536), .A2(n8321), .B1(n24530), .B2(n23912), .ZN(
        n23234) );
  AOI22_X1 U22944 ( .A1(n24560), .A2(n8064), .B1(n24554), .B2(n8256), .ZN(
        n23215) );
  AOI22_X1 U22945 ( .A1(n24536), .A2(n8320), .B1(n24530), .B2(n23914), .ZN(
        n23216) );
  AOI22_X1 U22946 ( .A1(n24560), .A2(n8063), .B1(n24554), .B2(n8255), .ZN(
        n23197) );
  AOI22_X1 U22947 ( .A1(n24536), .A2(n8319), .B1(n24530), .B2(n23916), .ZN(
        n23198) );
  AOI22_X1 U22948 ( .A1(n24560), .A2(n8062), .B1(n24554), .B2(n8254), .ZN(
        n23179) );
  AOI22_X1 U22949 ( .A1(n24536), .A2(n8318), .B1(n24530), .B2(n23918), .ZN(
        n23180) );
  AOI22_X1 U22950 ( .A1(n24560), .A2(n8061), .B1(n24554), .B2(n8253), .ZN(
        n23161) );
  AOI22_X1 U22951 ( .A1(n24536), .A2(n8317), .B1(n24530), .B2(n23920), .ZN(
        n23162) );
  AOI22_X1 U22952 ( .A1(n24560), .A2(n8060), .B1(n24554), .B2(n8252), .ZN(
        n23143) );
  AOI22_X1 U22953 ( .A1(n24536), .A2(n8316), .B1(n24530), .B2(n23922), .ZN(
        n23144) );
  AOI22_X1 U22954 ( .A1(n24560), .A2(n8059), .B1(n24554), .B2(n8251), .ZN(
        n23125) );
  AOI22_X1 U22955 ( .A1(n24536), .A2(n8315), .B1(n24530), .B2(n23924), .ZN(
        n23126) );
  AOI22_X1 U22956 ( .A1(n24560), .A2(n8058), .B1(n24554), .B2(n8250), .ZN(
        n23107) );
  AOI22_X1 U22957 ( .A1(n24536), .A2(n8314), .B1(n24530), .B2(n23926), .ZN(
        n23108) );
  AOI22_X1 U22958 ( .A1(n24561), .A2(n8057), .B1(n24555), .B2(n8249), .ZN(
        n23089) );
  AOI22_X1 U22959 ( .A1(n24537), .A2(n8313), .B1(n24531), .B2(n23928), .ZN(
        n23090) );
  AOI22_X1 U22960 ( .A1(n24561), .A2(n8056), .B1(n24555), .B2(n8248), .ZN(
        n23071) );
  AOI22_X1 U22961 ( .A1(n24537), .A2(n8312), .B1(n24531), .B2(n23930), .ZN(
        n23072) );
  AOI22_X1 U22962 ( .A1(n24561), .A2(n8055), .B1(n24555), .B2(n8247), .ZN(
        n23053) );
  AOI22_X1 U22963 ( .A1(n24537), .A2(n8311), .B1(n24531), .B2(n23932), .ZN(
        n23054) );
  AOI22_X1 U22964 ( .A1(n24561), .A2(n8054), .B1(n24555), .B2(n8246), .ZN(
        n23035) );
  AOI22_X1 U22965 ( .A1(n24537), .A2(n8310), .B1(n24531), .B2(n23934), .ZN(
        n23036) );
  OAI22_X1 U22966 ( .A1(n24831), .A2(n20249), .B1(n24819), .B2(n25359), .ZN(
        n5064) );
  OAI22_X1 U22967 ( .A1(n24831), .A2(n20248), .B1(n24819), .B2(n25362), .ZN(
        n5065) );
  OAI22_X1 U22968 ( .A1(n24831), .A2(n20247), .B1(n24819), .B2(n25365), .ZN(
        n5066) );
  OAI22_X1 U22969 ( .A1(n24831), .A2(n20246), .B1(n24819), .B2(n25368), .ZN(
        n5067) );
  OAI22_X1 U22970 ( .A1(n24831), .A2(n20245), .B1(n24819), .B2(n25371), .ZN(
        n5068) );
  OAI22_X1 U22971 ( .A1(n24830), .A2(n20244), .B1(n24819), .B2(n25374), .ZN(
        n5069) );
  OAI22_X1 U22972 ( .A1(n24830), .A2(n20243), .B1(n24819), .B2(n25377), .ZN(
        n5070) );
  OAI22_X1 U22973 ( .A1(n24830), .A2(n20242), .B1(n24819), .B2(n25380), .ZN(
        n5071) );
  OAI22_X1 U22974 ( .A1(n24830), .A2(n20241), .B1(n24819), .B2(n25383), .ZN(
        n5072) );
  OAI22_X1 U22975 ( .A1(n24830), .A2(n20240), .B1(n24819), .B2(n25386), .ZN(
        n5073) );
  OAI22_X1 U22976 ( .A1(n24829), .A2(n20239), .B1(n24819), .B2(n25389), .ZN(
        n5074) );
  OAI22_X1 U22977 ( .A1(n24829), .A2(n20238), .B1(n24819), .B2(n25392), .ZN(
        n5075) );
  OAI22_X1 U22978 ( .A1(n24829), .A2(n20237), .B1(n24817), .B2(n25395), .ZN(
        n5076) );
  OAI22_X1 U22979 ( .A1(n24829), .A2(n20236), .B1(n24819), .B2(n25398), .ZN(
        n5077) );
  OAI22_X1 U22980 ( .A1(n24829), .A2(n20235), .B1(n24818), .B2(n25401), .ZN(
        n5078) );
  OAI22_X1 U22981 ( .A1(n24828), .A2(n20234), .B1(n24817), .B2(n25404), .ZN(
        n5079) );
  OAI22_X1 U22982 ( .A1(n24828), .A2(n20233), .B1(n24819), .B2(n25407), .ZN(
        n5080) );
  OAI22_X1 U22983 ( .A1(n24828), .A2(n20232), .B1(n24818), .B2(n25410), .ZN(
        n5081) );
  OAI22_X1 U22984 ( .A1(n24828), .A2(n20231), .B1(n24817), .B2(n25413), .ZN(
        n5082) );
  OAI22_X1 U22985 ( .A1(n24828), .A2(n20230), .B1(n24819), .B2(n25416), .ZN(
        n5083) );
  OAI22_X1 U22986 ( .A1(n24827), .A2(n20229), .B1(n24818), .B2(n25419), .ZN(
        n5084) );
  OAI22_X1 U22987 ( .A1(n24827), .A2(n20228), .B1(n24817), .B2(n25422), .ZN(
        n5085) );
  OAI22_X1 U22988 ( .A1(n24827), .A2(n20227), .B1(n24819), .B2(n25425), .ZN(
        n5086) );
  OAI22_X1 U22989 ( .A1(n24827), .A2(n20226), .B1(n24818), .B2(n25428), .ZN(
        n5087) );
  OAI22_X1 U22990 ( .A1(n24827), .A2(n20225), .B1(n24818), .B2(n25431), .ZN(
        n5088) );
  OAI22_X1 U22991 ( .A1(n24826), .A2(n20224), .B1(n24817), .B2(n25434), .ZN(
        n5089) );
  OAI22_X1 U22992 ( .A1(n24826), .A2(n20223), .B1(n24819), .B2(n25437), .ZN(
        n5090) );
  OAI22_X1 U22993 ( .A1(n24826), .A2(n20222), .B1(n24818), .B2(n25440), .ZN(
        n5091) );
  OAI22_X1 U22994 ( .A1(n24826), .A2(n20221), .B1(n24818), .B2(n25443), .ZN(
        n5092) );
  OAI22_X1 U22995 ( .A1(n24826), .A2(n20220), .B1(n24817), .B2(n25446), .ZN(
        n5093) );
  OAI22_X1 U22996 ( .A1(n24825), .A2(n20219), .B1(n24819), .B2(n25449), .ZN(
        n5094) );
  OAI22_X1 U22997 ( .A1(n24825), .A2(n20218), .B1(n24817), .B2(n25452), .ZN(
        n5095) );
  OAI22_X1 U22998 ( .A1(n24825), .A2(n20217), .B1(n24818), .B2(n25455), .ZN(
        n5096) );
  OAI22_X1 U22999 ( .A1(n24825), .A2(n20216), .B1(n24817), .B2(n25458), .ZN(
        n5097) );
  OAI22_X1 U23000 ( .A1(n24825), .A2(n20215), .B1(n24819), .B2(n25461), .ZN(
        n5098) );
  OAI22_X1 U23001 ( .A1(n24824), .A2(n20214), .B1(n24819), .B2(n25464), .ZN(
        n5099) );
  OAI22_X1 U23002 ( .A1(n24832), .A2(n20526), .B1(n24818), .B2(n25347), .ZN(
        n5060) );
  OAI22_X1 U23003 ( .A1(n24832), .A2(n20189), .B1(n24817), .B2(n25350), .ZN(
        n5061) );
  OAI22_X1 U23004 ( .A1(n24832), .A2(n20188), .B1(n24819), .B2(n25353), .ZN(
        n5062) );
  OAI22_X1 U23005 ( .A1(n24832), .A2(n20187), .B1(n24818), .B2(n25356), .ZN(
        n5063) );
  OAI22_X1 U23006 ( .A1(n25337), .A2(n25450), .B1(n93), .B2(n25327), .ZN(n7015) );
  OAI22_X1 U23007 ( .A1(n25337), .A2(n25462), .B1(n89), .B2(n21255), .ZN(n7019) );
  OAI22_X1 U23008 ( .A1(n25338), .A2(n25468), .B1(n87), .B2(n25327), .ZN(n7021) );
  OAI22_X1 U23009 ( .A1(n25338), .A2(n25474), .B1(n85), .B2(n21255), .ZN(n7023) );
  OAI22_X1 U23010 ( .A1(n25338), .A2(n25477), .B1(n84), .B2(n25327), .ZN(n7024) );
  OAI22_X1 U23011 ( .A1(n25339), .A2(n25480), .B1(n83), .B2(n21255), .ZN(n7025) );
  OAI22_X1 U23012 ( .A1(n25339), .A2(n25483), .B1(n82), .B2(n25327), .ZN(n7026) );
  OAI22_X1 U23013 ( .A1(n25339), .A2(n25486), .B1(n81), .B2(n21255), .ZN(n7027) );
  OAI22_X1 U23014 ( .A1(n25339), .A2(n25489), .B1(n80), .B2(n25327), .ZN(n7028) );
  OAI22_X1 U23015 ( .A1(n25339), .A2(n25492), .B1(n79), .B2(n21255), .ZN(n7029) );
  OAI22_X1 U23016 ( .A1(n25340), .A2(n25495), .B1(n78), .B2(n25327), .ZN(n7030) );
  OAI22_X1 U23017 ( .A1(n25340), .A2(n25498), .B1(n77), .B2(n21255), .ZN(n7031) );
  OAI22_X1 U23018 ( .A1(n25262), .A2(n25345), .B1(n17410), .B2(n25260), .ZN(
        n6724) );
  OAI22_X1 U23019 ( .A1(n25262), .A2(n25348), .B1(n17407), .B2(n25260), .ZN(
        n6725) );
  OAI22_X1 U23020 ( .A1(n25262), .A2(n25351), .B1(n17404), .B2(n25260), .ZN(
        n6726) );
  OAI22_X1 U23021 ( .A1(n25262), .A2(n25354), .B1(n17401), .B2(n25260), .ZN(
        n6727) );
  OAI22_X1 U23022 ( .A1(n25262), .A2(n25357), .B1(n17398), .B2(n25260), .ZN(
        n6728) );
  OAI22_X1 U23023 ( .A1(n25263), .A2(n25360), .B1(n17395), .B2(n25260), .ZN(
        n6729) );
  OAI22_X1 U23024 ( .A1(n25263), .A2(n25363), .B1(n17392), .B2(n25260), .ZN(
        n6730) );
  OAI22_X1 U23025 ( .A1(n25263), .A2(n25366), .B1(n17389), .B2(n25260), .ZN(
        n6731) );
  OAI22_X1 U23026 ( .A1(n25263), .A2(n25369), .B1(n17386), .B2(n25260), .ZN(
        n6732) );
  OAI22_X1 U23027 ( .A1(n25263), .A2(n25372), .B1(n17383), .B2(n25260), .ZN(
        n6733) );
  OAI22_X1 U23028 ( .A1(n25264), .A2(n25375), .B1(n17380), .B2(n25260), .ZN(
        n6734) );
  OAI22_X1 U23029 ( .A1(n25264), .A2(n25378), .B1(n17377), .B2(n25260), .ZN(
        n6735) );
  OAI22_X1 U23030 ( .A1(n25264), .A2(n25381), .B1(n17374), .B2(n25261), .ZN(
        n6736) );
  OAI22_X1 U23031 ( .A1(n25264), .A2(n25384), .B1(n17371), .B2(n25261), .ZN(
        n6737) );
  OAI22_X1 U23032 ( .A1(n25264), .A2(n25387), .B1(n17368), .B2(n25261), .ZN(
        n6738) );
  OAI22_X1 U23033 ( .A1(n25265), .A2(n25390), .B1(n17365), .B2(n25261), .ZN(
        n6739) );
  OAI22_X1 U23034 ( .A1(n25265), .A2(n25393), .B1(n17362), .B2(n25261), .ZN(
        n6740) );
  OAI22_X1 U23035 ( .A1(n25265), .A2(n25396), .B1(n17359), .B2(n25261), .ZN(
        n6741) );
  OAI22_X1 U23036 ( .A1(n25265), .A2(n25399), .B1(n17356), .B2(n25261), .ZN(
        n6742) );
  OAI22_X1 U23037 ( .A1(n25265), .A2(n25402), .B1(n17353), .B2(n25261), .ZN(
        n6743) );
  OAI22_X1 U23038 ( .A1(n25266), .A2(n25405), .B1(n17350), .B2(n25261), .ZN(
        n6744) );
  OAI22_X1 U23039 ( .A1(n25266), .A2(n25408), .B1(n17347), .B2(n25261), .ZN(
        n6745) );
  OAI22_X1 U23040 ( .A1(n25266), .A2(n25411), .B1(n17344), .B2(n25261), .ZN(
        n6746) );
  OAI22_X1 U23041 ( .A1(n25266), .A2(n25414), .B1(n17341), .B2(n25261), .ZN(
        n6747) );
  OAI22_X1 U23042 ( .A1(n25177), .A2(n25345), .B1(n7554), .B2(n25175), .ZN(
        n6404) );
  OAI22_X1 U23043 ( .A1(n25177), .A2(n25348), .B1(n7552), .B2(n25175), .ZN(
        n6405) );
  OAI22_X1 U23044 ( .A1(n25177), .A2(n25351), .B1(n7550), .B2(n25175), .ZN(
        n6406) );
  OAI22_X1 U23045 ( .A1(n25177), .A2(n25354), .B1(n7548), .B2(n25175), .ZN(
        n6407) );
  OAI22_X1 U23046 ( .A1(n25177), .A2(n25357), .B1(n7546), .B2(n25175), .ZN(
        n6408) );
  OAI22_X1 U23047 ( .A1(n25178), .A2(n25360), .B1(n7544), .B2(n25175), .ZN(
        n6409) );
  OAI22_X1 U23048 ( .A1(n25178), .A2(n25363), .B1(n7542), .B2(n25175), .ZN(
        n6410) );
  OAI22_X1 U23049 ( .A1(n25178), .A2(n25366), .B1(n7540), .B2(n25175), .ZN(
        n6411) );
  OAI22_X1 U23050 ( .A1(n25178), .A2(n25369), .B1(n7538), .B2(n25175), .ZN(
        n6412) );
  OAI22_X1 U23051 ( .A1(n25178), .A2(n25372), .B1(n7536), .B2(n25175), .ZN(
        n6413) );
  OAI22_X1 U23052 ( .A1(n25179), .A2(n25375), .B1(n7534), .B2(n25175), .ZN(
        n6414) );
  OAI22_X1 U23053 ( .A1(n25179), .A2(n25378), .B1(n7532), .B2(n25175), .ZN(
        n6415) );
  OAI22_X1 U23054 ( .A1(n25179), .A2(n25381), .B1(n7530), .B2(n25176), .ZN(
        n6416) );
  OAI22_X1 U23055 ( .A1(n25179), .A2(n25384), .B1(n7528), .B2(n25176), .ZN(
        n6417) );
  OAI22_X1 U23056 ( .A1(n25179), .A2(n25387), .B1(n7526), .B2(n25176), .ZN(
        n6418) );
  OAI22_X1 U23057 ( .A1(n25180), .A2(n25390), .B1(n7524), .B2(n25176), .ZN(
        n6419) );
  OAI22_X1 U23058 ( .A1(n25180), .A2(n25393), .B1(n7522), .B2(n25176), .ZN(
        n6420) );
  OAI22_X1 U23059 ( .A1(n25180), .A2(n25396), .B1(n7520), .B2(n25176), .ZN(
        n6421) );
  OAI22_X1 U23060 ( .A1(n25180), .A2(n25399), .B1(n7518), .B2(n25176), .ZN(
        n6422) );
  OAI22_X1 U23061 ( .A1(n25180), .A2(n25402), .B1(n7516), .B2(n25176), .ZN(
        n6423) );
  OAI22_X1 U23062 ( .A1(n25181), .A2(n25405), .B1(n7514), .B2(n25176), .ZN(
        n6424) );
  OAI22_X1 U23063 ( .A1(n25181), .A2(n25408), .B1(n7512), .B2(n25176), .ZN(
        n6425) );
  OAI22_X1 U23064 ( .A1(n25181), .A2(n25411), .B1(n7510), .B2(n25176), .ZN(
        n6426) );
  OAI22_X1 U23065 ( .A1(n25181), .A2(n25414), .B1(n7508), .B2(n25176), .ZN(
        n6427) );
  OAI22_X1 U23066 ( .A1(n25092), .A2(n25346), .B1(n7426), .B2(n25090), .ZN(
        n6084) );
  OAI22_X1 U23067 ( .A1(n25092), .A2(n25349), .B1(n7424), .B2(n25090), .ZN(
        n6085) );
  OAI22_X1 U23068 ( .A1(n25092), .A2(n25352), .B1(n7422), .B2(n25090), .ZN(
        n6086) );
  OAI22_X1 U23069 ( .A1(n25092), .A2(n25355), .B1(n7420), .B2(n25090), .ZN(
        n6087) );
  OAI22_X1 U23070 ( .A1(n25092), .A2(n25358), .B1(n7418), .B2(n25090), .ZN(
        n6088) );
  OAI22_X1 U23071 ( .A1(n25093), .A2(n25361), .B1(n7416), .B2(n25090), .ZN(
        n6089) );
  OAI22_X1 U23072 ( .A1(n25093), .A2(n25364), .B1(n7414), .B2(n25090), .ZN(
        n6090) );
  OAI22_X1 U23073 ( .A1(n25093), .A2(n25367), .B1(n7412), .B2(n25090), .ZN(
        n6091) );
  OAI22_X1 U23074 ( .A1(n25093), .A2(n25370), .B1(n7410), .B2(n25090), .ZN(
        n6092) );
  OAI22_X1 U23075 ( .A1(n25093), .A2(n25373), .B1(n7408), .B2(n25090), .ZN(
        n6093) );
  OAI22_X1 U23076 ( .A1(n25094), .A2(n25376), .B1(n7406), .B2(n25090), .ZN(
        n6094) );
  OAI22_X1 U23077 ( .A1(n25094), .A2(n25379), .B1(n7404), .B2(n25090), .ZN(
        n6095) );
  OAI22_X1 U23078 ( .A1(n25094), .A2(n25382), .B1(n7402), .B2(n25091), .ZN(
        n6096) );
  OAI22_X1 U23079 ( .A1(n25094), .A2(n25385), .B1(n7400), .B2(n25091), .ZN(
        n6097) );
  OAI22_X1 U23080 ( .A1(n25094), .A2(n25388), .B1(n7398), .B2(n25091), .ZN(
        n6098) );
  OAI22_X1 U23081 ( .A1(n25095), .A2(n25391), .B1(n7396), .B2(n25091), .ZN(
        n6099) );
  OAI22_X1 U23082 ( .A1(n25095), .A2(n25394), .B1(n7394), .B2(n25091), .ZN(
        n6100) );
  OAI22_X1 U23083 ( .A1(n25095), .A2(n25397), .B1(n7392), .B2(n25091), .ZN(
        n6101) );
  OAI22_X1 U23084 ( .A1(n25095), .A2(n25400), .B1(n7390), .B2(n25091), .ZN(
        n6102) );
  OAI22_X1 U23085 ( .A1(n25095), .A2(n25403), .B1(n7388), .B2(n25091), .ZN(
        n6103) );
  OAI22_X1 U23086 ( .A1(n25096), .A2(n25406), .B1(n7386), .B2(n25091), .ZN(
        n6104) );
  OAI22_X1 U23087 ( .A1(n25096), .A2(n25409), .B1(n7384), .B2(n25091), .ZN(
        n6105) );
  OAI22_X1 U23088 ( .A1(n25096), .A2(n25412), .B1(n7382), .B2(n25091), .ZN(
        n6106) );
  OAI22_X1 U23089 ( .A1(n25096), .A2(n25415), .B1(n7380), .B2(n25091), .ZN(
        n6107) );
  OAI22_X1 U23090 ( .A1(n25041), .A2(n25346), .B1(n8861), .B2(n25039), .ZN(
        n5892) );
  OAI22_X1 U23091 ( .A1(n25041), .A2(n25349), .B1(n8859), .B2(n25039), .ZN(
        n5893) );
  OAI22_X1 U23092 ( .A1(n25041), .A2(n25352), .B1(n8857), .B2(n25039), .ZN(
        n5894) );
  OAI22_X1 U23093 ( .A1(n25041), .A2(n25355), .B1(n8855), .B2(n25039), .ZN(
        n5895) );
  OAI22_X1 U23094 ( .A1(n25041), .A2(n25358), .B1(n8853), .B2(n25039), .ZN(
        n5896) );
  OAI22_X1 U23095 ( .A1(n25042), .A2(n25361), .B1(n8851), .B2(n25039), .ZN(
        n5897) );
  OAI22_X1 U23096 ( .A1(n25042), .A2(n25364), .B1(n8849), .B2(n25039), .ZN(
        n5898) );
  OAI22_X1 U23097 ( .A1(n25042), .A2(n25367), .B1(n8847), .B2(n25039), .ZN(
        n5899) );
  OAI22_X1 U23098 ( .A1(n25042), .A2(n25370), .B1(n8845), .B2(n25039), .ZN(
        n5900) );
  OAI22_X1 U23099 ( .A1(n25042), .A2(n25373), .B1(n8843), .B2(n25039), .ZN(
        n5901) );
  OAI22_X1 U23100 ( .A1(n25043), .A2(n25376), .B1(n8841), .B2(n25039), .ZN(
        n5902) );
  OAI22_X1 U23101 ( .A1(n25043), .A2(n25379), .B1(n8839), .B2(n25039), .ZN(
        n5903) );
  OAI22_X1 U23102 ( .A1(n25043), .A2(n25382), .B1(n8837), .B2(n25040), .ZN(
        n5904) );
  OAI22_X1 U23103 ( .A1(n25043), .A2(n25385), .B1(n8835), .B2(n25040), .ZN(
        n5905) );
  OAI22_X1 U23104 ( .A1(n25043), .A2(n25388), .B1(n8833), .B2(n25040), .ZN(
        n5906) );
  OAI22_X1 U23105 ( .A1(n25044), .A2(n25391), .B1(n8831), .B2(n25040), .ZN(
        n5907) );
  OAI22_X1 U23106 ( .A1(n25044), .A2(n25394), .B1(n8829), .B2(n25040), .ZN(
        n5908) );
  OAI22_X1 U23107 ( .A1(n25044), .A2(n25397), .B1(n8827), .B2(n25040), .ZN(
        n5909) );
  OAI22_X1 U23108 ( .A1(n25044), .A2(n25400), .B1(n8825), .B2(n25040), .ZN(
        n5910) );
  OAI22_X1 U23109 ( .A1(n25044), .A2(n25403), .B1(n8823), .B2(n25040), .ZN(
        n5911) );
  OAI22_X1 U23110 ( .A1(n25045), .A2(n25406), .B1(n8821), .B2(n25040), .ZN(
        n5912) );
  OAI22_X1 U23111 ( .A1(n25045), .A2(n25409), .B1(n8819), .B2(n25040), .ZN(
        n5913) );
  OAI22_X1 U23112 ( .A1(n25045), .A2(n25412), .B1(n8817), .B2(n25040), .ZN(
        n5914) );
  OAI22_X1 U23113 ( .A1(n25045), .A2(n25415), .B1(n8815), .B2(n25040), .ZN(
        n5915) );
  OAI22_X1 U23114 ( .A1(n25024), .A2(n25346), .B1(n8989), .B2(n25022), .ZN(
        n5828) );
  OAI22_X1 U23115 ( .A1(n25024), .A2(n25349), .B1(n8987), .B2(n25022), .ZN(
        n5829) );
  OAI22_X1 U23116 ( .A1(n25024), .A2(n25352), .B1(n8985), .B2(n25022), .ZN(
        n5830) );
  OAI22_X1 U23117 ( .A1(n25024), .A2(n25355), .B1(n8983), .B2(n25022), .ZN(
        n5831) );
  OAI22_X1 U23118 ( .A1(n25024), .A2(n25358), .B1(n8981), .B2(n25022), .ZN(
        n5832) );
  OAI22_X1 U23119 ( .A1(n25025), .A2(n25361), .B1(n8979), .B2(n25022), .ZN(
        n5833) );
  OAI22_X1 U23120 ( .A1(n25025), .A2(n25364), .B1(n8977), .B2(n25022), .ZN(
        n5834) );
  OAI22_X1 U23121 ( .A1(n25025), .A2(n25367), .B1(n8975), .B2(n25022), .ZN(
        n5835) );
  OAI22_X1 U23122 ( .A1(n25025), .A2(n25370), .B1(n8973), .B2(n25022), .ZN(
        n5836) );
  OAI22_X1 U23123 ( .A1(n25025), .A2(n25373), .B1(n8971), .B2(n25022), .ZN(
        n5837) );
  OAI22_X1 U23124 ( .A1(n25026), .A2(n25376), .B1(n8969), .B2(n25022), .ZN(
        n5838) );
  OAI22_X1 U23125 ( .A1(n25026), .A2(n25379), .B1(n8967), .B2(n25022), .ZN(
        n5839) );
  OAI22_X1 U23126 ( .A1(n25026), .A2(n25382), .B1(n8965), .B2(n25023), .ZN(
        n5840) );
  OAI22_X1 U23127 ( .A1(n25026), .A2(n25385), .B1(n8963), .B2(n25023), .ZN(
        n5841) );
  OAI22_X1 U23128 ( .A1(n25026), .A2(n25388), .B1(n8961), .B2(n25023), .ZN(
        n5842) );
  OAI22_X1 U23129 ( .A1(n25027), .A2(n25391), .B1(n8959), .B2(n25023), .ZN(
        n5843) );
  OAI22_X1 U23130 ( .A1(n25027), .A2(n25394), .B1(n8957), .B2(n25023), .ZN(
        n5844) );
  OAI22_X1 U23131 ( .A1(n25027), .A2(n25397), .B1(n8955), .B2(n25023), .ZN(
        n5845) );
  OAI22_X1 U23132 ( .A1(n25027), .A2(n25400), .B1(n8953), .B2(n25023), .ZN(
        n5846) );
  OAI22_X1 U23133 ( .A1(n25027), .A2(n25403), .B1(n8951), .B2(n25023), .ZN(
        n5847) );
  OAI22_X1 U23134 ( .A1(n25028), .A2(n25406), .B1(n8949), .B2(n25023), .ZN(
        n5848) );
  OAI22_X1 U23135 ( .A1(n25028), .A2(n25409), .B1(n8947), .B2(n25023), .ZN(
        n5849) );
  OAI22_X1 U23136 ( .A1(n25028), .A2(n25412), .B1(n8945), .B2(n25023), .ZN(
        n5850) );
  OAI22_X1 U23137 ( .A1(n25028), .A2(n25415), .B1(n8943), .B2(n25023), .ZN(
        n5851) );
  OAI22_X1 U23138 ( .A1(n24854), .A2(n25347), .B1(n8988), .B2(n24852), .ZN(
        n5188) );
  OAI22_X1 U23139 ( .A1(n24854), .A2(n25350), .B1(n8986), .B2(n24852), .ZN(
        n5189) );
  OAI22_X1 U23140 ( .A1(n24854), .A2(n25353), .B1(n8984), .B2(n24852), .ZN(
        n5190) );
  OAI22_X1 U23141 ( .A1(n24854), .A2(n25356), .B1(n8982), .B2(n24852), .ZN(
        n5191) );
  OAI22_X1 U23142 ( .A1(n24854), .A2(n25359), .B1(n8980), .B2(n24852), .ZN(
        n5192) );
  OAI22_X1 U23143 ( .A1(n24855), .A2(n25362), .B1(n8978), .B2(n24852), .ZN(
        n5193) );
  OAI22_X1 U23144 ( .A1(n24855), .A2(n25365), .B1(n8976), .B2(n24852), .ZN(
        n5194) );
  OAI22_X1 U23145 ( .A1(n24855), .A2(n25368), .B1(n8974), .B2(n24852), .ZN(
        n5195) );
  OAI22_X1 U23146 ( .A1(n24855), .A2(n25371), .B1(n8972), .B2(n24852), .ZN(
        n5196) );
  OAI22_X1 U23147 ( .A1(n24855), .A2(n25374), .B1(n8970), .B2(n24852), .ZN(
        n5197) );
  OAI22_X1 U23148 ( .A1(n24856), .A2(n25377), .B1(n8968), .B2(n24852), .ZN(
        n5198) );
  OAI22_X1 U23149 ( .A1(n24856), .A2(n25380), .B1(n8966), .B2(n24852), .ZN(
        n5199) );
  OAI22_X1 U23150 ( .A1(n24856), .A2(n25383), .B1(n8964), .B2(n24853), .ZN(
        n5200) );
  OAI22_X1 U23151 ( .A1(n24856), .A2(n25386), .B1(n8962), .B2(n24853), .ZN(
        n5201) );
  OAI22_X1 U23152 ( .A1(n24856), .A2(n25389), .B1(n8960), .B2(n24853), .ZN(
        n5202) );
  OAI22_X1 U23153 ( .A1(n24857), .A2(n25392), .B1(n8958), .B2(n24853), .ZN(
        n5203) );
  OAI22_X1 U23154 ( .A1(n24857), .A2(n25395), .B1(n8956), .B2(n24853), .ZN(
        n5204) );
  OAI22_X1 U23155 ( .A1(n24857), .A2(n25398), .B1(n8954), .B2(n24853), .ZN(
        n5205) );
  OAI22_X1 U23156 ( .A1(n24857), .A2(n25401), .B1(n8952), .B2(n24853), .ZN(
        n5206) );
  OAI22_X1 U23157 ( .A1(n24857), .A2(n25404), .B1(n8950), .B2(n24853), .ZN(
        n5207) );
  OAI22_X1 U23158 ( .A1(n24858), .A2(n25407), .B1(n8948), .B2(n24853), .ZN(
        n5208) );
  OAI22_X1 U23159 ( .A1(n24858), .A2(n25410), .B1(n8946), .B2(n24853), .ZN(
        n5209) );
  OAI22_X1 U23160 ( .A1(n24858), .A2(n25413), .B1(n8944), .B2(n24853), .ZN(
        n5210) );
  OAI22_X1 U23161 ( .A1(n24858), .A2(n25416), .B1(n8942), .B2(n24853), .ZN(
        n5211) );
  OAI22_X1 U23162 ( .A1(n24922), .A2(n25347), .B1(n7427), .B2(n24920), .ZN(
        n5444) );
  OAI22_X1 U23163 ( .A1(n24922), .A2(n25350), .B1(n7425), .B2(n24920), .ZN(
        n5445) );
  OAI22_X1 U23164 ( .A1(n24922), .A2(n25353), .B1(n7423), .B2(n24920), .ZN(
        n5446) );
  OAI22_X1 U23165 ( .A1(n24922), .A2(n25356), .B1(n7421), .B2(n24920), .ZN(
        n5447) );
  OAI22_X1 U23166 ( .A1(n24922), .A2(n25359), .B1(n7419), .B2(n24920), .ZN(
        n5448) );
  OAI22_X1 U23167 ( .A1(n24923), .A2(n25362), .B1(n7417), .B2(n24920), .ZN(
        n5449) );
  OAI22_X1 U23168 ( .A1(n24923), .A2(n25365), .B1(n7415), .B2(n24920), .ZN(
        n5450) );
  OAI22_X1 U23169 ( .A1(n24923), .A2(n25368), .B1(n7413), .B2(n24920), .ZN(
        n5451) );
  OAI22_X1 U23170 ( .A1(n24923), .A2(n25371), .B1(n7411), .B2(n24920), .ZN(
        n5452) );
  OAI22_X1 U23171 ( .A1(n24923), .A2(n25374), .B1(n7409), .B2(n24920), .ZN(
        n5453) );
  OAI22_X1 U23172 ( .A1(n24924), .A2(n25377), .B1(n7407), .B2(n24920), .ZN(
        n5454) );
  OAI22_X1 U23173 ( .A1(n24924), .A2(n25380), .B1(n7405), .B2(n24920), .ZN(
        n5455) );
  OAI22_X1 U23174 ( .A1(n24924), .A2(n25383), .B1(n7403), .B2(n24921), .ZN(
        n5456) );
  OAI22_X1 U23175 ( .A1(n24924), .A2(n25386), .B1(n7401), .B2(n24921), .ZN(
        n5457) );
  OAI22_X1 U23176 ( .A1(n24924), .A2(n25389), .B1(n7399), .B2(n24921), .ZN(
        n5458) );
  OAI22_X1 U23177 ( .A1(n24925), .A2(n25392), .B1(n7397), .B2(n24921), .ZN(
        n5459) );
  OAI22_X1 U23178 ( .A1(n24925), .A2(n25395), .B1(n7395), .B2(n24921), .ZN(
        n5460) );
  OAI22_X1 U23179 ( .A1(n24925), .A2(n25398), .B1(n7393), .B2(n24921), .ZN(
        n5461) );
  OAI22_X1 U23180 ( .A1(n24925), .A2(n25401), .B1(n7391), .B2(n24921), .ZN(
        n5462) );
  OAI22_X1 U23181 ( .A1(n24925), .A2(n25404), .B1(n7389), .B2(n24921), .ZN(
        n5463) );
  OAI22_X1 U23182 ( .A1(n24926), .A2(n25407), .B1(n7387), .B2(n24921), .ZN(
        n5464) );
  OAI22_X1 U23183 ( .A1(n24926), .A2(n25410), .B1(n7385), .B2(n24921), .ZN(
        n5465) );
  OAI22_X1 U23184 ( .A1(n24926), .A2(n25413), .B1(n7383), .B2(n24921), .ZN(
        n5466) );
  OAI22_X1 U23185 ( .A1(n24926), .A2(n25416), .B1(n7381), .B2(n24921), .ZN(
        n5467) );
  OAI22_X1 U23186 ( .A1(n24956), .A2(n25346), .B1(n9245), .B2(n24954), .ZN(
        n5572) );
  OAI22_X1 U23187 ( .A1(n24956), .A2(n25349), .B1(n9243), .B2(n24954), .ZN(
        n5573) );
  OAI22_X1 U23188 ( .A1(n24956), .A2(n25352), .B1(n9241), .B2(n24954), .ZN(
        n5574) );
  OAI22_X1 U23189 ( .A1(n24956), .A2(n25355), .B1(n9239), .B2(n24954), .ZN(
        n5575) );
  OAI22_X1 U23190 ( .A1(n24956), .A2(n25358), .B1(n9237), .B2(n24954), .ZN(
        n5576) );
  OAI22_X1 U23191 ( .A1(n24957), .A2(n25361), .B1(n9235), .B2(n24954), .ZN(
        n5577) );
  OAI22_X1 U23192 ( .A1(n24957), .A2(n25364), .B1(n9233), .B2(n24954), .ZN(
        n5578) );
  OAI22_X1 U23193 ( .A1(n24957), .A2(n25367), .B1(n9231), .B2(n24954), .ZN(
        n5579) );
  OAI22_X1 U23194 ( .A1(n24957), .A2(n25370), .B1(n9229), .B2(n24954), .ZN(
        n5580) );
  OAI22_X1 U23195 ( .A1(n24957), .A2(n25373), .B1(n9227), .B2(n24954), .ZN(
        n5581) );
  OAI22_X1 U23196 ( .A1(n24958), .A2(n25376), .B1(n9225), .B2(n24954), .ZN(
        n5582) );
  OAI22_X1 U23197 ( .A1(n24958), .A2(n25379), .B1(n9223), .B2(n24954), .ZN(
        n5583) );
  OAI22_X1 U23198 ( .A1(n24958), .A2(n25382), .B1(n9221), .B2(n24955), .ZN(
        n5584) );
  OAI22_X1 U23199 ( .A1(n24958), .A2(n25385), .B1(n9219), .B2(n24955), .ZN(
        n5585) );
  OAI22_X1 U23200 ( .A1(n24958), .A2(n25388), .B1(n9217), .B2(n24955), .ZN(
        n5586) );
  OAI22_X1 U23201 ( .A1(n24959), .A2(n25391), .B1(n9215), .B2(n24955), .ZN(
        n5587) );
  OAI22_X1 U23202 ( .A1(n24959), .A2(n25394), .B1(n9213), .B2(n24955), .ZN(
        n5588) );
  OAI22_X1 U23203 ( .A1(n24959), .A2(n25397), .B1(n9211), .B2(n24955), .ZN(
        n5589) );
  OAI22_X1 U23204 ( .A1(n24959), .A2(n25400), .B1(n9209), .B2(n24955), .ZN(
        n5590) );
  OAI22_X1 U23205 ( .A1(n24959), .A2(n25403), .B1(n9207), .B2(n24955), .ZN(
        n5591) );
  OAI22_X1 U23206 ( .A1(n24960), .A2(n25406), .B1(n9205), .B2(n24955), .ZN(
        n5592) );
  OAI22_X1 U23207 ( .A1(n24960), .A2(n25409), .B1(n9203), .B2(n24955), .ZN(
        n5593) );
  OAI22_X1 U23208 ( .A1(n24960), .A2(n25412), .B1(n9201), .B2(n24955), .ZN(
        n5594) );
  OAI22_X1 U23209 ( .A1(n24960), .A2(n25415), .B1(n9199), .B2(n24955), .ZN(
        n5595) );
  OAI22_X1 U23210 ( .A1(n24973), .A2(n25346), .B1(n7555), .B2(n24971), .ZN(
        n5636) );
  OAI22_X1 U23211 ( .A1(n24973), .A2(n25349), .B1(n7553), .B2(n24971), .ZN(
        n5637) );
  OAI22_X1 U23212 ( .A1(n24973), .A2(n25352), .B1(n7551), .B2(n24971), .ZN(
        n5638) );
  OAI22_X1 U23213 ( .A1(n24973), .A2(n25355), .B1(n7549), .B2(n24971), .ZN(
        n5639) );
  OAI22_X1 U23214 ( .A1(n24973), .A2(n25358), .B1(n7547), .B2(n24971), .ZN(
        n5640) );
  OAI22_X1 U23215 ( .A1(n24974), .A2(n25361), .B1(n7545), .B2(n24971), .ZN(
        n5641) );
  OAI22_X1 U23216 ( .A1(n24974), .A2(n25364), .B1(n7543), .B2(n24971), .ZN(
        n5642) );
  OAI22_X1 U23217 ( .A1(n24974), .A2(n25367), .B1(n7541), .B2(n24971), .ZN(
        n5643) );
  OAI22_X1 U23218 ( .A1(n24974), .A2(n25370), .B1(n7539), .B2(n24971), .ZN(
        n5644) );
  OAI22_X1 U23219 ( .A1(n24974), .A2(n25373), .B1(n7537), .B2(n24971), .ZN(
        n5645) );
  OAI22_X1 U23220 ( .A1(n24975), .A2(n25376), .B1(n7535), .B2(n24971), .ZN(
        n5646) );
  OAI22_X1 U23221 ( .A1(n24975), .A2(n25379), .B1(n7533), .B2(n24971), .ZN(
        n5647) );
  OAI22_X1 U23222 ( .A1(n24975), .A2(n25382), .B1(n7531), .B2(n24972), .ZN(
        n5648) );
  OAI22_X1 U23223 ( .A1(n24975), .A2(n25385), .B1(n7529), .B2(n24972), .ZN(
        n5649) );
  OAI22_X1 U23224 ( .A1(n24975), .A2(n25388), .B1(n7527), .B2(n24972), .ZN(
        n5650) );
  OAI22_X1 U23225 ( .A1(n24976), .A2(n25391), .B1(n7525), .B2(n24972), .ZN(
        n5651) );
  OAI22_X1 U23226 ( .A1(n24976), .A2(n25394), .B1(n7523), .B2(n24972), .ZN(
        n5652) );
  OAI22_X1 U23227 ( .A1(n24976), .A2(n25397), .B1(n7521), .B2(n24972), .ZN(
        n5653) );
  OAI22_X1 U23228 ( .A1(n24976), .A2(n25400), .B1(n7519), .B2(n24972), .ZN(
        n5654) );
  OAI22_X1 U23229 ( .A1(n24976), .A2(n25403), .B1(n7517), .B2(n24972), .ZN(
        n5655) );
  OAI22_X1 U23230 ( .A1(n24977), .A2(n25406), .B1(n7515), .B2(n24972), .ZN(
        n5656) );
  OAI22_X1 U23231 ( .A1(n24977), .A2(n25409), .B1(n7513), .B2(n24972), .ZN(
        n5657) );
  OAI22_X1 U23232 ( .A1(n24977), .A2(n25412), .B1(n7511), .B2(n24972), .ZN(
        n5658) );
  OAI22_X1 U23233 ( .A1(n24977), .A2(n25415), .B1(n7509), .B2(n24972), .ZN(
        n5659) );
  OAI22_X1 U23234 ( .A1(n25109), .A2(n25346), .B1(n9116), .B2(n25107), .ZN(
        n6148) );
  OAI22_X1 U23235 ( .A1(n25109), .A2(n25349), .B1(n9114), .B2(n25107), .ZN(
        n6149) );
  OAI22_X1 U23236 ( .A1(n25109), .A2(n25352), .B1(n9112), .B2(n25107), .ZN(
        n6150) );
  OAI22_X1 U23237 ( .A1(n25109), .A2(n25355), .B1(n9110), .B2(n25107), .ZN(
        n6151) );
  OAI22_X1 U23238 ( .A1(n25109), .A2(n25358), .B1(n9108), .B2(n25107), .ZN(
        n6152) );
  OAI22_X1 U23239 ( .A1(n25110), .A2(n25361), .B1(n9106), .B2(n25107), .ZN(
        n6153) );
  OAI22_X1 U23240 ( .A1(n25110), .A2(n25364), .B1(n9104), .B2(n25107), .ZN(
        n6154) );
  OAI22_X1 U23241 ( .A1(n25110), .A2(n25367), .B1(n9102), .B2(n25107), .ZN(
        n6155) );
  OAI22_X1 U23242 ( .A1(n25110), .A2(n25370), .B1(n9100), .B2(n25107), .ZN(
        n6156) );
  OAI22_X1 U23243 ( .A1(n25110), .A2(n25373), .B1(n9098), .B2(n25107), .ZN(
        n6157) );
  OAI22_X1 U23244 ( .A1(n25111), .A2(n25376), .B1(n9096), .B2(n25107), .ZN(
        n6158) );
  OAI22_X1 U23245 ( .A1(n25111), .A2(n25379), .B1(n9094), .B2(n25107), .ZN(
        n6159) );
  OAI22_X1 U23246 ( .A1(n25111), .A2(n25382), .B1(n9092), .B2(n25108), .ZN(
        n6160) );
  OAI22_X1 U23247 ( .A1(n25111), .A2(n25385), .B1(n9090), .B2(n25108), .ZN(
        n6161) );
  OAI22_X1 U23248 ( .A1(n25111), .A2(n25388), .B1(n9088), .B2(n25108), .ZN(
        n6162) );
  OAI22_X1 U23249 ( .A1(n25112), .A2(n25391), .B1(n9086), .B2(n25108), .ZN(
        n6163) );
  OAI22_X1 U23250 ( .A1(n25112), .A2(n25394), .B1(n9084), .B2(n25108), .ZN(
        n6164) );
  OAI22_X1 U23251 ( .A1(n25112), .A2(n25397), .B1(n9082), .B2(n25108), .ZN(
        n6165) );
  OAI22_X1 U23252 ( .A1(n25112), .A2(n25400), .B1(n9080), .B2(n25108), .ZN(
        n6166) );
  OAI22_X1 U23253 ( .A1(n25112), .A2(n25403), .B1(n9078), .B2(n25108), .ZN(
        n6167) );
  OAI22_X1 U23254 ( .A1(n25113), .A2(n25406), .B1(n9076), .B2(n25108), .ZN(
        n6168) );
  OAI22_X1 U23255 ( .A1(n25113), .A2(n25409), .B1(n9074), .B2(n25108), .ZN(
        n6169) );
  OAI22_X1 U23256 ( .A1(n25113), .A2(n25412), .B1(n9072), .B2(n25108), .ZN(
        n6170) );
  OAI22_X1 U23257 ( .A1(n25113), .A2(n25415), .B1(n9070), .B2(n25108), .ZN(
        n6171) );
  OAI22_X1 U23258 ( .A1(n25126), .A2(n25346), .B1(n896), .B2(n25124), .ZN(
        n6212) );
  OAI22_X1 U23259 ( .A1(n25126), .A2(n25349), .B1(n895), .B2(n25124), .ZN(
        n6213) );
  OAI22_X1 U23260 ( .A1(n25126), .A2(n25352), .B1(n894), .B2(n25124), .ZN(
        n6214) );
  OAI22_X1 U23261 ( .A1(n25126), .A2(n25355), .B1(n893), .B2(n25124), .ZN(
        n6215) );
  OAI22_X1 U23262 ( .A1(n25126), .A2(n25358), .B1(n892), .B2(n25124), .ZN(
        n6216) );
  OAI22_X1 U23263 ( .A1(n25127), .A2(n25361), .B1(n891), .B2(n25124), .ZN(
        n6217) );
  OAI22_X1 U23264 ( .A1(n25127), .A2(n25364), .B1(n890), .B2(n25124), .ZN(
        n6218) );
  OAI22_X1 U23265 ( .A1(n25127), .A2(n25367), .B1(n889), .B2(n25124), .ZN(
        n6219) );
  OAI22_X1 U23266 ( .A1(n25127), .A2(n25370), .B1(n888), .B2(n25124), .ZN(
        n6220) );
  OAI22_X1 U23267 ( .A1(n25127), .A2(n25373), .B1(n887), .B2(n25124), .ZN(
        n6221) );
  OAI22_X1 U23268 ( .A1(n25128), .A2(n25376), .B1(n886), .B2(n25124), .ZN(
        n6222) );
  OAI22_X1 U23269 ( .A1(n25128), .A2(n25379), .B1(n885), .B2(n25124), .ZN(
        n6223) );
  OAI22_X1 U23270 ( .A1(n25128), .A2(n25382), .B1(n884), .B2(n25125), .ZN(
        n6224) );
  OAI22_X1 U23271 ( .A1(n25128), .A2(n25385), .B1(n883), .B2(n25125), .ZN(
        n6225) );
  OAI22_X1 U23272 ( .A1(n25128), .A2(n25388), .B1(n882), .B2(n25125), .ZN(
        n6226) );
  OAI22_X1 U23273 ( .A1(n25129), .A2(n25391), .B1(n881), .B2(n25125), .ZN(
        n6227) );
  OAI22_X1 U23274 ( .A1(n25129), .A2(n25394), .B1(n880), .B2(n25125), .ZN(
        n6228) );
  OAI22_X1 U23275 ( .A1(n25129), .A2(n25397), .B1(n879), .B2(n25125), .ZN(
        n6229) );
  OAI22_X1 U23276 ( .A1(n25129), .A2(n25400), .B1(n878), .B2(n25125), .ZN(
        n6230) );
  OAI22_X1 U23277 ( .A1(n25129), .A2(n25403), .B1(n877), .B2(n25125), .ZN(
        n6231) );
  OAI22_X1 U23278 ( .A1(n25130), .A2(n25406), .B1(n876), .B2(n25125), .ZN(
        n6232) );
  OAI22_X1 U23279 ( .A1(n25130), .A2(n25409), .B1(n875), .B2(n25125), .ZN(
        n6233) );
  OAI22_X1 U23280 ( .A1(n25130), .A2(n25412), .B1(n874), .B2(n25125), .ZN(
        n6234) );
  OAI22_X1 U23281 ( .A1(n25130), .A2(n25415), .B1(n873), .B2(n25125), .ZN(
        n6235) );
  OAI22_X1 U23282 ( .A1(n25160), .A2(n25345), .B1(n9244), .B2(n25158), .ZN(
        n6340) );
  OAI22_X1 U23283 ( .A1(n25160), .A2(n25348), .B1(n9242), .B2(n25158), .ZN(
        n6341) );
  OAI22_X1 U23284 ( .A1(n25160), .A2(n25351), .B1(n9240), .B2(n25158), .ZN(
        n6342) );
  OAI22_X1 U23285 ( .A1(n25160), .A2(n25354), .B1(n9238), .B2(n25158), .ZN(
        n6343) );
  OAI22_X1 U23286 ( .A1(n25160), .A2(n25357), .B1(n9236), .B2(n25158), .ZN(
        n6344) );
  OAI22_X1 U23287 ( .A1(n25161), .A2(n25360), .B1(n9234), .B2(n25158), .ZN(
        n6345) );
  OAI22_X1 U23288 ( .A1(n25161), .A2(n25363), .B1(n9232), .B2(n25158), .ZN(
        n6346) );
  OAI22_X1 U23289 ( .A1(n25161), .A2(n25366), .B1(n9230), .B2(n25158), .ZN(
        n6347) );
  OAI22_X1 U23290 ( .A1(n25161), .A2(n25369), .B1(n9228), .B2(n25158), .ZN(
        n6348) );
  OAI22_X1 U23291 ( .A1(n25161), .A2(n25372), .B1(n9226), .B2(n25158), .ZN(
        n6349) );
  OAI22_X1 U23292 ( .A1(n25162), .A2(n25375), .B1(n9224), .B2(n25158), .ZN(
        n6350) );
  OAI22_X1 U23293 ( .A1(n25162), .A2(n25378), .B1(n9222), .B2(n25158), .ZN(
        n6351) );
  OAI22_X1 U23294 ( .A1(n25162), .A2(n25381), .B1(n9220), .B2(n25159), .ZN(
        n6352) );
  OAI22_X1 U23295 ( .A1(n25162), .A2(n25384), .B1(n9218), .B2(n25159), .ZN(
        n6353) );
  OAI22_X1 U23296 ( .A1(n25162), .A2(n25387), .B1(n9216), .B2(n25159), .ZN(
        n6354) );
  OAI22_X1 U23297 ( .A1(n25163), .A2(n25390), .B1(n9214), .B2(n25159), .ZN(
        n6355) );
  OAI22_X1 U23298 ( .A1(n25163), .A2(n25393), .B1(n9212), .B2(n25159), .ZN(
        n6356) );
  OAI22_X1 U23299 ( .A1(n25163), .A2(n25396), .B1(n9210), .B2(n25159), .ZN(
        n6357) );
  OAI22_X1 U23300 ( .A1(n25163), .A2(n25399), .B1(n9208), .B2(n25159), .ZN(
        n6358) );
  OAI22_X1 U23301 ( .A1(n25163), .A2(n25402), .B1(n9206), .B2(n25159), .ZN(
        n6359) );
  OAI22_X1 U23302 ( .A1(n25164), .A2(n25405), .B1(n9204), .B2(n25159), .ZN(
        n6360) );
  OAI22_X1 U23303 ( .A1(n25164), .A2(n25408), .B1(n9202), .B2(n25159), .ZN(
        n6361) );
  OAI22_X1 U23304 ( .A1(n25164), .A2(n25411), .B1(n9200), .B2(n25159), .ZN(
        n6362) );
  OAI22_X1 U23305 ( .A1(n25164), .A2(n25414), .B1(n9198), .B2(n25159), .ZN(
        n6363) );
  OAI22_X1 U23306 ( .A1(n25335), .A2(n25432), .B1(n99), .B2(n21255), .ZN(n7009) );
  OAI22_X1 U23307 ( .A1(n25336), .A2(n25435), .B1(n98), .B2(n25327), .ZN(n7010) );
  OAI22_X1 U23308 ( .A1(n25336), .A2(n25438), .B1(n97), .B2(n21255), .ZN(n7011) );
  OAI22_X1 U23309 ( .A1(n25336), .A2(n25441), .B1(n96), .B2(n25327), .ZN(n7012) );
  OAI22_X1 U23310 ( .A1(n25336), .A2(n25444), .B1(n95), .B2(n21255), .ZN(n7013) );
  OAI22_X1 U23311 ( .A1(n25336), .A2(n25447), .B1(n94), .B2(n25327), .ZN(n7014) );
  OAI22_X1 U23312 ( .A1(n25337), .A2(n25453), .B1(n92), .B2(n21255), .ZN(n7016) );
  OAI22_X1 U23313 ( .A1(n25337), .A2(n25456), .B1(n91), .B2(n25327), .ZN(n7017) );
  OAI22_X1 U23314 ( .A1(n25337), .A2(n25459), .B1(n90), .B2(n25327), .ZN(n7018) );
  OAI22_X1 U23315 ( .A1(n25338), .A2(n25465), .B1(n88), .B2(n25327), .ZN(n7020) );
  OAI22_X1 U23316 ( .A1(n25338), .A2(n25471), .B1(n86), .B2(n25329), .ZN(n7022) );
  OAI22_X1 U23317 ( .A1(n25096), .A2(n25418), .B1(n7378), .B2(n25090), .ZN(
        n6108) );
  OAI22_X1 U23318 ( .A1(n25097), .A2(n25421), .B1(n7376), .B2(n25091), .ZN(
        n6109) );
  OAI22_X1 U23319 ( .A1(n25097), .A2(n25424), .B1(n7374), .B2(n25089), .ZN(
        n6110) );
  OAI22_X1 U23320 ( .A1(n25097), .A2(n25427), .B1(n7372), .B2(n25090), .ZN(
        n6111) );
  OAI22_X1 U23321 ( .A1(n25097), .A2(n25430), .B1(n7370), .B2(n25091), .ZN(
        n6112) );
  OAI22_X1 U23322 ( .A1(n25097), .A2(n25433), .B1(n7368), .B2(n25089), .ZN(
        n6113) );
  OAI22_X1 U23323 ( .A1(n25098), .A2(n25436), .B1(n7366), .B2(n25090), .ZN(
        n6114) );
  OAI22_X1 U23324 ( .A1(n25098), .A2(n25439), .B1(n7364), .B2(n25091), .ZN(
        n6115) );
  OAI22_X1 U23325 ( .A1(n25098), .A2(n25442), .B1(n7362), .B2(n25089), .ZN(
        n6116) );
  OAI22_X1 U23326 ( .A1(n25098), .A2(n25445), .B1(n7360), .B2(n25090), .ZN(
        n6117) );
  OAI22_X1 U23327 ( .A1(n25098), .A2(n25448), .B1(n7358), .B2(n25091), .ZN(
        n6118) );
  OAI22_X1 U23328 ( .A1(n25099), .A2(n25451), .B1(n7356), .B2(n25089), .ZN(
        n6119) );
  OAI22_X1 U23329 ( .A1(n25099), .A2(n25454), .B1(n7354), .B2(n21278), .ZN(
        n6120) );
  OAI22_X1 U23330 ( .A1(n25099), .A2(n25457), .B1(n7352), .B2(n25089), .ZN(
        n6121) );
  OAI22_X1 U23331 ( .A1(n25099), .A2(n25460), .B1(n7350), .B2(n21278), .ZN(
        n6122) );
  OAI22_X1 U23332 ( .A1(n25099), .A2(n25463), .B1(n7348), .B2(n25089), .ZN(
        n6123) );
  OAI22_X1 U23333 ( .A1(n25100), .A2(n25466), .B1(n7346), .B2(n21278), .ZN(
        n6124) );
  OAI22_X1 U23334 ( .A1(n25100), .A2(n25469), .B1(n7344), .B2(n25089), .ZN(
        n6125) );
  OAI22_X1 U23335 ( .A1(n25100), .A2(n25472), .B1(n7342), .B2(n25090), .ZN(
        n6126) );
  OAI22_X1 U23336 ( .A1(n25100), .A2(n25475), .B1(n7340), .B2(n25091), .ZN(
        n6127) );
  OAI22_X1 U23337 ( .A1(n25100), .A2(n25478), .B1(n7338), .B2(n25089), .ZN(
        n6128) );
  OAI22_X1 U23338 ( .A1(n25101), .A2(n25481), .B1(n7336), .B2(n25089), .ZN(
        n6129) );
  OAI22_X1 U23339 ( .A1(n25101), .A2(n25484), .B1(n7334), .B2(n25090), .ZN(
        n6130) );
  OAI22_X1 U23340 ( .A1(n25101), .A2(n25487), .B1(n7332), .B2(n25091), .ZN(
        n6131) );
  OAI22_X1 U23341 ( .A1(n25101), .A2(n25490), .B1(n7330), .B2(n25089), .ZN(
        n6132) );
  OAI22_X1 U23342 ( .A1(n25101), .A2(n25493), .B1(n7328), .B2(n25089), .ZN(
        n6133) );
  OAI22_X1 U23343 ( .A1(n25102), .A2(n25496), .B1(n7326), .B2(n21278), .ZN(
        n6134) );
  OAI22_X1 U23344 ( .A1(n25102), .A2(n25499), .B1(n7324), .B2(n25089), .ZN(
        n6135) );
  OAI22_X1 U23345 ( .A1(n25102), .A2(n25502), .B1(n7322), .B2(n21278), .ZN(
        n6136) );
  OAI22_X1 U23346 ( .A1(n25102), .A2(n25505), .B1(n7320), .B2(n25089), .ZN(
        n6137) );
  OAI22_X1 U23347 ( .A1(n25102), .A2(n25508), .B1(n7318), .B2(n21278), .ZN(
        n6138) );
  OAI22_X1 U23348 ( .A1(n25103), .A2(n25511), .B1(n7316), .B2(n25089), .ZN(
        n6139) );
  OAI22_X1 U23349 ( .A1(n25103), .A2(n25514), .B1(n7314), .B2(n21278), .ZN(
        n6140) );
  OAI22_X1 U23350 ( .A1(n25103), .A2(n25517), .B1(n7312), .B2(n25089), .ZN(
        n6141) );
  OAI22_X1 U23351 ( .A1(n25103), .A2(n25520), .B1(n7310), .B2(n21278), .ZN(
        n6142) );
  OAI22_X1 U23352 ( .A1(n25103), .A2(n25523), .B1(n7308), .B2(n25089), .ZN(
        n6143) );
  OAI22_X1 U23353 ( .A1(n25104), .A2(n25526), .B1(n7306), .B2(n21278), .ZN(
        n6144) );
  OAI22_X1 U23354 ( .A1(n25104), .A2(n25529), .B1(n7304), .B2(n21278), .ZN(
        n6145) );
  OAI22_X1 U23355 ( .A1(n25104), .A2(n25532), .B1(n7302), .B2(n25089), .ZN(
        n6146) );
  OAI22_X1 U23356 ( .A1(n25104), .A2(n25552), .B1(n7300), .B2(n21278), .ZN(
        n6147) );
  OAI22_X1 U23357 ( .A1(n25266), .A2(n25417), .B1(n17338), .B2(n25260), .ZN(
        n6748) );
  OAI22_X1 U23358 ( .A1(n25267), .A2(n25420), .B1(n17335), .B2(n25261), .ZN(
        n6749) );
  OAI22_X1 U23359 ( .A1(n25267), .A2(n25423), .B1(n17332), .B2(n25259), .ZN(
        n6750) );
  OAI22_X1 U23360 ( .A1(n25267), .A2(n25426), .B1(n17329), .B2(n25260), .ZN(
        n6751) );
  OAI22_X1 U23361 ( .A1(n25267), .A2(n25429), .B1(n17326), .B2(n25261), .ZN(
        n6752) );
  OAI22_X1 U23362 ( .A1(n25267), .A2(n25432), .B1(n17323), .B2(n25259), .ZN(
        n6753) );
  OAI22_X1 U23363 ( .A1(n25268), .A2(n25435), .B1(n17320), .B2(n25260), .ZN(
        n6754) );
  OAI22_X1 U23364 ( .A1(n25268), .A2(n25438), .B1(n17317), .B2(n25261), .ZN(
        n6755) );
  OAI22_X1 U23365 ( .A1(n25268), .A2(n25441), .B1(n17314), .B2(n25259), .ZN(
        n6756) );
  OAI22_X1 U23366 ( .A1(n25268), .A2(n25444), .B1(n17311), .B2(n25260), .ZN(
        n6757) );
  OAI22_X1 U23367 ( .A1(n25268), .A2(n25447), .B1(n17308), .B2(n25261), .ZN(
        n6758) );
  OAI22_X1 U23368 ( .A1(n25269), .A2(n25450), .B1(n17305), .B2(n25259), .ZN(
        n6759) );
  OAI22_X1 U23369 ( .A1(n25269), .A2(n25453), .B1(n17302), .B2(n21263), .ZN(
        n6760) );
  OAI22_X1 U23370 ( .A1(n25269), .A2(n25456), .B1(n17299), .B2(n25259), .ZN(
        n6761) );
  OAI22_X1 U23371 ( .A1(n25269), .A2(n25459), .B1(n17296), .B2(n21263), .ZN(
        n6762) );
  OAI22_X1 U23372 ( .A1(n25269), .A2(n25462), .B1(n17293), .B2(n25259), .ZN(
        n6763) );
  OAI22_X1 U23373 ( .A1(n25270), .A2(n25465), .B1(n17290), .B2(n21263), .ZN(
        n6764) );
  OAI22_X1 U23374 ( .A1(n25270), .A2(n25468), .B1(n17287), .B2(n25259), .ZN(
        n6765) );
  OAI22_X1 U23375 ( .A1(n25270), .A2(n25471), .B1(n17284), .B2(n25260), .ZN(
        n6766) );
  OAI22_X1 U23376 ( .A1(n25270), .A2(n25474), .B1(n17281), .B2(n25261), .ZN(
        n6767) );
  OAI22_X1 U23377 ( .A1(n25270), .A2(n25477), .B1(n17278), .B2(n25259), .ZN(
        n6768) );
  OAI22_X1 U23378 ( .A1(n25271), .A2(n25480), .B1(n17275), .B2(n25259), .ZN(
        n6769) );
  OAI22_X1 U23379 ( .A1(n25271), .A2(n25483), .B1(n17272), .B2(n25260), .ZN(
        n6770) );
  OAI22_X1 U23380 ( .A1(n25271), .A2(n25486), .B1(n17269), .B2(n25261), .ZN(
        n6771) );
  OAI22_X1 U23381 ( .A1(n25271), .A2(n25489), .B1(n17266), .B2(n25259), .ZN(
        n6772) );
  OAI22_X1 U23382 ( .A1(n25271), .A2(n25492), .B1(n17263), .B2(n25259), .ZN(
        n6773) );
  OAI22_X1 U23383 ( .A1(n25272), .A2(n25495), .B1(n17260), .B2(n21263), .ZN(
        n6774) );
  OAI22_X1 U23384 ( .A1(n25272), .A2(n25498), .B1(n17257), .B2(n25259), .ZN(
        n6775) );
  OAI22_X1 U23385 ( .A1(n25272), .A2(n25501), .B1(n17254), .B2(n21263), .ZN(
        n6776) );
  OAI22_X1 U23386 ( .A1(n25272), .A2(n25504), .B1(n17251), .B2(n25259), .ZN(
        n6777) );
  OAI22_X1 U23387 ( .A1(n25272), .A2(n25507), .B1(n17248), .B2(n21263), .ZN(
        n6778) );
  OAI22_X1 U23388 ( .A1(n25273), .A2(n25510), .B1(n17245), .B2(n25259), .ZN(
        n6779) );
  OAI22_X1 U23389 ( .A1(n25273), .A2(n25513), .B1(n17242), .B2(n21263), .ZN(
        n6780) );
  OAI22_X1 U23390 ( .A1(n25273), .A2(n25516), .B1(n17239), .B2(n25259), .ZN(
        n6781) );
  OAI22_X1 U23391 ( .A1(n25273), .A2(n25519), .B1(n17236), .B2(n21263), .ZN(
        n6782) );
  OAI22_X1 U23392 ( .A1(n25273), .A2(n25522), .B1(n17233), .B2(n25259), .ZN(
        n6783) );
  OAI22_X1 U23393 ( .A1(n25181), .A2(n25417), .B1(n7506), .B2(n25175), .ZN(
        n6428) );
  OAI22_X1 U23394 ( .A1(n25182), .A2(n25420), .B1(n7504), .B2(n25176), .ZN(
        n6429) );
  OAI22_X1 U23395 ( .A1(n25182), .A2(n25423), .B1(n7502), .B2(n25174), .ZN(
        n6430) );
  OAI22_X1 U23396 ( .A1(n25182), .A2(n25426), .B1(n7500), .B2(n25175), .ZN(
        n6431) );
  OAI22_X1 U23397 ( .A1(n25182), .A2(n25429), .B1(n7498), .B2(n25176), .ZN(
        n6432) );
  OAI22_X1 U23398 ( .A1(n25182), .A2(n25432), .B1(n7496), .B2(n25174), .ZN(
        n6433) );
  OAI22_X1 U23399 ( .A1(n25183), .A2(n25435), .B1(n7494), .B2(n25175), .ZN(
        n6434) );
  OAI22_X1 U23400 ( .A1(n25183), .A2(n25438), .B1(n7492), .B2(n25176), .ZN(
        n6435) );
  OAI22_X1 U23401 ( .A1(n25183), .A2(n25441), .B1(n7490), .B2(n25174), .ZN(
        n6436) );
  OAI22_X1 U23402 ( .A1(n25183), .A2(n25444), .B1(n7488), .B2(n25175), .ZN(
        n6437) );
  OAI22_X1 U23403 ( .A1(n25183), .A2(n25447), .B1(n7486), .B2(n25176), .ZN(
        n6438) );
  OAI22_X1 U23404 ( .A1(n25184), .A2(n25450), .B1(n7484), .B2(n25174), .ZN(
        n6439) );
  OAI22_X1 U23405 ( .A1(n25184), .A2(n25453), .B1(n7482), .B2(n21273), .ZN(
        n6440) );
  OAI22_X1 U23406 ( .A1(n25184), .A2(n25456), .B1(n7480), .B2(n25174), .ZN(
        n6441) );
  OAI22_X1 U23407 ( .A1(n25184), .A2(n25459), .B1(n7478), .B2(n21273), .ZN(
        n6442) );
  OAI22_X1 U23408 ( .A1(n25184), .A2(n25462), .B1(n7476), .B2(n25174), .ZN(
        n6443) );
  OAI22_X1 U23409 ( .A1(n25185), .A2(n25465), .B1(n7474), .B2(n21273), .ZN(
        n6444) );
  OAI22_X1 U23410 ( .A1(n25185), .A2(n25468), .B1(n7472), .B2(n25174), .ZN(
        n6445) );
  OAI22_X1 U23411 ( .A1(n25185), .A2(n25471), .B1(n7470), .B2(n25175), .ZN(
        n6446) );
  OAI22_X1 U23412 ( .A1(n25185), .A2(n25474), .B1(n7468), .B2(n25176), .ZN(
        n6447) );
  OAI22_X1 U23413 ( .A1(n25185), .A2(n25477), .B1(n7466), .B2(n25174), .ZN(
        n6448) );
  OAI22_X1 U23414 ( .A1(n25186), .A2(n25480), .B1(n7464), .B2(n25174), .ZN(
        n6449) );
  OAI22_X1 U23415 ( .A1(n25186), .A2(n25483), .B1(n7462), .B2(n25175), .ZN(
        n6450) );
  OAI22_X1 U23416 ( .A1(n25186), .A2(n25486), .B1(n7460), .B2(n25176), .ZN(
        n6451) );
  OAI22_X1 U23417 ( .A1(n25186), .A2(n25489), .B1(n7458), .B2(n25174), .ZN(
        n6452) );
  OAI22_X1 U23418 ( .A1(n25186), .A2(n25492), .B1(n7456), .B2(n25174), .ZN(
        n6453) );
  OAI22_X1 U23419 ( .A1(n25187), .A2(n25495), .B1(n7454), .B2(n21273), .ZN(
        n6454) );
  OAI22_X1 U23420 ( .A1(n25187), .A2(n25498), .B1(n7452), .B2(n25174), .ZN(
        n6455) );
  OAI22_X1 U23421 ( .A1(n25187), .A2(n25501), .B1(n7450), .B2(n21273), .ZN(
        n6456) );
  OAI22_X1 U23422 ( .A1(n25187), .A2(n25504), .B1(n7448), .B2(n25174), .ZN(
        n6457) );
  OAI22_X1 U23423 ( .A1(n25187), .A2(n25507), .B1(n7446), .B2(n21273), .ZN(
        n6458) );
  OAI22_X1 U23424 ( .A1(n25188), .A2(n25510), .B1(n7444), .B2(n25174), .ZN(
        n6459) );
  OAI22_X1 U23425 ( .A1(n25188), .A2(n25513), .B1(n7442), .B2(n21273), .ZN(
        n6460) );
  OAI22_X1 U23426 ( .A1(n25188), .A2(n25516), .B1(n7440), .B2(n25174), .ZN(
        n6461) );
  OAI22_X1 U23427 ( .A1(n25188), .A2(n25519), .B1(n7438), .B2(n21273), .ZN(
        n6462) );
  OAI22_X1 U23428 ( .A1(n25188), .A2(n25522), .B1(n7436), .B2(n25174), .ZN(
        n6463) );
  OAI22_X1 U23429 ( .A1(n25045), .A2(n25418), .B1(n8813), .B2(n25039), .ZN(
        n5916) );
  OAI22_X1 U23430 ( .A1(n25046), .A2(n25421), .B1(n8811), .B2(n25040), .ZN(
        n5917) );
  OAI22_X1 U23431 ( .A1(n25046), .A2(n25424), .B1(n8809), .B2(n25038), .ZN(
        n5918) );
  OAI22_X1 U23432 ( .A1(n25046), .A2(n25427), .B1(n8807), .B2(n25039), .ZN(
        n5919) );
  OAI22_X1 U23433 ( .A1(n25046), .A2(n25430), .B1(n8805), .B2(n25040), .ZN(
        n5920) );
  OAI22_X1 U23434 ( .A1(n25046), .A2(n25433), .B1(n8803), .B2(n25038), .ZN(
        n5921) );
  OAI22_X1 U23435 ( .A1(n25047), .A2(n25436), .B1(n8801), .B2(n25039), .ZN(
        n5922) );
  OAI22_X1 U23436 ( .A1(n25047), .A2(n25439), .B1(n8799), .B2(n25040), .ZN(
        n5923) );
  OAI22_X1 U23437 ( .A1(n25047), .A2(n25442), .B1(n8797), .B2(n25038), .ZN(
        n5924) );
  OAI22_X1 U23438 ( .A1(n25047), .A2(n25445), .B1(n8795), .B2(n25039), .ZN(
        n5925) );
  OAI22_X1 U23439 ( .A1(n25047), .A2(n25448), .B1(n8793), .B2(n25040), .ZN(
        n5926) );
  OAI22_X1 U23440 ( .A1(n25048), .A2(n25451), .B1(n8791), .B2(n25038), .ZN(
        n5927) );
  OAI22_X1 U23441 ( .A1(n25048), .A2(n25454), .B1(n8789), .B2(n21282), .ZN(
        n5928) );
  OAI22_X1 U23442 ( .A1(n25048), .A2(n25457), .B1(n8787), .B2(n25038), .ZN(
        n5929) );
  OAI22_X1 U23443 ( .A1(n25048), .A2(n25460), .B1(n8785), .B2(n21282), .ZN(
        n5930) );
  OAI22_X1 U23444 ( .A1(n25048), .A2(n25463), .B1(n8783), .B2(n25038), .ZN(
        n5931) );
  OAI22_X1 U23445 ( .A1(n25049), .A2(n25466), .B1(n8781), .B2(n21282), .ZN(
        n5932) );
  OAI22_X1 U23446 ( .A1(n25049), .A2(n25469), .B1(n8779), .B2(n25038), .ZN(
        n5933) );
  OAI22_X1 U23447 ( .A1(n25049), .A2(n25472), .B1(n8777), .B2(n25039), .ZN(
        n5934) );
  OAI22_X1 U23448 ( .A1(n25049), .A2(n25475), .B1(n8775), .B2(n25040), .ZN(
        n5935) );
  OAI22_X1 U23449 ( .A1(n25049), .A2(n25478), .B1(n8773), .B2(n25038), .ZN(
        n5936) );
  OAI22_X1 U23450 ( .A1(n25050), .A2(n25481), .B1(n8771), .B2(n25038), .ZN(
        n5937) );
  OAI22_X1 U23451 ( .A1(n25050), .A2(n25484), .B1(n8769), .B2(n25039), .ZN(
        n5938) );
  OAI22_X1 U23452 ( .A1(n25050), .A2(n25487), .B1(n8767), .B2(n25040), .ZN(
        n5939) );
  OAI22_X1 U23453 ( .A1(n25050), .A2(n25490), .B1(n8765), .B2(n25038), .ZN(
        n5940) );
  OAI22_X1 U23454 ( .A1(n25050), .A2(n25493), .B1(n8763), .B2(n25038), .ZN(
        n5941) );
  OAI22_X1 U23455 ( .A1(n25051), .A2(n25496), .B1(n8761), .B2(n21282), .ZN(
        n5942) );
  OAI22_X1 U23456 ( .A1(n25051), .A2(n25499), .B1(n8759), .B2(n25038), .ZN(
        n5943) );
  OAI22_X1 U23457 ( .A1(n25051), .A2(n25502), .B1(n8757), .B2(n21282), .ZN(
        n5944) );
  OAI22_X1 U23458 ( .A1(n25051), .A2(n25505), .B1(n8755), .B2(n25038), .ZN(
        n5945) );
  OAI22_X1 U23459 ( .A1(n25051), .A2(n25508), .B1(n8753), .B2(n21282), .ZN(
        n5946) );
  OAI22_X1 U23460 ( .A1(n25052), .A2(n25511), .B1(n8751), .B2(n25038), .ZN(
        n5947) );
  OAI22_X1 U23461 ( .A1(n25052), .A2(n25514), .B1(n8749), .B2(n21282), .ZN(
        n5948) );
  OAI22_X1 U23462 ( .A1(n25052), .A2(n25517), .B1(n8747), .B2(n25038), .ZN(
        n5949) );
  OAI22_X1 U23463 ( .A1(n25052), .A2(n25520), .B1(n8745), .B2(n21282), .ZN(
        n5950) );
  OAI22_X1 U23464 ( .A1(n25052), .A2(n25523), .B1(n8743), .B2(n25038), .ZN(
        n5951) );
  OAI22_X1 U23465 ( .A1(n25028), .A2(n25418), .B1(n8941), .B2(n25022), .ZN(
        n5852) );
  OAI22_X1 U23466 ( .A1(n25029), .A2(n25421), .B1(n8939), .B2(n25023), .ZN(
        n5853) );
  OAI22_X1 U23467 ( .A1(n25029), .A2(n25424), .B1(n8937), .B2(n25021), .ZN(
        n5854) );
  OAI22_X1 U23468 ( .A1(n25029), .A2(n25427), .B1(n8935), .B2(n25022), .ZN(
        n5855) );
  OAI22_X1 U23469 ( .A1(n25029), .A2(n25430), .B1(n8933), .B2(n25023), .ZN(
        n5856) );
  OAI22_X1 U23470 ( .A1(n25029), .A2(n25433), .B1(n8931), .B2(n25021), .ZN(
        n5857) );
  OAI22_X1 U23471 ( .A1(n25030), .A2(n25436), .B1(n8929), .B2(n25022), .ZN(
        n5858) );
  OAI22_X1 U23472 ( .A1(n25030), .A2(n25439), .B1(n8927), .B2(n25023), .ZN(
        n5859) );
  OAI22_X1 U23473 ( .A1(n25030), .A2(n25442), .B1(n8925), .B2(n25021), .ZN(
        n5860) );
  OAI22_X1 U23474 ( .A1(n25030), .A2(n25445), .B1(n8923), .B2(n25022), .ZN(
        n5861) );
  OAI22_X1 U23475 ( .A1(n25030), .A2(n25448), .B1(n8921), .B2(n25023), .ZN(
        n5862) );
  OAI22_X1 U23476 ( .A1(n25031), .A2(n25451), .B1(n8919), .B2(n25021), .ZN(
        n5863) );
  OAI22_X1 U23477 ( .A1(n25031), .A2(n25454), .B1(n8917), .B2(n21283), .ZN(
        n5864) );
  OAI22_X1 U23478 ( .A1(n25031), .A2(n25457), .B1(n8915), .B2(n25021), .ZN(
        n5865) );
  OAI22_X1 U23479 ( .A1(n25031), .A2(n25460), .B1(n8913), .B2(n21283), .ZN(
        n5866) );
  OAI22_X1 U23480 ( .A1(n25031), .A2(n25463), .B1(n8911), .B2(n25021), .ZN(
        n5867) );
  OAI22_X1 U23481 ( .A1(n25032), .A2(n25466), .B1(n8909), .B2(n21283), .ZN(
        n5868) );
  OAI22_X1 U23482 ( .A1(n25032), .A2(n25469), .B1(n8907), .B2(n25021), .ZN(
        n5869) );
  OAI22_X1 U23483 ( .A1(n25032), .A2(n25472), .B1(n8905), .B2(n25022), .ZN(
        n5870) );
  OAI22_X1 U23484 ( .A1(n25032), .A2(n25475), .B1(n8903), .B2(n25023), .ZN(
        n5871) );
  OAI22_X1 U23485 ( .A1(n25032), .A2(n25478), .B1(n8901), .B2(n25021), .ZN(
        n5872) );
  OAI22_X1 U23486 ( .A1(n25033), .A2(n25481), .B1(n8899), .B2(n25021), .ZN(
        n5873) );
  OAI22_X1 U23487 ( .A1(n25033), .A2(n25484), .B1(n8897), .B2(n25022), .ZN(
        n5874) );
  OAI22_X1 U23488 ( .A1(n25033), .A2(n25487), .B1(n8895), .B2(n25023), .ZN(
        n5875) );
  OAI22_X1 U23489 ( .A1(n25033), .A2(n25490), .B1(n8893), .B2(n25021), .ZN(
        n5876) );
  OAI22_X1 U23490 ( .A1(n25033), .A2(n25493), .B1(n8891), .B2(n25021), .ZN(
        n5877) );
  OAI22_X1 U23491 ( .A1(n25034), .A2(n25496), .B1(n8889), .B2(n21283), .ZN(
        n5878) );
  OAI22_X1 U23492 ( .A1(n25034), .A2(n25499), .B1(n8887), .B2(n25021), .ZN(
        n5879) );
  OAI22_X1 U23493 ( .A1(n25034), .A2(n25502), .B1(n8885), .B2(n21283), .ZN(
        n5880) );
  OAI22_X1 U23494 ( .A1(n25034), .A2(n25505), .B1(n8883), .B2(n25021), .ZN(
        n5881) );
  OAI22_X1 U23495 ( .A1(n25034), .A2(n25508), .B1(n8881), .B2(n21283), .ZN(
        n5882) );
  OAI22_X1 U23496 ( .A1(n25035), .A2(n25511), .B1(n8879), .B2(n25021), .ZN(
        n5883) );
  OAI22_X1 U23497 ( .A1(n25035), .A2(n25514), .B1(n8877), .B2(n21283), .ZN(
        n5884) );
  OAI22_X1 U23498 ( .A1(n25035), .A2(n25517), .B1(n8875), .B2(n25021), .ZN(
        n5885) );
  OAI22_X1 U23499 ( .A1(n25035), .A2(n25520), .B1(n8873), .B2(n21283), .ZN(
        n5886) );
  OAI22_X1 U23500 ( .A1(n25035), .A2(n25523), .B1(n8871), .B2(n25021), .ZN(
        n5887) );
  OAI22_X1 U23501 ( .A1(n24858), .A2(n25419), .B1(n8940), .B2(n24852), .ZN(
        n5212) );
  OAI22_X1 U23502 ( .A1(n24859), .A2(n25422), .B1(n8938), .B2(n24853), .ZN(
        n5213) );
  OAI22_X1 U23503 ( .A1(n24859), .A2(n25425), .B1(n8936), .B2(n24851), .ZN(
        n5214) );
  OAI22_X1 U23504 ( .A1(n24859), .A2(n25428), .B1(n8934), .B2(n24852), .ZN(
        n5215) );
  OAI22_X1 U23505 ( .A1(n24859), .A2(n25431), .B1(n8932), .B2(n24853), .ZN(
        n5216) );
  OAI22_X1 U23506 ( .A1(n24859), .A2(n25434), .B1(n8930), .B2(n24851), .ZN(
        n5217) );
  OAI22_X1 U23507 ( .A1(n24860), .A2(n25437), .B1(n8928), .B2(n24852), .ZN(
        n5218) );
  OAI22_X1 U23508 ( .A1(n24860), .A2(n25440), .B1(n8926), .B2(n24853), .ZN(
        n5219) );
  OAI22_X1 U23509 ( .A1(n24860), .A2(n25443), .B1(n8924), .B2(n24851), .ZN(
        n5220) );
  OAI22_X1 U23510 ( .A1(n24860), .A2(n25446), .B1(n8922), .B2(n24852), .ZN(
        n5221) );
  OAI22_X1 U23511 ( .A1(n24860), .A2(n25449), .B1(n8920), .B2(n24853), .ZN(
        n5222) );
  OAI22_X1 U23512 ( .A1(n24861), .A2(n25452), .B1(n8918), .B2(n24851), .ZN(
        n5223) );
  OAI22_X1 U23513 ( .A1(n24861), .A2(n25455), .B1(n8916), .B2(n21294), .ZN(
        n5224) );
  OAI22_X1 U23514 ( .A1(n24861), .A2(n25458), .B1(n8914), .B2(n24851), .ZN(
        n5225) );
  OAI22_X1 U23515 ( .A1(n24861), .A2(n25461), .B1(n8912), .B2(n21294), .ZN(
        n5226) );
  OAI22_X1 U23516 ( .A1(n24861), .A2(n25464), .B1(n8910), .B2(n24851), .ZN(
        n5227) );
  OAI22_X1 U23517 ( .A1(n24862), .A2(n25467), .B1(n8908), .B2(n21294), .ZN(
        n5228) );
  OAI22_X1 U23518 ( .A1(n24862), .A2(n25470), .B1(n8906), .B2(n24851), .ZN(
        n5229) );
  OAI22_X1 U23519 ( .A1(n24862), .A2(n25473), .B1(n8904), .B2(n24852), .ZN(
        n5230) );
  OAI22_X1 U23520 ( .A1(n24862), .A2(n25476), .B1(n8902), .B2(n24853), .ZN(
        n5231) );
  OAI22_X1 U23521 ( .A1(n24862), .A2(n25479), .B1(n8900), .B2(n24851), .ZN(
        n5232) );
  OAI22_X1 U23522 ( .A1(n24863), .A2(n25482), .B1(n8898), .B2(n24851), .ZN(
        n5233) );
  OAI22_X1 U23523 ( .A1(n24863), .A2(n25485), .B1(n8896), .B2(n24852), .ZN(
        n5234) );
  OAI22_X1 U23524 ( .A1(n24863), .A2(n25488), .B1(n8894), .B2(n24853), .ZN(
        n5235) );
  OAI22_X1 U23525 ( .A1(n24863), .A2(n25491), .B1(n8892), .B2(n24851), .ZN(
        n5236) );
  OAI22_X1 U23526 ( .A1(n24863), .A2(n25494), .B1(n8890), .B2(n24851), .ZN(
        n5237) );
  OAI22_X1 U23527 ( .A1(n24864), .A2(n25497), .B1(n8888), .B2(n21294), .ZN(
        n5238) );
  OAI22_X1 U23528 ( .A1(n24864), .A2(n25500), .B1(n8886), .B2(n24851), .ZN(
        n5239) );
  OAI22_X1 U23529 ( .A1(n24864), .A2(n25503), .B1(n8884), .B2(n21294), .ZN(
        n5240) );
  OAI22_X1 U23530 ( .A1(n24864), .A2(n25506), .B1(n8882), .B2(n24851), .ZN(
        n5241) );
  OAI22_X1 U23531 ( .A1(n24864), .A2(n25509), .B1(n8880), .B2(n21294), .ZN(
        n5242) );
  OAI22_X1 U23532 ( .A1(n24865), .A2(n25512), .B1(n8878), .B2(n24851), .ZN(
        n5243) );
  OAI22_X1 U23533 ( .A1(n24865), .A2(n25515), .B1(n8876), .B2(n21294), .ZN(
        n5244) );
  OAI22_X1 U23534 ( .A1(n24865), .A2(n25518), .B1(n8874), .B2(n24851), .ZN(
        n5245) );
  OAI22_X1 U23535 ( .A1(n24865), .A2(n25521), .B1(n8872), .B2(n21294), .ZN(
        n5246) );
  OAI22_X1 U23536 ( .A1(n24865), .A2(n25524), .B1(n8870), .B2(n24851), .ZN(
        n5247) );
  OAI22_X1 U23537 ( .A1(n24926), .A2(n25419), .B1(n7379), .B2(n24920), .ZN(
        n5468) );
  OAI22_X1 U23538 ( .A1(n24927), .A2(n25422), .B1(n7377), .B2(n24921), .ZN(
        n5469) );
  OAI22_X1 U23539 ( .A1(n24927), .A2(n25425), .B1(n7375), .B2(n24919), .ZN(
        n5470) );
  OAI22_X1 U23540 ( .A1(n24927), .A2(n25428), .B1(n7373), .B2(n24920), .ZN(
        n5471) );
  OAI22_X1 U23541 ( .A1(n24927), .A2(n25431), .B1(n7371), .B2(n24921), .ZN(
        n5472) );
  OAI22_X1 U23542 ( .A1(n24927), .A2(n25434), .B1(n7369), .B2(n24919), .ZN(
        n5473) );
  OAI22_X1 U23543 ( .A1(n24928), .A2(n25437), .B1(n7367), .B2(n24920), .ZN(
        n5474) );
  OAI22_X1 U23544 ( .A1(n24928), .A2(n25440), .B1(n7365), .B2(n24921), .ZN(
        n5475) );
  OAI22_X1 U23545 ( .A1(n24928), .A2(n25443), .B1(n7363), .B2(n24919), .ZN(
        n5476) );
  OAI22_X1 U23546 ( .A1(n24928), .A2(n25446), .B1(n7361), .B2(n24920), .ZN(
        n5477) );
  OAI22_X1 U23547 ( .A1(n24928), .A2(n25449), .B1(n7359), .B2(n24921), .ZN(
        n5478) );
  OAI22_X1 U23548 ( .A1(n24929), .A2(n25452), .B1(n7357), .B2(n24919), .ZN(
        n5479) );
  OAI22_X1 U23549 ( .A1(n24929), .A2(n25455), .B1(n7355), .B2(n21290), .ZN(
        n5480) );
  OAI22_X1 U23550 ( .A1(n24929), .A2(n25458), .B1(n7353), .B2(n24919), .ZN(
        n5481) );
  OAI22_X1 U23551 ( .A1(n24929), .A2(n25461), .B1(n7351), .B2(n21290), .ZN(
        n5482) );
  OAI22_X1 U23552 ( .A1(n24929), .A2(n25464), .B1(n7349), .B2(n24919), .ZN(
        n5483) );
  OAI22_X1 U23553 ( .A1(n24930), .A2(n25467), .B1(n7347), .B2(n21290), .ZN(
        n5484) );
  OAI22_X1 U23554 ( .A1(n24930), .A2(n25470), .B1(n7345), .B2(n24919), .ZN(
        n5485) );
  OAI22_X1 U23555 ( .A1(n24930), .A2(n25473), .B1(n7343), .B2(n24920), .ZN(
        n5486) );
  OAI22_X1 U23556 ( .A1(n24930), .A2(n25476), .B1(n7341), .B2(n24921), .ZN(
        n5487) );
  OAI22_X1 U23557 ( .A1(n24930), .A2(n25479), .B1(n7339), .B2(n24919), .ZN(
        n5488) );
  OAI22_X1 U23558 ( .A1(n24931), .A2(n25482), .B1(n7337), .B2(n24919), .ZN(
        n5489) );
  OAI22_X1 U23559 ( .A1(n24931), .A2(n25485), .B1(n7335), .B2(n24920), .ZN(
        n5490) );
  OAI22_X1 U23560 ( .A1(n24931), .A2(n25488), .B1(n7333), .B2(n24921), .ZN(
        n5491) );
  OAI22_X1 U23561 ( .A1(n24931), .A2(n25491), .B1(n7331), .B2(n24919), .ZN(
        n5492) );
  OAI22_X1 U23562 ( .A1(n24931), .A2(n25494), .B1(n7329), .B2(n24919), .ZN(
        n5493) );
  OAI22_X1 U23563 ( .A1(n24932), .A2(n25497), .B1(n7327), .B2(n21290), .ZN(
        n5494) );
  OAI22_X1 U23564 ( .A1(n24932), .A2(n25500), .B1(n7325), .B2(n24919), .ZN(
        n5495) );
  OAI22_X1 U23565 ( .A1(n24932), .A2(n25503), .B1(n7323), .B2(n21290), .ZN(
        n5496) );
  OAI22_X1 U23566 ( .A1(n24932), .A2(n25506), .B1(n7321), .B2(n24919), .ZN(
        n5497) );
  OAI22_X1 U23567 ( .A1(n24932), .A2(n25509), .B1(n7319), .B2(n21290), .ZN(
        n5498) );
  OAI22_X1 U23568 ( .A1(n24933), .A2(n25512), .B1(n7317), .B2(n24919), .ZN(
        n5499) );
  OAI22_X1 U23569 ( .A1(n24933), .A2(n25515), .B1(n7315), .B2(n21290), .ZN(
        n5500) );
  OAI22_X1 U23570 ( .A1(n24933), .A2(n25518), .B1(n7313), .B2(n24919), .ZN(
        n5501) );
  OAI22_X1 U23571 ( .A1(n24933), .A2(n25521), .B1(n7311), .B2(n21290), .ZN(
        n5502) );
  OAI22_X1 U23572 ( .A1(n24933), .A2(n25524), .B1(n7309), .B2(n24919), .ZN(
        n5503) );
  OAI22_X1 U23573 ( .A1(n24960), .A2(n25418), .B1(n9197), .B2(n24954), .ZN(
        n5596) );
  OAI22_X1 U23574 ( .A1(n24961), .A2(n25421), .B1(n9195), .B2(n24955), .ZN(
        n5597) );
  OAI22_X1 U23575 ( .A1(n24961), .A2(n25424), .B1(n9193), .B2(n24953), .ZN(
        n5598) );
  OAI22_X1 U23576 ( .A1(n24961), .A2(n25427), .B1(n9191), .B2(n24954), .ZN(
        n5599) );
  OAI22_X1 U23577 ( .A1(n24961), .A2(n25430), .B1(n9189), .B2(n24955), .ZN(
        n5600) );
  OAI22_X1 U23578 ( .A1(n24961), .A2(n25433), .B1(n9187), .B2(n24953), .ZN(
        n5601) );
  OAI22_X1 U23579 ( .A1(n24962), .A2(n25436), .B1(n9185), .B2(n24954), .ZN(
        n5602) );
  OAI22_X1 U23580 ( .A1(n24962), .A2(n25439), .B1(n9183), .B2(n24955), .ZN(
        n5603) );
  OAI22_X1 U23581 ( .A1(n24962), .A2(n25442), .B1(n9181), .B2(n24953), .ZN(
        n5604) );
  OAI22_X1 U23582 ( .A1(n24962), .A2(n25445), .B1(n9179), .B2(n24954), .ZN(
        n5605) );
  OAI22_X1 U23583 ( .A1(n24962), .A2(n25448), .B1(n9177), .B2(n24955), .ZN(
        n5606) );
  OAI22_X1 U23584 ( .A1(n24963), .A2(n25451), .B1(n9175), .B2(n24953), .ZN(
        n5607) );
  OAI22_X1 U23585 ( .A1(n24963), .A2(n25454), .B1(n9173), .B2(n21287), .ZN(
        n5608) );
  OAI22_X1 U23586 ( .A1(n24963), .A2(n25457), .B1(n9171), .B2(n24953), .ZN(
        n5609) );
  OAI22_X1 U23587 ( .A1(n24963), .A2(n25460), .B1(n9169), .B2(n21287), .ZN(
        n5610) );
  OAI22_X1 U23588 ( .A1(n24963), .A2(n25463), .B1(n9167), .B2(n24953), .ZN(
        n5611) );
  OAI22_X1 U23589 ( .A1(n24964), .A2(n25466), .B1(n9165), .B2(n21287), .ZN(
        n5612) );
  OAI22_X1 U23590 ( .A1(n24964), .A2(n25469), .B1(n9163), .B2(n24953), .ZN(
        n5613) );
  OAI22_X1 U23591 ( .A1(n24964), .A2(n25472), .B1(n9161), .B2(n24954), .ZN(
        n5614) );
  OAI22_X1 U23592 ( .A1(n24964), .A2(n25475), .B1(n9159), .B2(n24955), .ZN(
        n5615) );
  OAI22_X1 U23593 ( .A1(n24964), .A2(n25478), .B1(n9157), .B2(n24953), .ZN(
        n5616) );
  OAI22_X1 U23594 ( .A1(n24965), .A2(n25481), .B1(n9155), .B2(n24953), .ZN(
        n5617) );
  OAI22_X1 U23595 ( .A1(n24965), .A2(n25484), .B1(n9153), .B2(n24954), .ZN(
        n5618) );
  OAI22_X1 U23596 ( .A1(n24965), .A2(n25487), .B1(n9151), .B2(n24955), .ZN(
        n5619) );
  OAI22_X1 U23597 ( .A1(n24965), .A2(n25490), .B1(n9149), .B2(n24953), .ZN(
        n5620) );
  OAI22_X1 U23598 ( .A1(n24965), .A2(n25493), .B1(n9147), .B2(n24953), .ZN(
        n5621) );
  OAI22_X1 U23599 ( .A1(n24966), .A2(n25496), .B1(n9145), .B2(n21287), .ZN(
        n5622) );
  OAI22_X1 U23600 ( .A1(n24966), .A2(n25499), .B1(n9143), .B2(n24953), .ZN(
        n5623) );
  OAI22_X1 U23601 ( .A1(n24966), .A2(n25502), .B1(n9141), .B2(n21287), .ZN(
        n5624) );
  OAI22_X1 U23602 ( .A1(n24966), .A2(n25505), .B1(n9139), .B2(n24953), .ZN(
        n5625) );
  OAI22_X1 U23603 ( .A1(n24966), .A2(n25508), .B1(n9137), .B2(n21287), .ZN(
        n5626) );
  OAI22_X1 U23604 ( .A1(n24967), .A2(n25511), .B1(n9135), .B2(n24953), .ZN(
        n5627) );
  OAI22_X1 U23605 ( .A1(n24967), .A2(n25514), .B1(n9133), .B2(n21287), .ZN(
        n5628) );
  OAI22_X1 U23606 ( .A1(n24967), .A2(n25517), .B1(n9131), .B2(n24953), .ZN(
        n5629) );
  OAI22_X1 U23607 ( .A1(n24967), .A2(n25520), .B1(n9129), .B2(n21287), .ZN(
        n5630) );
  OAI22_X1 U23608 ( .A1(n24967), .A2(n25523), .B1(n9127), .B2(n24953), .ZN(
        n5631) );
  OAI22_X1 U23609 ( .A1(n24977), .A2(n25418), .B1(n7507), .B2(n24971), .ZN(
        n5660) );
  OAI22_X1 U23610 ( .A1(n24978), .A2(n25421), .B1(n7505), .B2(n24972), .ZN(
        n5661) );
  OAI22_X1 U23611 ( .A1(n24978), .A2(n25424), .B1(n7503), .B2(n24970), .ZN(
        n5662) );
  OAI22_X1 U23612 ( .A1(n24978), .A2(n25427), .B1(n7501), .B2(n24971), .ZN(
        n5663) );
  OAI22_X1 U23613 ( .A1(n24978), .A2(n25430), .B1(n7499), .B2(n24972), .ZN(
        n5664) );
  OAI22_X1 U23614 ( .A1(n24978), .A2(n25433), .B1(n7497), .B2(n24970), .ZN(
        n5665) );
  OAI22_X1 U23615 ( .A1(n24979), .A2(n25436), .B1(n7495), .B2(n24971), .ZN(
        n5666) );
  OAI22_X1 U23616 ( .A1(n24979), .A2(n25439), .B1(n7493), .B2(n24972), .ZN(
        n5667) );
  OAI22_X1 U23617 ( .A1(n24979), .A2(n25442), .B1(n7491), .B2(n24970), .ZN(
        n5668) );
  OAI22_X1 U23618 ( .A1(n24979), .A2(n25445), .B1(n7489), .B2(n24971), .ZN(
        n5669) );
  OAI22_X1 U23619 ( .A1(n24979), .A2(n25448), .B1(n7487), .B2(n24972), .ZN(
        n5670) );
  OAI22_X1 U23620 ( .A1(n24980), .A2(n25451), .B1(n7485), .B2(n24970), .ZN(
        n5671) );
  OAI22_X1 U23621 ( .A1(n24980), .A2(n25454), .B1(n7483), .B2(n21286), .ZN(
        n5672) );
  OAI22_X1 U23622 ( .A1(n24980), .A2(n25457), .B1(n7481), .B2(n24970), .ZN(
        n5673) );
  OAI22_X1 U23623 ( .A1(n24980), .A2(n25460), .B1(n7479), .B2(n21286), .ZN(
        n5674) );
  OAI22_X1 U23624 ( .A1(n24980), .A2(n25463), .B1(n7477), .B2(n24970), .ZN(
        n5675) );
  OAI22_X1 U23625 ( .A1(n24981), .A2(n25466), .B1(n7475), .B2(n21286), .ZN(
        n5676) );
  OAI22_X1 U23626 ( .A1(n24981), .A2(n25469), .B1(n7473), .B2(n24970), .ZN(
        n5677) );
  OAI22_X1 U23627 ( .A1(n24981), .A2(n25472), .B1(n7471), .B2(n24971), .ZN(
        n5678) );
  OAI22_X1 U23628 ( .A1(n24981), .A2(n25475), .B1(n7469), .B2(n24972), .ZN(
        n5679) );
  OAI22_X1 U23629 ( .A1(n24981), .A2(n25478), .B1(n7467), .B2(n24970), .ZN(
        n5680) );
  OAI22_X1 U23630 ( .A1(n24982), .A2(n25481), .B1(n7465), .B2(n24970), .ZN(
        n5681) );
  OAI22_X1 U23631 ( .A1(n24982), .A2(n25484), .B1(n7463), .B2(n24971), .ZN(
        n5682) );
  OAI22_X1 U23632 ( .A1(n24982), .A2(n25487), .B1(n7461), .B2(n24972), .ZN(
        n5683) );
  OAI22_X1 U23633 ( .A1(n24982), .A2(n25490), .B1(n7459), .B2(n24970), .ZN(
        n5684) );
  OAI22_X1 U23634 ( .A1(n24982), .A2(n25493), .B1(n7457), .B2(n24970), .ZN(
        n5685) );
  OAI22_X1 U23635 ( .A1(n24983), .A2(n25496), .B1(n7455), .B2(n21286), .ZN(
        n5686) );
  OAI22_X1 U23636 ( .A1(n24983), .A2(n25499), .B1(n7453), .B2(n24970), .ZN(
        n5687) );
  OAI22_X1 U23637 ( .A1(n24983), .A2(n25502), .B1(n7451), .B2(n21286), .ZN(
        n5688) );
  OAI22_X1 U23638 ( .A1(n24983), .A2(n25505), .B1(n7449), .B2(n24970), .ZN(
        n5689) );
  OAI22_X1 U23639 ( .A1(n24983), .A2(n25508), .B1(n7447), .B2(n21286), .ZN(
        n5690) );
  OAI22_X1 U23640 ( .A1(n24984), .A2(n25511), .B1(n7445), .B2(n24970), .ZN(
        n5691) );
  OAI22_X1 U23641 ( .A1(n24984), .A2(n25514), .B1(n7443), .B2(n21286), .ZN(
        n5692) );
  OAI22_X1 U23642 ( .A1(n24984), .A2(n25517), .B1(n7441), .B2(n24970), .ZN(
        n5693) );
  OAI22_X1 U23643 ( .A1(n24984), .A2(n25520), .B1(n7439), .B2(n21286), .ZN(
        n5694) );
  OAI22_X1 U23644 ( .A1(n24984), .A2(n25523), .B1(n7437), .B2(n24970), .ZN(
        n5695) );
  OAI22_X1 U23645 ( .A1(n25113), .A2(n25418), .B1(n9068), .B2(n25107), .ZN(
        n6172) );
  OAI22_X1 U23646 ( .A1(n25114), .A2(n25421), .B1(n9066), .B2(n25108), .ZN(
        n6173) );
  OAI22_X1 U23647 ( .A1(n25114), .A2(n25424), .B1(n9064), .B2(n25106), .ZN(
        n6174) );
  OAI22_X1 U23648 ( .A1(n25114), .A2(n25427), .B1(n9062), .B2(n25107), .ZN(
        n6175) );
  OAI22_X1 U23649 ( .A1(n25114), .A2(n25430), .B1(n9060), .B2(n25108), .ZN(
        n6176) );
  OAI22_X1 U23650 ( .A1(n25114), .A2(n25433), .B1(n9058), .B2(n25106), .ZN(
        n6177) );
  OAI22_X1 U23651 ( .A1(n25115), .A2(n25436), .B1(n9056), .B2(n25107), .ZN(
        n6178) );
  OAI22_X1 U23652 ( .A1(n25115), .A2(n25439), .B1(n9054), .B2(n25108), .ZN(
        n6179) );
  OAI22_X1 U23653 ( .A1(n25115), .A2(n25442), .B1(n9052), .B2(n25106), .ZN(
        n6180) );
  OAI22_X1 U23654 ( .A1(n25115), .A2(n25445), .B1(n9050), .B2(n25107), .ZN(
        n6181) );
  OAI22_X1 U23655 ( .A1(n25115), .A2(n25448), .B1(n9048), .B2(n25108), .ZN(
        n6182) );
  OAI22_X1 U23656 ( .A1(n25116), .A2(n25451), .B1(n9046), .B2(n25106), .ZN(
        n6183) );
  OAI22_X1 U23657 ( .A1(n25116), .A2(n25454), .B1(n9044), .B2(n21277), .ZN(
        n6184) );
  OAI22_X1 U23658 ( .A1(n25116), .A2(n25457), .B1(n9042), .B2(n25106), .ZN(
        n6185) );
  OAI22_X1 U23659 ( .A1(n25116), .A2(n25460), .B1(n9040), .B2(n21277), .ZN(
        n6186) );
  OAI22_X1 U23660 ( .A1(n25116), .A2(n25463), .B1(n9038), .B2(n25106), .ZN(
        n6187) );
  OAI22_X1 U23661 ( .A1(n25117), .A2(n25466), .B1(n9036), .B2(n21277), .ZN(
        n6188) );
  OAI22_X1 U23662 ( .A1(n25117), .A2(n25469), .B1(n9034), .B2(n25106), .ZN(
        n6189) );
  OAI22_X1 U23663 ( .A1(n25117), .A2(n25472), .B1(n9032), .B2(n25107), .ZN(
        n6190) );
  OAI22_X1 U23664 ( .A1(n25117), .A2(n25475), .B1(n9030), .B2(n25108), .ZN(
        n6191) );
  OAI22_X1 U23665 ( .A1(n25117), .A2(n25478), .B1(n9028), .B2(n25106), .ZN(
        n6192) );
  OAI22_X1 U23666 ( .A1(n25118), .A2(n25481), .B1(n9026), .B2(n25106), .ZN(
        n6193) );
  OAI22_X1 U23667 ( .A1(n25118), .A2(n25484), .B1(n9024), .B2(n25107), .ZN(
        n6194) );
  OAI22_X1 U23668 ( .A1(n25118), .A2(n25487), .B1(n9022), .B2(n25108), .ZN(
        n6195) );
  OAI22_X1 U23669 ( .A1(n25118), .A2(n25490), .B1(n9020), .B2(n25106), .ZN(
        n6196) );
  OAI22_X1 U23670 ( .A1(n25118), .A2(n25493), .B1(n9018), .B2(n25106), .ZN(
        n6197) );
  OAI22_X1 U23671 ( .A1(n25119), .A2(n25496), .B1(n9016), .B2(n21277), .ZN(
        n6198) );
  OAI22_X1 U23672 ( .A1(n25119), .A2(n25499), .B1(n9014), .B2(n25106), .ZN(
        n6199) );
  OAI22_X1 U23673 ( .A1(n25119), .A2(n25502), .B1(n9012), .B2(n21277), .ZN(
        n6200) );
  OAI22_X1 U23674 ( .A1(n25119), .A2(n25505), .B1(n9010), .B2(n25106), .ZN(
        n6201) );
  OAI22_X1 U23675 ( .A1(n25119), .A2(n25508), .B1(n9008), .B2(n21277), .ZN(
        n6202) );
  OAI22_X1 U23676 ( .A1(n25120), .A2(n25511), .B1(n9006), .B2(n25106), .ZN(
        n6203) );
  OAI22_X1 U23677 ( .A1(n25120), .A2(n25514), .B1(n9004), .B2(n21277), .ZN(
        n6204) );
  OAI22_X1 U23678 ( .A1(n25120), .A2(n25517), .B1(n9002), .B2(n25106), .ZN(
        n6205) );
  OAI22_X1 U23679 ( .A1(n25120), .A2(n25520), .B1(n9000), .B2(n21277), .ZN(
        n6206) );
  OAI22_X1 U23680 ( .A1(n25120), .A2(n25523), .B1(n8998), .B2(n25106), .ZN(
        n6207) );
  OAI22_X1 U23681 ( .A1(n25130), .A2(n25418), .B1(n872), .B2(n25124), .ZN(
        n6236) );
  OAI22_X1 U23682 ( .A1(n25131), .A2(n25421), .B1(n871), .B2(n25125), .ZN(
        n6237) );
  OAI22_X1 U23683 ( .A1(n25131), .A2(n25424), .B1(n870), .B2(n25123), .ZN(
        n6238) );
  OAI22_X1 U23684 ( .A1(n25131), .A2(n25427), .B1(n869), .B2(n25124), .ZN(
        n6239) );
  OAI22_X1 U23685 ( .A1(n25131), .A2(n25430), .B1(n868), .B2(n25125), .ZN(
        n6240) );
  OAI22_X1 U23686 ( .A1(n25131), .A2(n25433), .B1(n867), .B2(n25123), .ZN(
        n6241) );
  OAI22_X1 U23687 ( .A1(n25132), .A2(n25436), .B1(n866), .B2(n25124), .ZN(
        n6242) );
  OAI22_X1 U23688 ( .A1(n25132), .A2(n25439), .B1(n865), .B2(n25125), .ZN(
        n6243) );
  OAI22_X1 U23689 ( .A1(n25132), .A2(n25442), .B1(n864), .B2(n25123), .ZN(
        n6244) );
  OAI22_X1 U23690 ( .A1(n25132), .A2(n25445), .B1(n863), .B2(n25124), .ZN(
        n6245) );
  OAI22_X1 U23691 ( .A1(n25132), .A2(n25448), .B1(n862), .B2(n25125), .ZN(
        n6246) );
  OAI22_X1 U23692 ( .A1(n25133), .A2(n25451), .B1(n861), .B2(n25123), .ZN(
        n6247) );
  OAI22_X1 U23693 ( .A1(n25133), .A2(n25454), .B1(n860), .B2(n21276), .ZN(
        n6248) );
  OAI22_X1 U23694 ( .A1(n25133), .A2(n25457), .B1(n859), .B2(n25123), .ZN(
        n6249) );
  OAI22_X1 U23695 ( .A1(n25133), .A2(n25460), .B1(n858), .B2(n21276), .ZN(
        n6250) );
  OAI22_X1 U23696 ( .A1(n25133), .A2(n25463), .B1(n857), .B2(n25123), .ZN(
        n6251) );
  OAI22_X1 U23697 ( .A1(n25134), .A2(n25466), .B1(n856), .B2(n21276), .ZN(
        n6252) );
  OAI22_X1 U23698 ( .A1(n25134), .A2(n25469), .B1(n855), .B2(n25123), .ZN(
        n6253) );
  OAI22_X1 U23699 ( .A1(n25134), .A2(n25472), .B1(n854), .B2(n25124), .ZN(
        n6254) );
  OAI22_X1 U23700 ( .A1(n25134), .A2(n25475), .B1(n853), .B2(n25125), .ZN(
        n6255) );
  OAI22_X1 U23701 ( .A1(n25134), .A2(n25478), .B1(n852), .B2(n25123), .ZN(
        n6256) );
  OAI22_X1 U23702 ( .A1(n25135), .A2(n25481), .B1(n851), .B2(n25123), .ZN(
        n6257) );
  OAI22_X1 U23703 ( .A1(n25135), .A2(n25484), .B1(n850), .B2(n25124), .ZN(
        n6258) );
  OAI22_X1 U23704 ( .A1(n25135), .A2(n25487), .B1(n849), .B2(n25125), .ZN(
        n6259) );
  OAI22_X1 U23705 ( .A1(n25135), .A2(n25490), .B1(n848), .B2(n25123), .ZN(
        n6260) );
  OAI22_X1 U23706 ( .A1(n25135), .A2(n25493), .B1(n847), .B2(n25123), .ZN(
        n6261) );
  OAI22_X1 U23707 ( .A1(n25136), .A2(n25496), .B1(n846), .B2(n21276), .ZN(
        n6262) );
  OAI22_X1 U23708 ( .A1(n25136), .A2(n25499), .B1(n845), .B2(n25123), .ZN(
        n6263) );
  OAI22_X1 U23709 ( .A1(n25136), .A2(n25502), .B1(n844), .B2(n21276), .ZN(
        n6264) );
  OAI22_X1 U23710 ( .A1(n25136), .A2(n25505), .B1(n843), .B2(n25123), .ZN(
        n6265) );
  OAI22_X1 U23711 ( .A1(n25136), .A2(n25508), .B1(n842), .B2(n21276), .ZN(
        n6266) );
  OAI22_X1 U23712 ( .A1(n25137), .A2(n25511), .B1(n841), .B2(n25123), .ZN(
        n6267) );
  OAI22_X1 U23713 ( .A1(n25137), .A2(n25514), .B1(n840), .B2(n21276), .ZN(
        n6268) );
  OAI22_X1 U23714 ( .A1(n25137), .A2(n25517), .B1(n839), .B2(n25123), .ZN(
        n6269) );
  OAI22_X1 U23715 ( .A1(n25137), .A2(n25520), .B1(n838), .B2(n21276), .ZN(
        n6270) );
  OAI22_X1 U23716 ( .A1(n25137), .A2(n25523), .B1(n837), .B2(n25123), .ZN(
        n6271) );
  OAI22_X1 U23717 ( .A1(n25164), .A2(n25417), .B1(n9196), .B2(n25158), .ZN(
        n6364) );
  OAI22_X1 U23718 ( .A1(n25165), .A2(n25420), .B1(n9194), .B2(n25159), .ZN(
        n6365) );
  OAI22_X1 U23719 ( .A1(n25165), .A2(n25423), .B1(n9192), .B2(n25157), .ZN(
        n6366) );
  OAI22_X1 U23720 ( .A1(n25165), .A2(n25426), .B1(n9190), .B2(n25158), .ZN(
        n6367) );
  OAI22_X1 U23721 ( .A1(n25165), .A2(n25429), .B1(n9188), .B2(n25159), .ZN(
        n6368) );
  OAI22_X1 U23722 ( .A1(n25165), .A2(n25432), .B1(n9186), .B2(n25157), .ZN(
        n6369) );
  OAI22_X1 U23723 ( .A1(n25166), .A2(n25435), .B1(n9184), .B2(n25158), .ZN(
        n6370) );
  OAI22_X1 U23724 ( .A1(n25166), .A2(n25438), .B1(n9182), .B2(n25159), .ZN(
        n6371) );
  OAI22_X1 U23725 ( .A1(n25166), .A2(n25441), .B1(n9180), .B2(n25157), .ZN(
        n6372) );
  OAI22_X1 U23726 ( .A1(n25166), .A2(n25444), .B1(n9178), .B2(n25158), .ZN(
        n6373) );
  OAI22_X1 U23727 ( .A1(n25166), .A2(n25447), .B1(n9176), .B2(n25159), .ZN(
        n6374) );
  OAI22_X1 U23728 ( .A1(n25167), .A2(n25450), .B1(n9174), .B2(n25157), .ZN(
        n6375) );
  OAI22_X1 U23729 ( .A1(n25167), .A2(n25453), .B1(n9172), .B2(n21274), .ZN(
        n6376) );
  OAI22_X1 U23730 ( .A1(n25167), .A2(n25456), .B1(n9170), .B2(n25157), .ZN(
        n6377) );
  OAI22_X1 U23731 ( .A1(n25167), .A2(n25459), .B1(n9168), .B2(n21274), .ZN(
        n6378) );
  OAI22_X1 U23732 ( .A1(n25167), .A2(n25462), .B1(n9166), .B2(n25157), .ZN(
        n6379) );
  OAI22_X1 U23733 ( .A1(n25168), .A2(n25465), .B1(n9164), .B2(n21274), .ZN(
        n6380) );
  OAI22_X1 U23734 ( .A1(n25168), .A2(n25468), .B1(n9162), .B2(n25157), .ZN(
        n6381) );
  OAI22_X1 U23735 ( .A1(n25168), .A2(n25471), .B1(n9160), .B2(n25158), .ZN(
        n6382) );
  OAI22_X1 U23736 ( .A1(n25168), .A2(n25474), .B1(n9158), .B2(n25159), .ZN(
        n6383) );
  OAI22_X1 U23737 ( .A1(n25168), .A2(n25477), .B1(n9156), .B2(n25157), .ZN(
        n6384) );
  OAI22_X1 U23738 ( .A1(n25169), .A2(n25480), .B1(n9154), .B2(n25157), .ZN(
        n6385) );
  OAI22_X1 U23739 ( .A1(n25169), .A2(n25483), .B1(n9152), .B2(n25158), .ZN(
        n6386) );
  OAI22_X1 U23740 ( .A1(n25169), .A2(n25486), .B1(n9150), .B2(n25159), .ZN(
        n6387) );
  OAI22_X1 U23741 ( .A1(n25169), .A2(n25489), .B1(n9148), .B2(n25157), .ZN(
        n6388) );
  OAI22_X1 U23742 ( .A1(n25169), .A2(n25492), .B1(n9146), .B2(n25157), .ZN(
        n6389) );
  OAI22_X1 U23743 ( .A1(n25170), .A2(n25495), .B1(n9144), .B2(n21274), .ZN(
        n6390) );
  OAI22_X1 U23744 ( .A1(n25170), .A2(n25498), .B1(n9142), .B2(n25157), .ZN(
        n6391) );
  OAI22_X1 U23745 ( .A1(n25170), .A2(n25501), .B1(n9140), .B2(n21274), .ZN(
        n6392) );
  OAI22_X1 U23746 ( .A1(n25170), .A2(n25504), .B1(n9138), .B2(n25157), .ZN(
        n6393) );
  OAI22_X1 U23747 ( .A1(n25170), .A2(n25507), .B1(n9136), .B2(n21274), .ZN(
        n6394) );
  OAI22_X1 U23748 ( .A1(n25171), .A2(n25510), .B1(n9134), .B2(n25157), .ZN(
        n6395) );
  OAI22_X1 U23749 ( .A1(n25171), .A2(n25513), .B1(n9132), .B2(n21274), .ZN(
        n6396) );
  OAI22_X1 U23750 ( .A1(n25171), .A2(n25516), .B1(n9130), .B2(n25157), .ZN(
        n6397) );
  OAI22_X1 U23751 ( .A1(n25171), .A2(n25519), .B1(n9128), .B2(n21274), .ZN(
        n6398) );
  OAI22_X1 U23752 ( .A1(n25171), .A2(n25522), .B1(n9126), .B2(n25157), .ZN(
        n6399) );
  OAI22_X1 U23753 ( .A1(n25274), .A2(n25525), .B1(n17230), .B2(n21263), .ZN(
        n6784) );
  OAI22_X1 U23754 ( .A1(n25274), .A2(n25528), .B1(n17227), .B2(n21263), .ZN(
        n6785) );
  OAI22_X1 U23755 ( .A1(n25274), .A2(n25531), .B1(n17224), .B2(n25259), .ZN(
        n6786) );
  OAI22_X1 U23756 ( .A1(n25274), .A2(n25551), .B1(n17221), .B2(n21263), .ZN(
        n6787) );
  OAI22_X1 U23757 ( .A1(n24968), .A2(n25526), .B1(n9125), .B2(n21287), .ZN(
        n5632) );
  OAI22_X1 U23758 ( .A1(n24968), .A2(n25529), .B1(n9123), .B2(n21287), .ZN(
        n5633) );
  OAI22_X1 U23759 ( .A1(n24968), .A2(n25532), .B1(n9121), .B2(n24953), .ZN(
        n5634) );
  OAI22_X1 U23760 ( .A1(n24968), .A2(n25552), .B1(n9119), .B2(n21287), .ZN(
        n5635) );
  OAI22_X1 U23761 ( .A1(n25036), .A2(n25526), .B1(n8869), .B2(n21283), .ZN(
        n5888) );
  OAI22_X1 U23762 ( .A1(n25036), .A2(n25529), .B1(n8867), .B2(n21283), .ZN(
        n5889) );
  OAI22_X1 U23763 ( .A1(n25036), .A2(n25532), .B1(n8865), .B2(n25021), .ZN(
        n5890) );
  OAI22_X1 U23764 ( .A1(n25036), .A2(n25552), .B1(n8863), .B2(n21283), .ZN(
        n5891) );
  OAI22_X1 U23765 ( .A1(n24866), .A2(n25527), .B1(n8868), .B2(n21294), .ZN(
        n5248) );
  OAI22_X1 U23766 ( .A1(n24866), .A2(n25530), .B1(n8866), .B2(n21294), .ZN(
        n5249) );
  OAI22_X1 U23767 ( .A1(n24866), .A2(n25533), .B1(n8864), .B2(n24851), .ZN(
        n5250) );
  OAI22_X1 U23768 ( .A1(n24866), .A2(n25553), .B1(n8862), .B2(n21294), .ZN(
        n5251) );
  OAI22_X1 U23769 ( .A1(n25172), .A2(n25525), .B1(n9124), .B2(n21274), .ZN(
        n6400) );
  OAI22_X1 U23770 ( .A1(n25172), .A2(n25528), .B1(n9122), .B2(n21274), .ZN(
        n6401) );
  OAI22_X1 U23771 ( .A1(n25172), .A2(n25531), .B1(n9120), .B2(n25157), .ZN(
        n6402) );
  OAI22_X1 U23772 ( .A1(n25172), .A2(n25551), .B1(n9118), .B2(n21274), .ZN(
        n6403) );
  OAI22_X1 U23773 ( .A1(n25189), .A2(n25525), .B1(n7434), .B2(n21273), .ZN(
        n6464) );
  OAI22_X1 U23774 ( .A1(n25189), .A2(n25528), .B1(n7432), .B2(n21273), .ZN(
        n6465) );
  OAI22_X1 U23775 ( .A1(n25189), .A2(n25531), .B1(n7430), .B2(n25174), .ZN(
        n6466) );
  OAI22_X1 U23776 ( .A1(n25189), .A2(n25551), .B1(n7428), .B2(n21273), .ZN(
        n6467) );
  OAI22_X1 U23777 ( .A1(n24934), .A2(n25527), .B1(n7307), .B2(n21290), .ZN(
        n5504) );
  OAI22_X1 U23778 ( .A1(n24934), .A2(n25530), .B1(n7305), .B2(n21290), .ZN(
        n5505) );
  OAI22_X1 U23779 ( .A1(n24934), .A2(n25533), .B1(n7303), .B2(n24919), .ZN(
        n5506) );
  OAI22_X1 U23780 ( .A1(n24934), .A2(n25553), .B1(n7301), .B2(n21290), .ZN(
        n5507) );
  OAI22_X1 U23781 ( .A1(n25138), .A2(n25526), .B1(n836), .B2(n21276), .ZN(
        n6272) );
  OAI22_X1 U23782 ( .A1(n25138), .A2(n25529), .B1(n835), .B2(n21276), .ZN(
        n6273) );
  OAI22_X1 U23783 ( .A1(n25138), .A2(n25532), .B1(n834), .B2(n25123), .ZN(
        n6274) );
  OAI22_X1 U23784 ( .A1(n25138), .A2(n25552), .B1(n833), .B2(n21276), .ZN(
        n6275) );
  OAI22_X1 U23785 ( .A1(n25053), .A2(n25526), .B1(n8741), .B2(n21282), .ZN(
        n5952) );
  OAI22_X1 U23786 ( .A1(n25053), .A2(n25529), .B1(n8739), .B2(n21282), .ZN(
        n5953) );
  OAI22_X1 U23787 ( .A1(n25053), .A2(n25532), .B1(n8737), .B2(n25038), .ZN(
        n5954) );
  OAI22_X1 U23788 ( .A1(n25053), .A2(n25552), .B1(n8735), .B2(n21282), .ZN(
        n5955) );
  OAI22_X1 U23789 ( .A1(n24985), .A2(n25526), .B1(n7435), .B2(n21286), .ZN(
        n5696) );
  OAI22_X1 U23790 ( .A1(n24985), .A2(n25529), .B1(n7433), .B2(n21286), .ZN(
        n5697) );
  OAI22_X1 U23791 ( .A1(n24985), .A2(n25532), .B1(n7431), .B2(n24970), .ZN(
        n5698) );
  OAI22_X1 U23792 ( .A1(n24985), .A2(n25552), .B1(n7429), .B2(n21286), .ZN(
        n5699) );
  OAI22_X1 U23793 ( .A1(n25121), .A2(n25526), .B1(n8996), .B2(n21277), .ZN(
        n6208) );
  OAI22_X1 U23794 ( .A1(n25121), .A2(n25529), .B1(n8994), .B2(n21277), .ZN(
        n6209) );
  OAI22_X1 U23795 ( .A1(n25121), .A2(n25532), .B1(n8992), .B2(n25106), .ZN(
        n6210) );
  OAI22_X1 U23796 ( .A1(n25121), .A2(n25552), .B1(n8990), .B2(n21277), .ZN(
        n6211) );
  OAI22_X1 U23797 ( .A1(n24900), .A2(n25527), .B1(n21292), .B2(n20530), .ZN(
        n5376) );
  OAI22_X1 U23798 ( .A1(n24900), .A2(n25530), .B1(n21292), .B2(n20529), .ZN(
        n5377) );
  OAI22_X1 U23799 ( .A1(n24900), .A2(n25533), .B1(n24885), .B2(n20528), .ZN(
        n5378) );
  OAI22_X1 U23800 ( .A1(n24900), .A2(n25553), .B1(n21292), .B2(n20527), .ZN(
        n5379) );
  OAI221_X1 U23801 ( .B1(n19207), .B2(n24809), .C1(n11843), .C2(n24798), .A(
        n21389), .ZN(n5056) );
  OAI21_X1 U23802 ( .B1(n21390), .B2(n21391), .A(n24797), .ZN(n21389) );
  NAND4_X1 U23803 ( .A1(n21400), .A2(n21401), .A3(n21402), .A4(n21403), .ZN(
        n21390) );
  NAND4_X1 U23804 ( .A1(n21392), .A2(n21393), .A3(n21394), .A4(n21395), .ZN(
        n21391) );
  OAI221_X1 U23805 ( .B1(n19206), .B2(n24809), .C1(n11844), .C2(n24798), .A(
        n21370), .ZN(n5057) );
  OAI21_X1 U23806 ( .B1(n21371), .B2(n21372), .A(n24797), .ZN(n21370) );
  NAND4_X1 U23807 ( .A1(n21381), .A2(n21382), .A3(n21383), .A4(n21384), .ZN(
        n21371) );
  NAND4_X1 U23808 ( .A1(n21373), .A2(n21374), .A3(n21375), .A4(n21376), .ZN(
        n21372) );
  OAI221_X1 U23809 ( .B1(n19205), .B2(n24809), .C1(n11845), .C2(n24798), .A(
        n21351), .ZN(n5058) );
  OAI21_X1 U23810 ( .B1(n21352), .B2(n21353), .A(n24797), .ZN(n21351) );
  NAND4_X1 U23811 ( .A1(n21362), .A2(n21363), .A3(n21364), .A4(n21365), .ZN(
        n21352) );
  NAND4_X1 U23812 ( .A1(n21354), .A2(n21355), .A3(n21356), .A4(n21357), .ZN(
        n21353) );
  OAI221_X1 U23813 ( .B1(n19204), .B2(n24809), .C1(n11846), .C2(n24800), .A(
        n21299), .ZN(n5059) );
  OAI21_X1 U23814 ( .B1(n21300), .B2(n21301), .A(n24797), .ZN(n21299) );
  NAND4_X1 U23815 ( .A1(n21327), .A2(n21328), .A3(n21329), .A4(n21330), .ZN(
        n21300) );
  NAND4_X1 U23816 ( .A1(n21303), .A2(n21304), .A3(n21305), .A4(n21306), .ZN(
        n21301) );
  OAI221_X1 U23817 ( .B1(n19267), .B2(n24804), .C1(n11783), .C2(n24803), .A(
        n22529), .ZN(n4996) );
  OAI21_X1 U23818 ( .B1(n22530), .B2(n22531), .A(n24792), .ZN(n22529) );
  NAND4_X1 U23819 ( .A1(n22548), .A2(n22549), .A3(n22550), .A4(n22551), .ZN(
        n22530) );
  NAND4_X1 U23820 ( .A1(n22532), .A2(n22533), .A3(n22534), .A4(n22535), .ZN(
        n22531) );
  OAI221_X1 U23821 ( .B1(n19266), .B2(n24804), .C1(n11784), .C2(n24803), .A(
        n22510), .ZN(n4997) );
  OAI21_X1 U23822 ( .B1(n22511), .B2(n22512), .A(n24792), .ZN(n22510) );
  NAND4_X1 U23823 ( .A1(n22521), .A2(n22522), .A3(n22523), .A4(n22524), .ZN(
        n22511) );
  NAND4_X1 U23824 ( .A1(n22513), .A2(n22514), .A3(n22515), .A4(n22516), .ZN(
        n22512) );
  OAI221_X1 U23825 ( .B1(n19265), .B2(n24804), .C1(n11785), .C2(n24803), .A(
        n22491), .ZN(n4998) );
  OAI21_X1 U23826 ( .B1(n22492), .B2(n22493), .A(n24792), .ZN(n22491) );
  NAND4_X1 U23827 ( .A1(n22502), .A2(n22503), .A3(n22504), .A4(n22505), .ZN(
        n22492) );
  NAND4_X1 U23828 ( .A1(n22494), .A2(n22495), .A3(n22496), .A4(n22497), .ZN(
        n22493) );
  OAI221_X1 U23829 ( .B1(n19264), .B2(n24804), .C1(n11786), .C2(n24803), .A(
        n22472), .ZN(n4999) );
  OAI21_X1 U23830 ( .B1(n22473), .B2(n22474), .A(n24792), .ZN(n22472) );
  NAND4_X1 U23831 ( .A1(n22483), .A2(n22484), .A3(n22485), .A4(n22486), .ZN(
        n22473) );
  NAND4_X1 U23832 ( .A1(n22475), .A2(n22476), .A3(n22477), .A4(n22478), .ZN(
        n22474) );
  OAI221_X1 U23833 ( .B1(n19263), .B2(n24804), .C1(n11787), .C2(n24802), .A(
        n22453), .ZN(n5000) );
  OAI21_X1 U23834 ( .B1(n22454), .B2(n22455), .A(n24792), .ZN(n22453) );
  NAND4_X1 U23835 ( .A1(n22464), .A2(n22465), .A3(n22466), .A4(n22467), .ZN(
        n22454) );
  NAND4_X1 U23836 ( .A1(n22456), .A2(n22457), .A3(n22458), .A4(n22459), .ZN(
        n22455) );
  OAI221_X1 U23837 ( .B1(n19262), .B2(n24804), .C1(n11788), .C2(n24802), .A(
        n22434), .ZN(n5001) );
  OAI21_X1 U23838 ( .B1(n22435), .B2(n22436), .A(n24792), .ZN(n22434) );
  NAND4_X1 U23839 ( .A1(n22445), .A2(n22446), .A3(n22447), .A4(n22448), .ZN(
        n22435) );
  NAND4_X1 U23840 ( .A1(n22437), .A2(n22438), .A3(n22439), .A4(n22440), .ZN(
        n22436) );
  OAI221_X1 U23841 ( .B1(n19261), .B2(n24804), .C1(n11789), .C2(n24802), .A(
        n22415), .ZN(n5002) );
  OAI21_X1 U23842 ( .B1(n22416), .B2(n22417), .A(n24792), .ZN(n22415) );
  NAND4_X1 U23843 ( .A1(n22426), .A2(n22427), .A3(n22428), .A4(n22429), .ZN(
        n22416) );
  NAND4_X1 U23844 ( .A1(n22418), .A2(n22419), .A3(n22420), .A4(n22421), .ZN(
        n22417) );
  OAI221_X1 U23845 ( .B1(n19260), .B2(n24804), .C1(n11790), .C2(n24802), .A(
        n22396), .ZN(n5003) );
  OAI21_X1 U23846 ( .B1(n22397), .B2(n22398), .A(n24792), .ZN(n22396) );
  NAND4_X1 U23847 ( .A1(n22407), .A2(n22408), .A3(n22409), .A4(n22410), .ZN(
        n22397) );
  NAND4_X1 U23848 ( .A1(n22399), .A2(n22400), .A3(n22401), .A4(n22402), .ZN(
        n22398) );
  OAI221_X1 U23849 ( .B1(n19259), .B2(n24804), .C1(n11791), .C2(n24802), .A(
        n22377), .ZN(n5004) );
  OAI21_X1 U23850 ( .B1(n22378), .B2(n22379), .A(n24792), .ZN(n22377) );
  NAND4_X1 U23851 ( .A1(n22388), .A2(n22389), .A3(n22390), .A4(n22391), .ZN(
        n22378) );
  NAND4_X1 U23852 ( .A1(n22380), .A2(n22381), .A3(n22382), .A4(n22383), .ZN(
        n22379) );
  OAI221_X1 U23853 ( .B1(n19258), .B2(n24804), .C1(n11792), .C2(n24802), .A(
        n22358), .ZN(n5005) );
  OAI21_X1 U23854 ( .B1(n22359), .B2(n22360), .A(n24792), .ZN(n22358) );
  NAND4_X1 U23855 ( .A1(n22369), .A2(n22370), .A3(n22371), .A4(n22372), .ZN(
        n22359) );
  NAND4_X1 U23856 ( .A1(n22361), .A2(n22362), .A3(n22363), .A4(n22364), .ZN(
        n22360) );
  OAI221_X1 U23857 ( .B1(n19257), .B2(n24804), .C1(n11793), .C2(n24802), .A(
        n22339), .ZN(n5006) );
  OAI21_X1 U23858 ( .B1(n22340), .B2(n22341), .A(n24792), .ZN(n22339) );
  NAND4_X1 U23859 ( .A1(n22350), .A2(n22351), .A3(n22352), .A4(n22353), .ZN(
        n22340) );
  NAND4_X1 U23860 ( .A1(n22342), .A2(n22343), .A3(n22344), .A4(n22345), .ZN(
        n22341) );
  OAI221_X1 U23861 ( .B1(n19256), .B2(n24804), .C1(n11794), .C2(n24802), .A(
        n22320), .ZN(n5007) );
  OAI21_X1 U23862 ( .B1(n22321), .B2(n22322), .A(n24792), .ZN(n22320) );
  NAND4_X1 U23863 ( .A1(n22331), .A2(n22332), .A3(n22333), .A4(n22334), .ZN(
        n22321) );
  NAND4_X1 U23864 ( .A1(n22323), .A2(n22324), .A3(n22325), .A4(n22326), .ZN(
        n22322) );
  OAI221_X1 U23865 ( .B1(n19255), .B2(n24805), .C1(n11795), .C2(n24802), .A(
        n22301), .ZN(n5008) );
  OAI21_X1 U23866 ( .B1(n22302), .B2(n22303), .A(n24793), .ZN(n22301) );
  NAND4_X1 U23867 ( .A1(n22312), .A2(n22313), .A3(n22314), .A4(n22315), .ZN(
        n22302) );
  NAND4_X1 U23868 ( .A1(n22304), .A2(n22305), .A3(n22306), .A4(n22307), .ZN(
        n22303) );
  OAI221_X1 U23869 ( .B1(n19254), .B2(n24805), .C1(n11796), .C2(n24802), .A(
        n22282), .ZN(n5009) );
  OAI21_X1 U23870 ( .B1(n22283), .B2(n22284), .A(n24793), .ZN(n22282) );
  NAND4_X1 U23871 ( .A1(n22293), .A2(n22294), .A3(n22295), .A4(n22296), .ZN(
        n22283) );
  NAND4_X1 U23872 ( .A1(n22285), .A2(n22286), .A3(n22287), .A4(n22288), .ZN(
        n22284) );
  OAI221_X1 U23873 ( .B1(n19253), .B2(n24805), .C1(n11797), .C2(n24802), .A(
        n22263), .ZN(n5010) );
  OAI21_X1 U23874 ( .B1(n22264), .B2(n22265), .A(n24793), .ZN(n22263) );
  NAND4_X1 U23875 ( .A1(n22274), .A2(n22275), .A3(n22276), .A4(n22277), .ZN(
        n22264) );
  NAND4_X1 U23876 ( .A1(n22266), .A2(n22267), .A3(n22268), .A4(n22269), .ZN(
        n22265) );
  OAI221_X1 U23877 ( .B1(n19252), .B2(n24805), .C1(n11798), .C2(n24802), .A(
        n22244), .ZN(n5011) );
  OAI21_X1 U23878 ( .B1(n22245), .B2(n22246), .A(n24793), .ZN(n22244) );
  NAND4_X1 U23879 ( .A1(n22255), .A2(n22256), .A3(n22257), .A4(n22258), .ZN(
        n22245) );
  NAND4_X1 U23880 ( .A1(n22247), .A2(n22248), .A3(n22249), .A4(n22250), .ZN(
        n22246) );
  OAI221_X1 U23881 ( .B1(n19251), .B2(n24805), .C1(n11799), .C2(n24801), .A(
        n22225), .ZN(n5012) );
  OAI21_X1 U23882 ( .B1(n22226), .B2(n22227), .A(n24793), .ZN(n22225) );
  NAND4_X1 U23883 ( .A1(n22236), .A2(n22237), .A3(n22238), .A4(n22239), .ZN(
        n22226) );
  NAND4_X1 U23884 ( .A1(n22228), .A2(n22229), .A3(n22230), .A4(n22231), .ZN(
        n22227) );
  OAI221_X1 U23885 ( .B1(n19250), .B2(n24805), .C1(n11800), .C2(n24801), .A(
        n22206), .ZN(n5013) );
  OAI21_X1 U23886 ( .B1(n22207), .B2(n22208), .A(n24793), .ZN(n22206) );
  NAND4_X1 U23887 ( .A1(n22217), .A2(n22218), .A3(n22219), .A4(n22220), .ZN(
        n22207) );
  NAND4_X1 U23888 ( .A1(n22209), .A2(n22210), .A3(n22211), .A4(n22212), .ZN(
        n22208) );
  OAI221_X1 U23889 ( .B1(n19249), .B2(n24805), .C1(n11801), .C2(n24801), .A(
        n22187), .ZN(n5014) );
  OAI21_X1 U23890 ( .B1(n22188), .B2(n22189), .A(n24793), .ZN(n22187) );
  NAND4_X1 U23891 ( .A1(n22198), .A2(n22199), .A3(n22200), .A4(n22201), .ZN(
        n22188) );
  NAND4_X1 U23892 ( .A1(n22190), .A2(n22191), .A3(n22192), .A4(n22193), .ZN(
        n22189) );
  OAI221_X1 U23893 ( .B1(n19248), .B2(n24805), .C1(n11802), .C2(n24801), .A(
        n22168), .ZN(n5015) );
  OAI21_X1 U23894 ( .B1(n22169), .B2(n22170), .A(n24793), .ZN(n22168) );
  NAND4_X1 U23895 ( .A1(n22179), .A2(n22180), .A3(n22181), .A4(n22182), .ZN(
        n22169) );
  NAND4_X1 U23896 ( .A1(n22171), .A2(n22172), .A3(n22173), .A4(n22174), .ZN(
        n22170) );
  OAI221_X1 U23897 ( .B1(n19247), .B2(n24805), .C1(n11803), .C2(n24801), .A(
        n22149), .ZN(n5016) );
  OAI21_X1 U23898 ( .B1(n22150), .B2(n22151), .A(n24793), .ZN(n22149) );
  NAND4_X1 U23899 ( .A1(n22160), .A2(n22161), .A3(n22162), .A4(n22163), .ZN(
        n22150) );
  NAND4_X1 U23900 ( .A1(n22152), .A2(n22153), .A3(n22154), .A4(n22155), .ZN(
        n22151) );
  OAI221_X1 U23901 ( .B1(n19246), .B2(n24805), .C1(n11804), .C2(n24801), .A(
        n22130), .ZN(n5017) );
  OAI21_X1 U23902 ( .B1(n22131), .B2(n22132), .A(n24793), .ZN(n22130) );
  NAND4_X1 U23903 ( .A1(n22141), .A2(n22142), .A3(n22143), .A4(n22144), .ZN(
        n22131) );
  NAND4_X1 U23904 ( .A1(n22133), .A2(n22134), .A3(n22135), .A4(n22136), .ZN(
        n22132) );
  OAI221_X1 U23905 ( .B1(n19245), .B2(n24805), .C1(n11805), .C2(n24801), .A(
        n22111), .ZN(n5018) );
  OAI21_X1 U23906 ( .B1(n22112), .B2(n22113), .A(n24793), .ZN(n22111) );
  NAND4_X1 U23907 ( .A1(n22122), .A2(n22123), .A3(n22124), .A4(n22125), .ZN(
        n22112) );
  NAND4_X1 U23908 ( .A1(n22114), .A2(n22115), .A3(n22116), .A4(n22117), .ZN(
        n22113) );
  OAI221_X1 U23909 ( .B1(n19244), .B2(n24805), .C1(n11806), .C2(n24801), .A(
        n22092), .ZN(n5019) );
  OAI21_X1 U23910 ( .B1(n22093), .B2(n22094), .A(n24793), .ZN(n22092) );
  NAND4_X1 U23911 ( .A1(n22103), .A2(n22104), .A3(n22105), .A4(n22106), .ZN(
        n22093) );
  NAND4_X1 U23912 ( .A1(n22095), .A2(n22096), .A3(n22097), .A4(n22098), .ZN(
        n22094) );
  OAI221_X1 U23913 ( .B1(n19243), .B2(n24806), .C1(n11807), .C2(n24801), .A(
        n22073), .ZN(n5020) );
  OAI21_X1 U23914 ( .B1(n22074), .B2(n22075), .A(n24794), .ZN(n22073) );
  NAND4_X1 U23915 ( .A1(n22084), .A2(n22085), .A3(n22086), .A4(n22087), .ZN(
        n22074) );
  NAND4_X1 U23916 ( .A1(n22076), .A2(n22077), .A3(n22078), .A4(n22079), .ZN(
        n22075) );
  OAI221_X1 U23917 ( .B1(n19242), .B2(n24806), .C1(n11808), .C2(n24801), .A(
        n22054), .ZN(n5021) );
  OAI21_X1 U23918 ( .B1(n22055), .B2(n22056), .A(n24794), .ZN(n22054) );
  NAND4_X1 U23919 ( .A1(n22065), .A2(n22066), .A3(n22067), .A4(n22068), .ZN(
        n22055) );
  NAND4_X1 U23920 ( .A1(n22057), .A2(n22058), .A3(n22059), .A4(n22060), .ZN(
        n22056) );
  OAI221_X1 U23921 ( .B1(n19241), .B2(n24806), .C1(n11809), .C2(n24801), .A(
        n22035), .ZN(n5022) );
  OAI21_X1 U23922 ( .B1(n22036), .B2(n22037), .A(n24794), .ZN(n22035) );
  NAND4_X1 U23923 ( .A1(n22046), .A2(n22047), .A3(n22048), .A4(n22049), .ZN(
        n22036) );
  NAND4_X1 U23924 ( .A1(n22038), .A2(n22039), .A3(n22040), .A4(n22041), .ZN(
        n22037) );
  OAI221_X1 U23925 ( .B1(n19240), .B2(n24806), .C1(n11810), .C2(n24801), .A(
        n22016), .ZN(n5023) );
  OAI21_X1 U23926 ( .B1(n22017), .B2(n22018), .A(n24794), .ZN(n22016) );
  NAND4_X1 U23927 ( .A1(n22027), .A2(n22028), .A3(n22029), .A4(n22030), .ZN(
        n22017) );
  NAND4_X1 U23928 ( .A1(n22019), .A2(n22020), .A3(n22021), .A4(n22022), .ZN(
        n22018) );
  OAI221_X1 U23929 ( .B1(n19239), .B2(n24806), .C1(n11811), .C2(n24800), .A(
        n21997), .ZN(n5024) );
  OAI21_X1 U23930 ( .B1(n21998), .B2(n21999), .A(n24794), .ZN(n21997) );
  NAND4_X1 U23931 ( .A1(n22008), .A2(n22009), .A3(n22010), .A4(n22011), .ZN(
        n21998) );
  NAND4_X1 U23932 ( .A1(n22000), .A2(n22001), .A3(n22002), .A4(n22003), .ZN(
        n21999) );
  OAI221_X1 U23933 ( .B1(n19238), .B2(n24806), .C1(n11812), .C2(n24800), .A(
        n21978), .ZN(n5025) );
  OAI21_X1 U23934 ( .B1(n21979), .B2(n21980), .A(n24794), .ZN(n21978) );
  NAND4_X1 U23935 ( .A1(n21989), .A2(n21990), .A3(n21991), .A4(n21992), .ZN(
        n21979) );
  NAND4_X1 U23936 ( .A1(n21981), .A2(n21982), .A3(n21983), .A4(n21984), .ZN(
        n21980) );
  OAI221_X1 U23937 ( .B1(n19237), .B2(n24806), .C1(n11813), .C2(n24800), .A(
        n21959), .ZN(n5026) );
  OAI21_X1 U23938 ( .B1(n21960), .B2(n21961), .A(n24794), .ZN(n21959) );
  NAND4_X1 U23939 ( .A1(n21970), .A2(n21971), .A3(n21972), .A4(n21973), .ZN(
        n21960) );
  NAND4_X1 U23940 ( .A1(n21962), .A2(n21963), .A3(n21964), .A4(n21965), .ZN(
        n21961) );
  OAI221_X1 U23941 ( .B1(n19236), .B2(n24806), .C1(n11814), .C2(n24800), .A(
        n21940), .ZN(n5027) );
  OAI21_X1 U23942 ( .B1(n21941), .B2(n21942), .A(n24794), .ZN(n21940) );
  NAND4_X1 U23943 ( .A1(n21951), .A2(n21952), .A3(n21953), .A4(n21954), .ZN(
        n21941) );
  NAND4_X1 U23944 ( .A1(n21943), .A2(n21944), .A3(n21945), .A4(n21946), .ZN(
        n21942) );
  OAI221_X1 U23945 ( .B1(n19235), .B2(n24806), .C1(n11815), .C2(n24800), .A(
        n21921), .ZN(n5028) );
  OAI21_X1 U23946 ( .B1(n21922), .B2(n21923), .A(n24794), .ZN(n21921) );
  NAND4_X1 U23947 ( .A1(n21932), .A2(n21933), .A3(n21934), .A4(n21935), .ZN(
        n21922) );
  NAND4_X1 U23948 ( .A1(n21924), .A2(n21925), .A3(n21926), .A4(n21927), .ZN(
        n21923) );
  OAI221_X1 U23949 ( .B1(n19234), .B2(n24806), .C1(n11816), .C2(n24800), .A(
        n21902), .ZN(n5029) );
  OAI21_X1 U23950 ( .B1(n21903), .B2(n21904), .A(n24794), .ZN(n21902) );
  NAND4_X1 U23951 ( .A1(n21913), .A2(n21914), .A3(n21915), .A4(n21916), .ZN(
        n21903) );
  NAND4_X1 U23952 ( .A1(n21905), .A2(n21906), .A3(n21907), .A4(n21908), .ZN(
        n21904) );
  OAI221_X1 U23953 ( .B1(n19233), .B2(n24806), .C1(n11817), .C2(n24800), .A(
        n21883), .ZN(n5030) );
  OAI21_X1 U23954 ( .B1(n21884), .B2(n21885), .A(n24794), .ZN(n21883) );
  NAND4_X1 U23955 ( .A1(n21894), .A2(n21895), .A3(n21896), .A4(n21897), .ZN(
        n21884) );
  NAND4_X1 U23956 ( .A1(n21886), .A2(n21887), .A3(n21888), .A4(n21889), .ZN(
        n21885) );
  OAI221_X1 U23957 ( .B1(n19232), .B2(n24806), .C1(n11818), .C2(n24800), .A(
        n21864), .ZN(n5031) );
  OAI21_X1 U23958 ( .B1(n21865), .B2(n21866), .A(n24794), .ZN(n21864) );
  NAND4_X1 U23959 ( .A1(n21875), .A2(n21876), .A3(n21877), .A4(n21878), .ZN(
        n21865) );
  NAND4_X1 U23960 ( .A1(n21867), .A2(n21868), .A3(n21869), .A4(n21870), .ZN(
        n21866) );
  OAI221_X1 U23961 ( .B1(n19231), .B2(n24807), .C1(n11819), .C2(n24800), .A(
        n21845), .ZN(n5032) );
  OAI21_X1 U23962 ( .B1(n21846), .B2(n21847), .A(n24795), .ZN(n21845) );
  NAND4_X1 U23963 ( .A1(n21856), .A2(n21857), .A3(n21858), .A4(n21859), .ZN(
        n21846) );
  NAND4_X1 U23964 ( .A1(n21848), .A2(n21849), .A3(n21850), .A4(n21851), .ZN(
        n21847) );
  OAI221_X1 U23965 ( .B1(n19230), .B2(n24807), .C1(n11820), .C2(n24800), .A(
        n21826), .ZN(n5033) );
  OAI21_X1 U23966 ( .B1(n21827), .B2(n21828), .A(n24795), .ZN(n21826) );
  NAND4_X1 U23967 ( .A1(n21837), .A2(n21838), .A3(n21839), .A4(n21840), .ZN(
        n21827) );
  NAND4_X1 U23968 ( .A1(n21829), .A2(n21830), .A3(n21831), .A4(n21832), .ZN(
        n21828) );
  OAI221_X1 U23969 ( .B1(n19229), .B2(n24807), .C1(n11821), .C2(n24800), .A(
        n21807), .ZN(n5034) );
  OAI21_X1 U23970 ( .B1(n21808), .B2(n21809), .A(n24795), .ZN(n21807) );
  NAND4_X1 U23971 ( .A1(n21818), .A2(n21819), .A3(n21820), .A4(n21821), .ZN(
        n21808) );
  NAND4_X1 U23972 ( .A1(n21810), .A2(n21811), .A3(n21812), .A4(n21813), .ZN(
        n21809) );
  OAI221_X1 U23973 ( .B1(n19228), .B2(n24807), .C1(n11822), .C2(n24799), .A(
        n21788), .ZN(n5035) );
  OAI21_X1 U23974 ( .B1(n21789), .B2(n21790), .A(n24795), .ZN(n21788) );
  NAND4_X1 U23975 ( .A1(n21799), .A2(n21800), .A3(n21801), .A4(n21802), .ZN(
        n21789) );
  NAND4_X1 U23976 ( .A1(n21791), .A2(n21792), .A3(n21793), .A4(n21794), .ZN(
        n21790) );
  OAI221_X1 U23977 ( .B1(n19227), .B2(n24807), .C1(n11823), .C2(n24799), .A(
        n21769), .ZN(n5036) );
  OAI21_X1 U23978 ( .B1(n21770), .B2(n21771), .A(n24795), .ZN(n21769) );
  NAND4_X1 U23979 ( .A1(n21780), .A2(n21781), .A3(n21782), .A4(n21783), .ZN(
        n21770) );
  NAND4_X1 U23980 ( .A1(n21772), .A2(n21773), .A3(n21774), .A4(n21775), .ZN(
        n21771) );
  OAI221_X1 U23981 ( .B1(n19226), .B2(n24807), .C1(n11824), .C2(n24799), .A(
        n21750), .ZN(n5037) );
  OAI21_X1 U23982 ( .B1(n21751), .B2(n21752), .A(n24795), .ZN(n21750) );
  NAND4_X1 U23983 ( .A1(n21761), .A2(n21762), .A3(n21763), .A4(n21764), .ZN(
        n21751) );
  NAND4_X1 U23984 ( .A1(n21753), .A2(n21754), .A3(n21755), .A4(n21756), .ZN(
        n21752) );
  OAI221_X1 U23985 ( .B1(n19225), .B2(n24807), .C1(n11825), .C2(n24799), .A(
        n21731), .ZN(n5038) );
  OAI21_X1 U23986 ( .B1(n21732), .B2(n21733), .A(n24795), .ZN(n21731) );
  NAND4_X1 U23987 ( .A1(n21742), .A2(n21743), .A3(n21744), .A4(n21745), .ZN(
        n21732) );
  NAND4_X1 U23988 ( .A1(n21734), .A2(n21735), .A3(n21736), .A4(n21737), .ZN(
        n21733) );
  OAI221_X1 U23989 ( .B1(n19224), .B2(n24807), .C1(n11826), .C2(n24799), .A(
        n21712), .ZN(n5039) );
  OAI21_X1 U23990 ( .B1(n21713), .B2(n21714), .A(n24795), .ZN(n21712) );
  NAND4_X1 U23991 ( .A1(n21723), .A2(n21724), .A3(n21725), .A4(n21726), .ZN(
        n21713) );
  NAND4_X1 U23992 ( .A1(n21715), .A2(n21716), .A3(n21717), .A4(n21718), .ZN(
        n21714) );
  OAI221_X1 U23993 ( .B1(n19223), .B2(n24807), .C1(n11827), .C2(n24799), .A(
        n21693), .ZN(n5040) );
  OAI21_X1 U23994 ( .B1(n21694), .B2(n21695), .A(n24795), .ZN(n21693) );
  NAND4_X1 U23995 ( .A1(n21704), .A2(n21705), .A3(n21706), .A4(n21707), .ZN(
        n21694) );
  NAND4_X1 U23996 ( .A1(n21696), .A2(n21697), .A3(n21698), .A4(n21699), .ZN(
        n21695) );
  OAI221_X1 U23997 ( .B1(n19222), .B2(n24807), .C1(n11828), .C2(n24799), .A(
        n21674), .ZN(n5041) );
  OAI21_X1 U23998 ( .B1(n21675), .B2(n21676), .A(n24795), .ZN(n21674) );
  NAND4_X1 U23999 ( .A1(n21685), .A2(n21686), .A3(n21687), .A4(n21688), .ZN(
        n21675) );
  NAND4_X1 U24000 ( .A1(n21677), .A2(n21678), .A3(n21679), .A4(n21680), .ZN(
        n21676) );
  OAI221_X1 U24001 ( .B1(n19221), .B2(n24807), .C1(n11829), .C2(n24799), .A(
        n21655), .ZN(n5042) );
  OAI21_X1 U24002 ( .B1(n21656), .B2(n21657), .A(n24795), .ZN(n21655) );
  NAND4_X1 U24003 ( .A1(n21666), .A2(n21667), .A3(n21668), .A4(n21669), .ZN(
        n21656) );
  NAND4_X1 U24004 ( .A1(n21658), .A2(n21659), .A3(n21660), .A4(n21661), .ZN(
        n21657) );
  OAI221_X1 U24005 ( .B1(n19220), .B2(n24807), .C1(n11830), .C2(n24799), .A(
        n21636), .ZN(n5043) );
  OAI21_X1 U24006 ( .B1(n21637), .B2(n21638), .A(n24795), .ZN(n21636) );
  NAND4_X1 U24007 ( .A1(n21647), .A2(n21648), .A3(n21649), .A4(n21650), .ZN(
        n21637) );
  NAND4_X1 U24008 ( .A1(n21639), .A2(n21640), .A3(n21641), .A4(n21642), .ZN(
        n21638) );
  OAI221_X1 U24009 ( .B1(n19219), .B2(n24808), .C1(n11831), .C2(n24799), .A(
        n21617), .ZN(n5044) );
  OAI21_X1 U24010 ( .B1(n21618), .B2(n21619), .A(n24796), .ZN(n21617) );
  NAND4_X1 U24011 ( .A1(n21628), .A2(n21629), .A3(n21630), .A4(n21631), .ZN(
        n21618) );
  NAND4_X1 U24012 ( .A1(n21620), .A2(n21621), .A3(n21622), .A4(n21623), .ZN(
        n21619) );
  OAI221_X1 U24013 ( .B1(n19218), .B2(n24808), .C1(n11832), .C2(n24799), .A(
        n21598), .ZN(n5045) );
  OAI21_X1 U24014 ( .B1(n21599), .B2(n21600), .A(n24796), .ZN(n21598) );
  NAND4_X1 U24015 ( .A1(n21609), .A2(n21610), .A3(n21611), .A4(n21612), .ZN(
        n21599) );
  NAND4_X1 U24016 ( .A1(n21601), .A2(n21602), .A3(n21603), .A4(n21604), .ZN(
        n21600) );
  OAI221_X1 U24017 ( .B1(n19217), .B2(n24808), .C1(n11833), .C2(n24799), .A(
        n21579), .ZN(n5046) );
  OAI21_X1 U24018 ( .B1(n21580), .B2(n21581), .A(n24796), .ZN(n21579) );
  NAND4_X1 U24019 ( .A1(n21590), .A2(n21591), .A3(n21592), .A4(n21593), .ZN(
        n21580) );
  NAND4_X1 U24020 ( .A1(n21582), .A2(n21583), .A3(n21584), .A4(n21585), .ZN(
        n21581) );
  OAI221_X1 U24021 ( .B1(n19216), .B2(n24808), .C1(n11834), .C2(n24798), .A(
        n21560), .ZN(n5047) );
  OAI21_X1 U24022 ( .B1(n21561), .B2(n21562), .A(n24796), .ZN(n21560) );
  NAND4_X1 U24023 ( .A1(n21571), .A2(n21572), .A3(n21573), .A4(n21574), .ZN(
        n21561) );
  NAND4_X1 U24024 ( .A1(n21563), .A2(n21564), .A3(n21565), .A4(n21566), .ZN(
        n21562) );
  OAI221_X1 U24025 ( .B1(n19215), .B2(n24808), .C1(n11835), .C2(n24798), .A(
        n21541), .ZN(n5048) );
  OAI21_X1 U24026 ( .B1(n21542), .B2(n21543), .A(n24796), .ZN(n21541) );
  NAND4_X1 U24027 ( .A1(n21552), .A2(n21553), .A3(n21554), .A4(n21555), .ZN(
        n21542) );
  NAND4_X1 U24028 ( .A1(n21544), .A2(n21545), .A3(n21546), .A4(n21547), .ZN(
        n21543) );
  OAI221_X1 U24029 ( .B1(n19214), .B2(n24808), .C1(n11836), .C2(n24798), .A(
        n21522), .ZN(n5049) );
  OAI21_X1 U24030 ( .B1(n21523), .B2(n21524), .A(n24796), .ZN(n21522) );
  NAND4_X1 U24031 ( .A1(n21533), .A2(n21534), .A3(n21535), .A4(n21536), .ZN(
        n21523) );
  NAND4_X1 U24032 ( .A1(n21525), .A2(n21526), .A3(n21527), .A4(n21528), .ZN(
        n21524) );
  OAI221_X1 U24033 ( .B1(n19213), .B2(n24808), .C1(n11837), .C2(n24798), .A(
        n21503), .ZN(n5050) );
  OAI21_X1 U24034 ( .B1(n21504), .B2(n21505), .A(n24796), .ZN(n21503) );
  NAND4_X1 U24035 ( .A1(n21514), .A2(n21515), .A3(n21516), .A4(n21517), .ZN(
        n21504) );
  NAND4_X1 U24036 ( .A1(n21506), .A2(n21507), .A3(n21508), .A4(n21509), .ZN(
        n21505) );
  OAI221_X1 U24037 ( .B1(n19212), .B2(n24808), .C1(n11838), .C2(n24798), .A(
        n21484), .ZN(n5051) );
  OAI21_X1 U24038 ( .B1(n21485), .B2(n21486), .A(n24796), .ZN(n21484) );
  NAND4_X1 U24039 ( .A1(n21495), .A2(n21496), .A3(n21497), .A4(n21498), .ZN(
        n21485) );
  NAND4_X1 U24040 ( .A1(n21487), .A2(n21488), .A3(n21489), .A4(n21490), .ZN(
        n21486) );
  OAI221_X1 U24041 ( .B1(n19211), .B2(n24808), .C1(n11839), .C2(n24798), .A(
        n21465), .ZN(n5052) );
  OAI21_X1 U24042 ( .B1(n21466), .B2(n21467), .A(n24796), .ZN(n21465) );
  NAND4_X1 U24043 ( .A1(n21476), .A2(n21477), .A3(n21478), .A4(n21479), .ZN(
        n21466) );
  NAND4_X1 U24044 ( .A1(n21468), .A2(n21469), .A3(n21470), .A4(n21471), .ZN(
        n21467) );
  OAI221_X1 U24045 ( .B1(n19210), .B2(n24808), .C1(n11840), .C2(n24798), .A(
        n21446), .ZN(n5053) );
  OAI21_X1 U24046 ( .B1(n21447), .B2(n21448), .A(n24796), .ZN(n21446) );
  NAND4_X1 U24047 ( .A1(n21457), .A2(n21458), .A3(n21459), .A4(n21460), .ZN(
        n21447) );
  NAND4_X1 U24048 ( .A1(n21449), .A2(n21450), .A3(n21451), .A4(n21452), .ZN(
        n21448) );
  OAI221_X1 U24049 ( .B1(n19209), .B2(n24808), .C1(n11841), .C2(n24798), .A(
        n21427), .ZN(n5054) );
  OAI21_X1 U24050 ( .B1(n21428), .B2(n21429), .A(n24796), .ZN(n21427) );
  NAND4_X1 U24051 ( .A1(n21438), .A2(n21439), .A3(n21440), .A4(n21441), .ZN(
        n21428) );
  NAND4_X1 U24052 ( .A1(n21430), .A2(n21431), .A3(n21432), .A4(n21433), .ZN(
        n21429) );
  OAI221_X1 U24053 ( .B1(n19208), .B2(n24808), .C1(n11842), .C2(n24798), .A(
        n21408), .ZN(n5055) );
  OAI21_X1 U24054 ( .B1(n21409), .B2(n21410), .A(n24796), .ZN(n21408) );
  NAND4_X1 U24055 ( .A1(n21419), .A2(n21420), .A3(n21421), .A4(n21422), .ZN(
        n21409) );
  NAND4_X1 U24056 ( .A1(n21411), .A2(n21412), .A3(n21413), .A4(n21414), .ZN(
        n21410) );
  NAND4_X1 U24057 ( .A1(n23008), .A2(n23009), .A3(n23010), .A4(n23011), .ZN(
        n4972) );
  AOI221_X1 U24058 ( .B1(n24441), .B2(n24332), .C1(n24435), .C2(n19877), .A(
        n23024), .ZN(n23009) );
  AOI221_X1 U24059 ( .B1(n24417), .B2(n19483), .C1(n24410), .C2(OUT2[40]), .A(
        n23025), .ZN(n23008) );
  NOR4_X1 U24060 ( .A1(n23020), .A2(n23021), .A3(n23022), .A4(n23023), .ZN(
        n23010) );
  NAND4_X1 U24061 ( .A1(n22990), .A2(n22991), .A3(n22992), .A4(n22993), .ZN(
        n4973) );
  AOI221_X1 U24062 ( .B1(n24441), .B2(n24333), .C1(n24435), .C2(n19876), .A(
        n23006), .ZN(n22991) );
  AOI221_X1 U24063 ( .B1(n24417), .B2(n19482), .C1(n24409), .C2(OUT2[41]), .A(
        n23007), .ZN(n22990) );
  NOR4_X1 U24064 ( .A1(n23002), .A2(n23003), .A3(n23004), .A4(n23005), .ZN(
        n22992) );
  NAND4_X1 U24065 ( .A1(n22972), .A2(n22973), .A3(n22974), .A4(n22975), .ZN(
        n4974) );
  AOI221_X1 U24066 ( .B1(n24441), .B2(n24334), .C1(n24435), .C2(n19875), .A(
        n22988), .ZN(n22973) );
  AOI221_X1 U24067 ( .B1(n24417), .B2(n19481), .C1(n24409), .C2(OUT2[42]), .A(
        n22989), .ZN(n22972) );
  NOR4_X1 U24068 ( .A1(n22984), .A2(n22985), .A3(n22986), .A4(n22987), .ZN(
        n22974) );
  NAND4_X1 U24069 ( .A1(n22954), .A2(n22955), .A3(n22956), .A4(n22957), .ZN(
        n4975) );
  AOI221_X1 U24070 ( .B1(n24441), .B2(n24335), .C1(n24435), .C2(n19874), .A(
        n22970), .ZN(n22955) );
  AOI221_X1 U24071 ( .B1(n24417), .B2(n19480), .C1(n24409), .C2(OUT2[43]), .A(
        n22971), .ZN(n22954) );
  NOR4_X1 U24072 ( .A1(n22966), .A2(n22967), .A3(n22968), .A4(n22969), .ZN(
        n22956) );
  NAND4_X1 U24073 ( .A1(n22936), .A2(n22937), .A3(n22938), .A4(n22939), .ZN(
        n4976) );
  AOI221_X1 U24074 ( .B1(n24441), .B2(n24336), .C1(n24435), .C2(n19873), .A(
        n22952), .ZN(n22937) );
  AOI221_X1 U24075 ( .B1(n24417), .B2(n19479), .C1(n24409), .C2(OUT2[44]), .A(
        n22953), .ZN(n22936) );
  NOR4_X1 U24076 ( .A1(n22948), .A2(n22949), .A3(n22950), .A4(n22951), .ZN(
        n22938) );
  NAND4_X1 U24077 ( .A1(n22918), .A2(n22919), .A3(n22920), .A4(n22921), .ZN(
        n4977) );
  AOI221_X1 U24078 ( .B1(n24441), .B2(n24337), .C1(n24435), .C2(n19872), .A(
        n22934), .ZN(n22919) );
  AOI221_X1 U24079 ( .B1(n24417), .B2(n19478), .C1(n24409), .C2(OUT2[45]), .A(
        n22935), .ZN(n22918) );
  NOR4_X1 U24080 ( .A1(n22930), .A2(n22931), .A3(n22932), .A4(n22933), .ZN(
        n22920) );
  NAND4_X1 U24081 ( .A1(n22900), .A2(n22901), .A3(n22902), .A4(n22903), .ZN(
        n4978) );
  AOI221_X1 U24082 ( .B1(n24441), .B2(n24338), .C1(n24435), .C2(n19871), .A(
        n22916), .ZN(n22901) );
  AOI221_X1 U24083 ( .B1(n24417), .B2(n19477), .C1(n24409), .C2(OUT2[46]), .A(
        n22917), .ZN(n22900) );
  NOR4_X1 U24084 ( .A1(n22912), .A2(n22913), .A3(n22914), .A4(n22915), .ZN(
        n22902) );
  NAND4_X1 U24085 ( .A1(n22882), .A2(n22883), .A3(n22884), .A4(n22885), .ZN(
        n4979) );
  AOI221_X1 U24086 ( .B1(n24441), .B2(n24339), .C1(n24435), .C2(n19870), .A(
        n22898), .ZN(n22883) );
  AOI221_X1 U24087 ( .B1(n24417), .B2(n19476), .C1(n24409), .C2(OUT2[47]), .A(
        n22899), .ZN(n22882) );
  NOR4_X1 U24088 ( .A1(n22894), .A2(n22895), .A3(n22896), .A4(n22897), .ZN(
        n22884) );
  NAND4_X1 U24089 ( .A1(n22864), .A2(n22865), .A3(n22866), .A4(n22867), .ZN(
        n4980) );
  AOI221_X1 U24090 ( .B1(n24442), .B2(n24340), .C1(n24436), .C2(n19869), .A(
        n22880), .ZN(n22865) );
  AOI221_X1 U24091 ( .B1(n24418), .B2(n19475), .C1(n24409), .C2(OUT2[48]), .A(
        n22881), .ZN(n22864) );
  NOR4_X1 U24092 ( .A1(n22876), .A2(n22877), .A3(n22878), .A4(n22879), .ZN(
        n22866) );
  NAND4_X1 U24093 ( .A1(n22846), .A2(n22847), .A3(n22848), .A4(n22849), .ZN(
        n4981) );
  AOI221_X1 U24094 ( .B1(n24442), .B2(n24341), .C1(n24436), .C2(n19868), .A(
        n22862), .ZN(n22847) );
  AOI221_X1 U24095 ( .B1(n24418), .B2(n19474), .C1(n24409), .C2(OUT2[49]), .A(
        n22863), .ZN(n22846) );
  NOR4_X1 U24096 ( .A1(n22858), .A2(n22859), .A3(n22860), .A4(n22861), .ZN(
        n22848) );
  NAND4_X1 U24097 ( .A1(n22828), .A2(n22829), .A3(n22830), .A4(n22831), .ZN(
        n4982) );
  AOI221_X1 U24098 ( .B1(n24442), .B2(n24342), .C1(n24436), .C2(n19867), .A(
        n22844), .ZN(n22829) );
  AOI221_X1 U24099 ( .B1(n24418), .B2(n19473), .C1(n24409), .C2(OUT2[50]), .A(
        n22845), .ZN(n22828) );
  NOR4_X1 U24100 ( .A1(n22840), .A2(n22841), .A3(n22842), .A4(n22843), .ZN(
        n22830) );
  NAND4_X1 U24101 ( .A1(n22810), .A2(n22811), .A3(n22812), .A4(n22813), .ZN(
        n4983) );
  AOI221_X1 U24102 ( .B1(n24442), .B2(n24343), .C1(n24436), .C2(n19866), .A(
        n22826), .ZN(n22811) );
  AOI221_X1 U24103 ( .B1(n24418), .B2(n19472), .C1(n24409), .C2(OUT2[51]), .A(
        n22827), .ZN(n22810) );
  NOR4_X1 U24104 ( .A1(n22822), .A2(n22823), .A3(n22824), .A4(n22825), .ZN(
        n22812) );
  NAND4_X1 U24105 ( .A1(n22792), .A2(n22793), .A3(n22794), .A4(n22795), .ZN(
        n4984) );
  AOI221_X1 U24106 ( .B1(n24442), .B2(n24344), .C1(n24436), .C2(n19865), .A(
        n22808), .ZN(n22793) );
  AOI221_X1 U24107 ( .B1(n24418), .B2(n19471), .C1(n24409), .C2(OUT2[52]), .A(
        n22809), .ZN(n22792) );
  NOR4_X1 U24108 ( .A1(n22804), .A2(n22805), .A3(n22806), .A4(n22807), .ZN(
        n22794) );
  NAND4_X1 U24109 ( .A1(n22774), .A2(n22775), .A3(n22776), .A4(n22777), .ZN(
        n4985) );
  AOI221_X1 U24110 ( .B1(n24442), .B2(n24345), .C1(n24436), .C2(n19864), .A(
        n22790), .ZN(n22775) );
  AOI221_X1 U24111 ( .B1(n24418), .B2(n19470), .C1(n24408), .C2(OUT2[53]), .A(
        n22791), .ZN(n22774) );
  NOR4_X1 U24112 ( .A1(n22786), .A2(n22787), .A3(n22788), .A4(n22789), .ZN(
        n22776) );
  NAND4_X1 U24113 ( .A1(n22756), .A2(n22757), .A3(n22758), .A4(n22759), .ZN(
        n4986) );
  AOI221_X1 U24114 ( .B1(n24442), .B2(n24346), .C1(n24436), .C2(n19863), .A(
        n22772), .ZN(n22757) );
  AOI221_X1 U24115 ( .B1(n24418), .B2(n19469), .C1(n24408), .C2(OUT2[54]), .A(
        n22773), .ZN(n22756) );
  NOR4_X1 U24116 ( .A1(n22768), .A2(n22769), .A3(n22770), .A4(n22771), .ZN(
        n22758) );
  NAND4_X1 U24117 ( .A1(n22738), .A2(n22739), .A3(n22740), .A4(n22741), .ZN(
        n4987) );
  AOI221_X1 U24118 ( .B1(n24442), .B2(n24347), .C1(n24436), .C2(n19862), .A(
        n22754), .ZN(n22739) );
  AOI221_X1 U24119 ( .B1(n24418), .B2(n19468), .C1(n24408), .C2(OUT2[55]), .A(
        n22755), .ZN(n22738) );
  NOR4_X1 U24120 ( .A1(n22750), .A2(n22751), .A3(n22752), .A4(n22753), .ZN(
        n22740) );
  NAND4_X1 U24121 ( .A1(n22720), .A2(n22721), .A3(n22722), .A4(n22723), .ZN(
        n4988) );
  AOI221_X1 U24122 ( .B1(n24442), .B2(n24348), .C1(n24436), .C2(n19861), .A(
        n22736), .ZN(n22721) );
  AOI221_X1 U24123 ( .B1(n24418), .B2(n19467), .C1(n24408), .C2(OUT2[56]), .A(
        n22737), .ZN(n22720) );
  NOR4_X1 U24124 ( .A1(n22732), .A2(n22733), .A3(n22734), .A4(n22735), .ZN(
        n22722) );
  NAND4_X1 U24125 ( .A1(n22702), .A2(n22703), .A3(n22704), .A4(n22705), .ZN(
        n4989) );
  AOI221_X1 U24126 ( .B1(n24442), .B2(n24349), .C1(n24436), .C2(n19860), .A(
        n22718), .ZN(n22703) );
  AOI221_X1 U24127 ( .B1(n24418), .B2(n19466), .C1(n24408), .C2(OUT2[57]), .A(
        n22719), .ZN(n22702) );
  NOR4_X1 U24128 ( .A1(n22714), .A2(n22715), .A3(n22716), .A4(n22717), .ZN(
        n22704) );
  NAND4_X1 U24129 ( .A1(n22684), .A2(n22685), .A3(n22686), .A4(n22687), .ZN(
        n4990) );
  AOI221_X1 U24130 ( .B1(n24442), .B2(n24350), .C1(n24436), .C2(n19859), .A(
        n22700), .ZN(n22685) );
  AOI221_X1 U24131 ( .B1(n24418), .B2(n19465), .C1(n24408), .C2(OUT2[58]), .A(
        n22701), .ZN(n22684) );
  NOR4_X1 U24132 ( .A1(n22696), .A2(n22697), .A3(n22698), .A4(n22699), .ZN(
        n22686) );
  NAND4_X1 U24133 ( .A1(n22666), .A2(n22667), .A3(n22668), .A4(n22669), .ZN(
        n4991) );
  AOI221_X1 U24134 ( .B1(n24442), .B2(n24351), .C1(n24436), .C2(n19858), .A(
        n22682), .ZN(n22667) );
  AOI221_X1 U24135 ( .B1(n24418), .B2(n19464), .C1(n24408), .C2(OUT2[59]), .A(
        n22683), .ZN(n22666) );
  NOR4_X1 U24136 ( .A1(n22678), .A2(n22679), .A3(n22680), .A4(n22681), .ZN(
        n22668) );
  NAND4_X1 U24137 ( .A1(n22648), .A2(n22649), .A3(n22650), .A4(n22651), .ZN(
        n4992) );
  AOI221_X1 U24138 ( .B1(n24443), .B2(n24352), .C1(n24437), .C2(n19809), .A(
        n22664), .ZN(n22649) );
  AOI221_X1 U24139 ( .B1(n24419), .B2(n19463), .C1(n24408), .C2(OUT2[60]), .A(
        n22665), .ZN(n22648) );
  NOR4_X1 U24140 ( .A1(n22660), .A2(n22661), .A3(n22662), .A4(n22663), .ZN(
        n22650) );
  NAND4_X1 U24141 ( .A1(n22630), .A2(n22631), .A3(n22632), .A4(n22633), .ZN(
        n4993) );
  AOI221_X1 U24142 ( .B1(n24443), .B2(n24353), .C1(n24437), .C2(n19808), .A(
        n22646), .ZN(n22631) );
  AOI221_X1 U24143 ( .B1(n24419), .B2(n19462), .C1(n24408), .C2(OUT2[61]), .A(
        n22647), .ZN(n22630) );
  NOR4_X1 U24144 ( .A1(n22642), .A2(n22643), .A3(n22644), .A4(n22645), .ZN(
        n22632) );
  NAND4_X1 U24145 ( .A1(n22612), .A2(n22613), .A3(n22614), .A4(n22615), .ZN(
        n4994) );
  AOI221_X1 U24146 ( .B1(n24443), .B2(n24354), .C1(n24437), .C2(n19807), .A(
        n22628), .ZN(n22613) );
  AOI221_X1 U24147 ( .B1(n24419), .B2(n19461), .C1(n24408), .C2(OUT2[62]), .A(
        n22629), .ZN(n22612) );
  NOR4_X1 U24148 ( .A1(n22624), .A2(n22625), .A3(n22626), .A4(n22627), .ZN(
        n22614) );
  NAND4_X1 U24149 ( .A1(n22560), .A2(n22561), .A3(n22562), .A4(n22563), .ZN(
        n4995) );
  AOI221_X1 U24150 ( .B1(n24443), .B2(n24355), .C1(n24437), .C2(n19806), .A(
        n22604), .ZN(n22561) );
  AOI221_X1 U24151 ( .B1(n24419), .B2(n19460), .C1(n24410), .C2(OUT2[63]), .A(
        n22609), .ZN(n22560) );
  NOR4_X1 U24152 ( .A1(n22589), .A2(n22590), .A3(n22591), .A4(n22592), .ZN(
        n22562) );
  NAND4_X1 U24153 ( .A1(n23728), .A2(n23729), .A3(n23730), .A4(n23731), .ZN(
        n4932) );
  AOI221_X1 U24154 ( .B1(n24438), .B2(n24356), .C1(n24432), .C2(n20049), .A(
        n23762), .ZN(n23729) );
  AOI221_X1 U24155 ( .B1(n24414), .B2(n19523), .C1(n24408), .C2(OUT2[0]), .A(
        n23763), .ZN(n23728) );
  NOR4_X1 U24156 ( .A1(n23750), .A2(n23751), .A3(n23752), .A4(n23753), .ZN(
        n23730) );
  NAND4_X1 U24157 ( .A1(n23710), .A2(n23711), .A3(n23712), .A4(n23713), .ZN(
        n4933) );
  AOI221_X1 U24158 ( .B1(n24438), .B2(n24357), .C1(n24432), .C2(n20048), .A(
        n23726), .ZN(n23711) );
  AOI221_X1 U24159 ( .B1(n24414), .B2(n19522), .C1(n24413), .C2(OUT2[1]), .A(
        n23727), .ZN(n23710) );
  NOR4_X1 U24160 ( .A1(n23722), .A2(n23723), .A3(n23724), .A4(n23725), .ZN(
        n23712) );
  NAND4_X1 U24161 ( .A1(n23692), .A2(n23693), .A3(n23694), .A4(n23695), .ZN(
        n4934) );
  AOI221_X1 U24162 ( .B1(n24438), .B2(n24358), .C1(n24432), .C2(n20047), .A(
        n23708), .ZN(n23693) );
  AOI221_X1 U24163 ( .B1(n24414), .B2(n19521), .C1(n24413), .C2(OUT2[2]), .A(
        n23709), .ZN(n23692) );
  NOR4_X1 U24164 ( .A1(n23704), .A2(n23705), .A3(n23706), .A4(n23707), .ZN(
        n23694) );
  NAND4_X1 U24165 ( .A1(n23674), .A2(n23675), .A3(n23676), .A4(n23677), .ZN(
        n4935) );
  AOI221_X1 U24166 ( .B1(n24438), .B2(n24359), .C1(n24432), .C2(n20046), .A(
        n23690), .ZN(n23675) );
  AOI221_X1 U24167 ( .B1(n24414), .B2(n19520), .C1(n24413), .C2(OUT2[3]), .A(
        n23691), .ZN(n23674) );
  NOR4_X1 U24168 ( .A1(n23686), .A2(n23687), .A3(n23688), .A4(n23689), .ZN(
        n23676) );
  NAND4_X1 U24169 ( .A1(n23656), .A2(n23657), .A3(n23658), .A4(n23659), .ZN(
        n4936) );
  AOI221_X1 U24170 ( .B1(n24438), .B2(n24360), .C1(n24432), .C2(n20045), .A(
        n23672), .ZN(n23657) );
  AOI221_X1 U24171 ( .B1(n24414), .B2(n19519), .C1(n24413), .C2(OUT2[4]), .A(
        n23673), .ZN(n23656) );
  NOR4_X1 U24172 ( .A1(n23668), .A2(n23669), .A3(n23670), .A4(n23671), .ZN(
        n23658) );
  NAND4_X1 U24173 ( .A1(n23638), .A2(n23639), .A3(n23640), .A4(n23641), .ZN(
        n4937) );
  AOI221_X1 U24174 ( .B1(n24438), .B2(n24361), .C1(n24432), .C2(n20044), .A(
        n23654), .ZN(n23639) );
  AOI221_X1 U24175 ( .B1(n24414), .B2(n19518), .C1(n24413), .C2(OUT2[5]), .A(
        n23655), .ZN(n23638) );
  NOR4_X1 U24176 ( .A1(n23650), .A2(n23651), .A3(n23652), .A4(n23653), .ZN(
        n23640) );
  NAND4_X1 U24177 ( .A1(n23620), .A2(n23621), .A3(n23622), .A4(n23623), .ZN(
        n4938) );
  AOI221_X1 U24178 ( .B1(n24438), .B2(n24362), .C1(n24432), .C2(n20043), .A(
        n23636), .ZN(n23621) );
  AOI221_X1 U24179 ( .B1(n24414), .B2(n19517), .C1(n24412), .C2(OUT2[6]), .A(
        n23637), .ZN(n23620) );
  NOR4_X1 U24180 ( .A1(n23632), .A2(n23633), .A3(n23634), .A4(n23635), .ZN(
        n23622) );
  NAND4_X1 U24181 ( .A1(n23602), .A2(n23603), .A3(n23604), .A4(n23605), .ZN(
        n4939) );
  AOI221_X1 U24182 ( .B1(n24438), .B2(n24363), .C1(n24432), .C2(n20042), .A(
        n23618), .ZN(n23603) );
  AOI221_X1 U24183 ( .B1(n24414), .B2(n19516), .C1(n24412), .C2(OUT2[7]), .A(
        n23619), .ZN(n23602) );
  NOR4_X1 U24184 ( .A1(n23614), .A2(n23615), .A3(n23616), .A4(n23617), .ZN(
        n23604) );
  NAND4_X1 U24185 ( .A1(n23584), .A2(n23585), .A3(n23586), .A4(n23587), .ZN(
        n4940) );
  AOI221_X1 U24186 ( .B1(n24438), .B2(n24364), .C1(n24432), .C2(n20041), .A(
        n23600), .ZN(n23585) );
  AOI221_X1 U24187 ( .B1(n24414), .B2(n19515), .C1(n24412), .C2(OUT2[8]), .A(
        n23601), .ZN(n23584) );
  NOR4_X1 U24188 ( .A1(n23596), .A2(n23597), .A3(n23598), .A4(n23599), .ZN(
        n23586) );
  NAND4_X1 U24189 ( .A1(n23566), .A2(n23567), .A3(n23568), .A4(n23569), .ZN(
        n4941) );
  AOI221_X1 U24190 ( .B1(n24438), .B2(n24365), .C1(n24432), .C2(n20040), .A(
        n23582), .ZN(n23567) );
  AOI221_X1 U24191 ( .B1(n24414), .B2(n19514), .C1(n24412), .C2(OUT2[9]), .A(
        n23583), .ZN(n23566) );
  NOR4_X1 U24192 ( .A1(n23578), .A2(n23579), .A3(n23580), .A4(n23581), .ZN(
        n23568) );
  NAND4_X1 U24193 ( .A1(n23548), .A2(n23549), .A3(n23550), .A4(n23551), .ZN(
        n4942) );
  AOI221_X1 U24194 ( .B1(n24438), .B2(n24366), .C1(n24432), .C2(n20039), .A(
        n23564), .ZN(n23549) );
  AOI221_X1 U24195 ( .B1(n24414), .B2(n19513), .C1(n24412), .C2(OUT2[10]), .A(
        n23565), .ZN(n23548) );
  NOR4_X1 U24196 ( .A1(n23560), .A2(n23561), .A3(n23562), .A4(n23563), .ZN(
        n23550) );
  NAND4_X1 U24197 ( .A1(n23530), .A2(n23531), .A3(n23532), .A4(n23533), .ZN(
        n4943) );
  AOI221_X1 U24198 ( .B1(n24438), .B2(n24367), .C1(n24432), .C2(n20038), .A(
        n23546), .ZN(n23531) );
  AOI221_X1 U24199 ( .B1(n24414), .B2(n19512), .C1(n24412), .C2(OUT2[11]), .A(
        n23547), .ZN(n23530) );
  NOR4_X1 U24200 ( .A1(n23542), .A2(n23543), .A3(n23544), .A4(n23545), .ZN(
        n23532) );
  NAND4_X1 U24201 ( .A1(n23512), .A2(n23513), .A3(n23514), .A4(n23515), .ZN(
        n4944) );
  AOI221_X1 U24202 ( .B1(n24439), .B2(n24368), .C1(n24433), .C2(n20037), .A(
        n23528), .ZN(n23513) );
  AOI221_X1 U24203 ( .B1(n24415), .B2(n19511), .C1(n24412), .C2(OUT2[12]), .A(
        n23529), .ZN(n23512) );
  NOR4_X1 U24204 ( .A1(n23524), .A2(n23525), .A3(n23526), .A4(n23527), .ZN(
        n23514) );
  NAND4_X1 U24205 ( .A1(n23494), .A2(n23495), .A3(n23496), .A4(n23497), .ZN(
        n4945) );
  AOI221_X1 U24206 ( .B1(n24439), .B2(n24369), .C1(n24433), .C2(n20036), .A(
        n23510), .ZN(n23495) );
  AOI221_X1 U24207 ( .B1(n24415), .B2(n19510), .C1(n24412), .C2(OUT2[13]), .A(
        n23511), .ZN(n23494) );
  NOR4_X1 U24208 ( .A1(n23506), .A2(n23507), .A3(n23508), .A4(n23509), .ZN(
        n23496) );
  NAND4_X1 U24209 ( .A1(n23476), .A2(n23477), .A3(n23478), .A4(n23479), .ZN(
        n4946) );
  AOI221_X1 U24210 ( .B1(n24439), .B2(n24370), .C1(n24433), .C2(n20035), .A(
        n23492), .ZN(n23477) );
  AOI221_X1 U24211 ( .B1(n24415), .B2(n19509), .C1(n24412), .C2(OUT2[14]), .A(
        n23493), .ZN(n23476) );
  NOR4_X1 U24212 ( .A1(n23488), .A2(n23489), .A3(n23490), .A4(n23491), .ZN(
        n23478) );
  NAND4_X1 U24213 ( .A1(n23458), .A2(n23459), .A3(n23460), .A4(n23461), .ZN(
        n4947) );
  AOI221_X1 U24214 ( .B1(n24439), .B2(n24371), .C1(n24433), .C2(n20034), .A(
        n23474), .ZN(n23459) );
  AOI221_X1 U24215 ( .B1(n24415), .B2(n19508), .C1(n24412), .C2(OUT2[15]), .A(
        n23475), .ZN(n23458) );
  NOR4_X1 U24216 ( .A1(n23470), .A2(n23471), .A3(n23472), .A4(n23473), .ZN(
        n23460) );
  NAND4_X1 U24217 ( .A1(n23440), .A2(n23441), .A3(n23442), .A4(n23443), .ZN(
        n4948) );
  AOI221_X1 U24218 ( .B1(n24439), .B2(n24372), .C1(n24433), .C2(n20033), .A(
        n23456), .ZN(n23441) );
  AOI221_X1 U24219 ( .B1(n24415), .B2(n19507), .C1(n24412), .C2(OUT2[16]), .A(
        n23457), .ZN(n23440) );
  NOR4_X1 U24220 ( .A1(n23452), .A2(n23453), .A3(n23454), .A4(n23455), .ZN(
        n23442) );
  NAND4_X1 U24221 ( .A1(n23422), .A2(n23423), .A3(n23424), .A4(n23425), .ZN(
        n4949) );
  AOI221_X1 U24222 ( .B1(n24439), .B2(n24373), .C1(n24433), .C2(n20032), .A(
        n23438), .ZN(n23423) );
  AOI221_X1 U24223 ( .B1(n24415), .B2(n19506), .C1(n24412), .C2(OUT2[17]), .A(
        n23439), .ZN(n23422) );
  NOR4_X1 U24224 ( .A1(n23434), .A2(n23435), .A3(n23436), .A4(n23437), .ZN(
        n23424) );
  NAND4_X1 U24225 ( .A1(n23404), .A2(n23405), .A3(n23406), .A4(n23407), .ZN(
        n4950) );
  AOI221_X1 U24226 ( .B1(n24439), .B2(n24374), .C1(n24433), .C2(n20031), .A(
        n23420), .ZN(n23405) );
  AOI221_X1 U24227 ( .B1(n24415), .B2(n19505), .C1(n24411), .C2(OUT2[18]), .A(
        n23421), .ZN(n23404) );
  NOR4_X1 U24228 ( .A1(n23416), .A2(n23417), .A3(n23418), .A4(n23419), .ZN(
        n23406) );
  NAND4_X1 U24229 ( .A1(n23386), .A2(n23387), .A3(n23388), .A4(n23389), .ZN(
        n4951) );
  AOI221_X1 U24230 ( .B1(n24439), .B2(n24375), .C1(n24433), .C2(n20030), .A(
        n23402), .ZN(n23387) );
  AOI221_X1 U24231 ( .B1(n24415), .B2(n19504), .C1(n24411), .C2(OUT2[19]), .A(
        n23403), .ZN(n23386) );
  NOR4_X1 U24232 ( .A1(n23398), .A2(n23399), .A3(n23400), .A4(n23401), .ZN(
        n23388) );
  NAND4_X1 U24233 ( .A1(n23368), .A2(n23369), .A3(n23370), .A4(n23371), .ZN(
        n4952) );
  AOI221_X1 U24234 ( .B1(n24439), .B2(n24376), .C1(n24433), .C2(n20029), .A(
        n23384), .ZN(n23369) );
  AOI221_X1 U24235 ( .B1(n24415), .B2(n19503), .C1(n24411), .C2(OUT2[20]), .A(
        n23385), .ZN(n23368) );
  NOR4_X1 U24236 ( .A1(n23380), .A2(n23381), .A3(n23382), .A4(n23383), .ZN(
        n23370) );
  NAND4_X1 U24237 ( .A1(n23350), .A2(n23351), .A3(n23352), .A4(n23353), .ZN(
        n4953) );
  AOI221_X1 U24238 ( .B1(n24439), .B2(n24377), .C1(n24433), .C2(n20028), .A(
        n23366), .ZN(n23351) );
  AOI221_X1 U24239 ( .B1(n24415), .B2(n19502), .C1(n24411), .C2(OUT2[21]), .A(
        n23367), .ZN(n23350) );
  NOR4_X1 U24240 ( .A1(n23362), .A2(n23363), .A3(n23364), .A4(n23365), .ZN(
        n23352) );
  NAND4_X1 U24241 ( .A1(n23332), .A2(n23333), .A3(n23334), .A4(n23335), .ZN(
        n4954) );
  AOI221_X1 U24242 ( .B1(n24439), .B2(n24378), .C1(n24433), .C2(n20027), .A(
        n23348), .ZN(n23333) );
  AOI221_X1 U24243 ( .B1(n24415), .B2(n19501), .C1(n24411), .C2(OUT2[22]), .A(
        n23349), .ZN(n23332) );
  NOR4_X1 U24244 ( .A1(n23344), .A2(n23345), .A3(n23346), .A4(n23347), .ZN(
        n23334) );
  NAND4_X1 U24245 ( .A1(n23314), .A2(n23315), .A3(n23316), .A4(n23317), .ZN(
        n4955) );
  AOI221_X1 U24246 ( .B1(n24439), .B2(n24379), .C1(n24433), .C2(n20026), .A(
        n23330), .ZN(n23315) );
  AOI221_X1 U24247 ( .B1(n24415), .B2(n19500), .C1(n24411), .C2(OUT2[23]), .A(
        n23331), .ZN(n23314) );
  NOR4_X1 U24248 ( .A1(n23326), .A2(n23327), .A3(n23328), .A4(n23329), .ZN(
        n23316) );
  NAND4_X1 U24249 ( .A1(n23296), .A2(n23297), .A3(n23298), .A4(n23299), .ZN(
        n4956) );
  AOI221_X1 U24250 ( .B1(n24440), .B2(n24380), .C1(n24434), .C2(n19893), .A(
        n23312), .ZN(n23297) );
  AOI221_X1 U24251 ( .B1(n24416), .B2(n19499), .C1(n24411), .C2(OUT2[24]), .A(
        n23313), .ZN(n23296) );
  NOR4_X1 U24252 ( .A1(n23308), .A2(n23309), .A3(n23310), .A4(n23311), .ZN(
        n23298) );
  NAND4_X1 U24253 ( .A1(n23278), .A2(n23279), .A3(n23280), .A4(n23281), .ZN(
        n4957) );
  AOI221_X1 U24254 ( .B1(n24440), .B2(n24381), .C1(n24434), .C2(n19892), .A(
        n23294), .ZN(n23279) );
  AOI221_X1 U24255 ( .B1(n24416), .B2(n19498), .C1(n24411), .C2(OUT2[25]), .A(
        n23295), .ZN(n23278) );
  NOR4_X1 U24256 ( .A1(n23290), .A2(n23291), .A3(n23292), .A4(n23293), .ZN(
        n23280) );
  NAND4_X1 U24257 ( .A1(n23260), .A2(n23261), .A3(n23262), .A4(n23263), .ZN(
        n4958) );
  AOI221_X1 U24258 ( .B1(n24440), .B2(n24382), .C1(n24434), .C2(n19891), .A(
        n23276), .ZN(n23261) );
  AOI221_X1 U24259 ( .B1(n24416), .B2(n19497), .C1(n24411), .C2(OUT2[26]), .A(
        n23277), .ZN(n23260) );
  NOR4_X1 U24260 ( .A1(n23272), .A2(n23273), .A3(n23274), .A4(n23275), .ZN(
        n23262) );
  NAND4_X1 U24261 ( .A1(n23242), .A2(n23243), .A3(n23244), .A4(n23245), .ZN(
        n4959) );
  AOI221_X1 U24262 ( .B1(n24440), .B2(n24383), .C1(n24434), .C2(n19890), .A(
        n23258), .ZN(n23243) );
  AOI221_X1 U24263 ( .B1(n24416), .B2(n19496), .C1(n24411), .C2(OUT2[27]), .A(
        n23259), .ZN(n23242) );
  NOR4_X1 U24264 ( .A1(n23254), .A2(n23255), .A3(n23256), .A4(n23257), .ZN(
        n23244) );
  NAND4_X1 U24265 ( .A1(n23224), .A2(n23225), .A3(n23226), .A4(n23227), .ZN(
        n4960) );
  AOI221_X1 U24266 ( .B1(n24440), .B2(n24384), .C1(n24434), .C2(n19889), .A(
        n23240), .ZN(n23225) );
  AOI221_X1 U24267 ( .B1(n24416), .B2(n19495), .C1(n24411), .C2(OUT2[28]), .A(
        n23241), .ZN(n23224) );
  NOR4_X1 U24268 ( .A1(n23236), .A2(n23237), .A3(n23238), .A4(n23239), .ZN(
        n23226) );
  NAND4_X1 U24269 ( .A1(n23206), .A2(n23207), .A3(n23208), .A4(n23209), .ZN(
        n4961) );
  AOI221_X1 U24270 ( .B1(n24440), .B2(n24385), .C1(n24434), .C2(n19888), .A(
        n23222), .ZN(n23207) );
  AOI221_X1 U24271 ( .B1(n24416), .B2(n19494), .C1(n24411), .C2(OUT2[29]), .A(
        n23223), .ZN(n23206) );
  NOR4_X1 U24272 ( .A1(n23218), .A2(n23219), .A3(n23220), .A4(n23221), .ZN(
        n23208) );
  NAND4_X1 U24273 ( .A1(n23188), .A2(n23189), .A3(n23190), .A4(n23191), .ZN(
        n4962) );
  AOI221_X1 U24274 ( .B1(n24440), .B2(n24386), .C1(n24434), .C2(n19887), .A(
        n23204), .ZN(n23189) );
  AOI221_X1 U24275 ( .B1(n24416), .B2(n19493), .C1(n24410), .C2(OUT2[30]), .A(
        n23205), .ZN(n23188) );
  NOR4_X1 U24276 ( .A1(n23200), .A2(n23201), .A3(n23202), .A4(n23203), .ZN(
        n23190) );
  NAND4_X1 U24277 ( .A1(n23170), .A2(n23171), .A3(n23172), .A4(n23173), .ZN(
        n4963) );
  AOI221_X1 U24278 ( .B1(n24440), .B2(n24387), .C1(n24434), .C2(n19886), .A(
        n23186), .ZN(n23171) );
  AOI221_X1 U24279 ( .B1(n24416), .B2(n19492), .C1(n24410), .C2(OUT2[31]), .A(
        n23187), .ZN(n23170) );
  NOR4_X1 U24280 ( .A1(n23182), .A2(n23183), .A3(n23184), .A4(n23185), .ZN(
        n23172) );
  NAND4_X1 U24281 ( .A1(n23152), .A2(n23153), .A3(n23154), .A4(n23155), .ZN(
        n4964) );
  AOI221_X1 U24282 ( .B1(n24440), .B2(n24388), .C1(n24434), .C2(n19885), .A(
        n23168), .ZN(n23153) );
  AOI221_X1 U24283 ( .B1(n24416), .B2(n19491), .C1(n24410), .C2(OUT2[32]), .A(
        n23169), .ZN(n23152) );
  NOR4_X1 U24284 ( .A1(n23164), .A2(n23165), .A3(n23166), .A4(n23167), .ZN(
        n23154) );
  NAND4_X1 U24285 ( .A1(n23134), .A2(n23135), .A3(n23136), .A4(n23137), .ZN(
        n4965) );
  AOI221_X1 U24286 ( .B1(n24440), .B2(n24389), .C1(n24434), .C2(n19884), .A(
        n23150), .ZN(n23135) );
  AOI221_X1 U24287 ( .B1(n24416), .B2(n19490), .C1(n24410), .C2(OUT2[33]), .A(
        n23151), .ZN(n23134) );
  NOR4_X1 U24288 ( .A1(n23146), .A2(n23147), .A3(n23148), .A4(n23149), .ZN(
        n23136) );
  NAND4_X1 U24289 ( .A1(n23116), .A2(n23117), .A3(n23118), .A4(n23119), .ZN(
        n4966) );
  AOI221_X1 U24290 ( .B1(n24440), .B2(n24390), .C1(n24434), .C2(n19883), .A(
        n23132), .ZN(n23117) );
  AOI221_X1 U24291 ( .B1(n24416), .B2(n19489), .C1(n24410), .C2(OUT2[34]), .A(
        n23133), .ZN(n23116) );
  NOR4_X1 U24292 ( .A1(n23128), .A2(n23129), .A3(n23130), .A4(n23131), .ZN(
        n23118) );
  NAND4_X1 U24293 ( .A1(n23098), .A2(n23099), .A3(n23100), .A4(n23101), .ZN(
        n4967) );
  AOI221_X1 U24294 ( .B1(n24440), .B2(n24391), .C1(n24434), .C2(n19882), .A(
        n23114), .ZN(n23099) );
  AOI221_X1 U24295 ( .B1(n24416), .B2(n19488), .C1(n24410), .C2(OUT2[35]), .A(
        n23115), .ZN(n23098) );
  NOR4_X1 U24296 ( .A1(n23110), .A2(n23111), .A3(n23112), .A4(n23113), .ZN(
        n23100) );
  NAND4_X1 U24297 ( .A1(n23080), .A2(n23081), .A3(n23082), .A4(n23083), .ZN(
        n4968) );
  AOI221_X1 U24298 ( .B1(n24441), .B2(n24392), .C1(n24435), .C2(n19881), .A(
        n23096), .ZN(n23081) );
  AOI221_X1 U24299 ( .B1(n24417), .B2(n19487), .C1(n24410), .C2(OUT2[36]), .A(
        n23097), .ZN(n23080) );
  NOR4_X1 U24300 ( .A1(n23092), .A2(n23093), .A3(n23094), .A4(n23095), .ZN(
        n23082) );
  NAND4_X1 U24301 ( .A1(n23062), .A2(n23063), .A3(n23064), .A4(n23065), .ZN(
        n4969) );
  AOI221_X1 U24302 ( .B1(n24441), .B2(n24393), .C1(n24435), .C2(n19880), .A(
        n23078), .ZN(n23063) );
  AOI221_X1 U24303 ( .B1(n24417), .B2(n19486), .C1(n24410), .C2(OUT2[37]), .A(
        n23079), .ZN(n23062) );
  NOR4_X1 U24304 ( .A1(n23074), .A2(n23075), .A3(n23076), .A4(n23077), .ZN(
        n23064) );
  NAND4_X1 U24305 ( .A1(n23044), .A2(n23045), .A3(n23046), .A4(n23047), .ZN(
        n4970) );
  AOI221_X1 U24306 ( .B1(n24441), .B2(n24394), .C1(n24435), .C2(n19879), .A(
        n23060), .ZN(n23045) );
  AOI221_X1 U24307 ( .B1(n24417), .B2(n19485), .C1(n24410), .C2(OUT2[38]), .A(
        n23061), .ZN(n23044) );
  NOR4_X1 U24308 ( .A1(n23056), .A2(n23057), .A3(n23058), .A4(n23059), .ZN(
        n23046) );
  NAND4_X1 U24309 ( .A1(n23026), .A2(n23027), .A3(n23028), .A4(n23029), .ZN(
        n4971) );
  AOI221_X1 U24310 ( .B1(n24441), .B2(n24395), .C1(n24435), .C2(n19878), .A(
        n23042), .ZN(n23027) );
  AOI221_X1 U24311 ( .B1(n24417), .B2(n19484), .C1(n24410), .C2(OUT2[39]), .A(
        n23043), .ZN(n23026) );
  NOR4_X1 U24312 ( .A1(n23038), .A2(n23039), .A3(n23040), .A4(n23041), .ZN(
        n23028) );
  OAI22_X1 U24313 ( .A1(n24888), .A2(n25347), .B1(n24886), .B2(n20906), .ZN(
        n5316) );
  OAI22_X1 U24314 ( .A1(n24888), .A2(n25350), .B1(n24886), .B2(n20905), .ZN(
        n5317) );
  OAI22_X1 U24315 ( .A1(n24888), .A2(n25353), .B1(n24886), .B2(n20904), .ZN(
        n5318) );
  OAI22_X1 U24316 ( .A1(n24888), .A2(n25356), .B1(n24886), .B2(n20903), .ZN(
        n5319) );
  OAI22_X1 U24317 ( .A1(n24888), .A2(n25359), .B1(n24886), .B2(n20902), .ZN(
        n5320) );
  OAI22_X1 U24318 ( .A1(n24889), .A2(n25362), .B1(n24886), .B2(n20901), .ZN(
        n5321) );
  OAI22_X1 U24319 ( .A1(n24889), .A2(n25365), .B1(n24886), .B2(n20900), .ZN(
        n5322) );
  OAI22_X1 U24320 ( .A1(n24889), .A2(n25368), .B1(n24886), .B2(n20899), .ZN(
        n5323) );
  OAI22_X1 U24321 ( .A1(n24889), .A2(n25371), .B1(n24886), .B2(n20898), .ZN(
        n5324) );
  OAI22_X1 U24322 ( .A1(n24889), .A2(n25374), .B1(n24886), .B2(n20897), .ZN(
        n5325) );
  OAI22_X1 U24323 ( .A1(n24890), .A2(n25377), .B1(n24886), .B2(n20896), .ZN(
        n5326) );
  OAI22_X1 U24324 ( .A1(n24890), .A2(n25380), .B1(n24886), .B2(n20895), .ZN(
        n5327) );
  OAI22_X1 U24325 ( .A1(n24890), .A2(n25383), .B1(n24887), .B2(n20894), .ZN(
        n5328) );
  OAI22_X1 U24326 ( .A1(n24890), .A2(n25386), .B1(n24887), .B2(n20893), .ZN(
        n5329) );
  OAI22_X1 U24327 ( .A1(n24890), .A2(n25389), .B1(n24887), .B2(n20892), .ZN(
        n5330) );
  OAI22_X1 U24328 ( .A1(n24891), .A2(n25392), .B1(n24887), .B2(n20891), .ZN(
        n5331) );
  OAI22_X1 U24329 ( .A1(n24891), .A2(n25395), .B1(n24887), .B2(n20890), .ZN(
        n5332) );
  OAI22_X1 U24330 ( .A1(n24891), .A2(n25398), .B1(n24887), .B2(n20889), .ZN(
        n5333) );
  OAI22_X1 U24331 ( .A1(n24891), .A2(n25401), .B1(n24887), .B2(n20888), .ZN(
        n5334) );
  OAI22_X1 U24332 ( .A1(n24891), .A2(n25404), .B1(n24887), .B2(n20887), .ZN(
        n5335) );
  OAI22_X1 U24333 ( .A1(n24892), .A2(n25407), .B1(n24887), .B2(n20886), .ZN(
        n5336) );
  OAI22_X1 U24334 ( .A1(n24892), .A2(n25410), .B1(n24887), .B2(n20885), .ZN(
        n5337) );
  OAI22_X1 U24335 ( .A1(n24892), .A2(n25413), .B1(n24887), .B2(n20884), .ZN(
        n5338) );
  OAI22_X1 U24336 ( .A1(n24892), .A2(n25416), .B1(n24887), .B2(n20883), .ZN(
        n5339) );
  OAI22_X1 U24337 ( .A1(n24892), .A2(n25419), .B1(n24886), .B2(n20882), .ZN(
        n5340) );
  OAI22_X1 U24338 ( .A1(n24893), .A2(n25422), .B1(n24887), .B2(n20881), .ZN(
        n5341) );
  OAI22_X1 U24339 ( .A1(n24893), .A2(n25425), .B1(n24885), .B2(n20880), .ZN(
        n5342) );
  OAI22_X1 U24340 ( .A1(n24893), .A2(n25428), .B1(n24886), .B2(n20879), .ZN(
        n5343) );
  OAI22_X1 U24341 ( .A1(n24893), .A2(n25431), .B1(n24887), .B2(n20878), .ZN(
        n5344) );
  OAI22_X1 U24342 ( .A1(n24893), .A2(n25434), .B1(n24885), .B2(n20877), .ZN(
        n5345) );
  OAI22_X1 U24343 ( .A1(n24894), .A2(n25437), .B1(n24886), .B2(n20876), .ZN(
        n5346) );
  OAI22_X1 U24344 ( .A1(n24894), .A2(n25440), .B1(n24887), .B2(n20875), .ZN(
        n5347) );
  OAI22_X1 U24345 ( .A1(n24894), .A2(n25443), .B1(n24885), .B2(n20874), .ZN(
        n5348) );
  OAI22_X1 U24346 ( .A1(n24894), .A2(n25446), .B1(n24886), .B2(n20873), .ZN(
        n5349) );
  OAI22_X1 U24347 ( .A1(n24894), .A2(n25449), .B1(n24887), .B2(n20872), .ZN(
        n5350) );
  OAI22_X1 U24348 ( .A1(n24895), .A2(n25452), .B1(n24885), .B2(n20871), .ZN(
        n5351) );
  OAI22_X1 U24349 ( .A1(n24895), .A2(n25455), .B1(n21292), .B2(n20870), .ZN(
        n5352) );
  OAI22_X1 U24350 ( .A1(n24895), .A2(n25458), .B1(n24885), .B2(n20869), .ZN(
        n5353) );
  OAI22_X1 U24351 ( .A1(n24895), .A2(n25461), .B1(n21292), .B2(n20868), .ZN(
        n5354) );
  OAI22_X1 U24352 ( .A1(n24895), .A2(n25464), .B1(n24885), .B2(n20867), .ZN(
        n5355) );
  OAI22_X1 U24353 ( .A1(n24896), .A2(n25467), .B1(n21292), .B2(n20866), .ZN(
        n5356) );
  OAI22_X1 U24354 ( .A1(n24896), .A2(n25470), .B1(n24885), .B2(n20865), .ZN(
        n5357) );
  OAI22_X1 U24355 ( .A1(n24896), .A2(n25473), .B1(n24886), .B2(n20864), .ZN(
        n5358) );
  OAI22_X1 U24356 ( .A1(n24896), .A2(n25476), .B1(n24887), .B2(n20863), .ZN(
        n5359) );
  OAI22_X1 U24357 ( .A1(n24896), .A2(n25479), .B1(n24885), .B2(n20862), .ZN(
        n5360) );
  OAI22_X1 U24358 ( .A1(n24897), .A2(n25482), .B1(n24885), .B2(n20861), .ZN(
        n5361) );
  OAI22_X1 U24359 ( .A1(n24897), .A2(n25485), .B1(n24886), .B2(n20860), .ZN(
        n5362) );
  OAI22_X1 U24360 ( .A1(n24897), .A2(n25488), .B1(n24887), .B2(n20859), .ZN(
        n5363) );
  OAI22_X1 U24361 ( .A1(n24897), .A2(n25491), .B1(n24885), .B2(n20858), .ZN(
        n5364) );
  OAI22_X1 U24362 ( .A1(n24897), .A2(n25494), .B1(n24885), .B2(n20857), .ZN(
        n5365) );
  OAI22_X1 U24363 ( .A1(n24898), .A2(n25497), .B1(n21292), .B2(n20856), .ZN(
        n5366) );
  OAI22_X1 U24364 ( .A1(n24898), .A2(n25500), .B1(n24885), .B2(n20855), .ZN(
        n5367) );
  OAI22_X1 U24365 ( .A1(n24898), .A2(n25503), .B1(n21292), .B2(n20854), .ZN(
        n5368) );
  OAI22_X1 U24366 ( .A1(n24898), .A2(n25506), .B1(n24885), .B2(n20853), .ZN(
        n5369) );
  OAI22_X1 U24367 ( .A1(n24898), .A2(n25509), .B1(n21292), .B2(n20852), .ZN(
        n5370) );
  OAI22_X1 U24368 ( .A1(n24899), .A2(n25512), .B1(n24885), .B2(n20851), .ZN(
        n5371) );
  OAI22_X1 U24369 ( .A1(n24899), .A2(n25515), .B1(n21292), .B2(n20850), .ZN(
        n5372) );
  OAI22_X1 U24370 ( .A1(n24899), .A2(n25518), .B1(n24885), .B2(n20849), .ZN(
        n5373) );
  OAI22_X1 U24371 ( .A1(n24899), .A2(n25521), .B1(n21292), .B2(n20848), .ZN(
        n5374) );
  OAI22_X1 U24372 ( .A1(n24899), .A2(n25524), .B1(n24885), .B2(n20847), .ZN(
        n5375) );
  NOR3_X1 U24373 ( .A1(n19199), .A2(ADD_RD2[0]), .A3(n19200), .ZN(n23748) );
  NOR3_X1 U24374 ( .A1(n19199), .A2(ADD_RD2[3]), .A3(n19203), .ZN(n23745) );
  NOR3_X1 U24375 ( .A1(n19203), .A2(ADD_RD2[4]), .A3(n19200), .ZN(n23742) );
  NOR3_X1 U24376 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n19196), .ZN(n22553)
         );
  NOR2_X1 U24377 ( .A1(n19197), .A2(ADD_RD1[2]), .ZN(n22543) );
  NOR3_X1 U24378 ( .A1(n19196), .A2(ADD_RD1[4]), .A3(n19198), .ZN(n22554) );
  NOR3_X1 U24379 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(
        n22558) );
  NOR3_X1 U24380 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n19198), .ZN(n22557)
         );
  NOR3_X1 U24381 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n19199), .ZN(n23738)
         );
  NOR3_X1 U24382 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n19200), .ZN(n23741)
         );
  AND2_X1 U24383 ( .A1(ADD_RD1[2]), .A2(n19197), .ZN(n22538) );
  NOR2_X1 U24384 ( .A1(n24408), .A2(WR), .ZN(n23761) );
  NOR2_X1 U24385 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n23757) );
  NOR2_X1 U24386 ( .A1(n19201), .A2(ADD_RD2[1]), .ZN(n23759) );
  NOR2_X1 U24387 ( .A1(n19202), .A2(ADD_RD2[2]), .ZN(n23758) );
  AND2_X1 U24388 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n22540) );
  NAND2_X1 U24389 ( .A1(n24803), .A2(WR), .ZN(n21297) );
  INV_X1 U24390 ( .A(ADD_RD2[3]), .ZN(n19200) );
  INV_X1 U24391 ( .A(ADD_RD2[4]), .ZN(n19199) );
  NAND2_X1 U24392 ( .A1(RD2), .A2(ENABLE), .ZN(n22608) );
  AND2_X1 U24393 ( .A1(n23760), .A2(ADD_RD2[0]), .ZN(n23756) );
  AND3_X1 U24394 ( .A1(n19198), .A2(n19196), .A3(ADD_RD1[4]), .ZN(n22545) );
  AND3_X1 U24395 ( .A1(ADD_RD1[3]), .A2(n19198), .A3(ADD_RD1[4]), .ZN(n22537)
         );
  AND3_X1 U24396 ( .A1(ADD_RD1[0]), .A2(n19196), .A3(ADD_RD1[4]), .ZN(n22546)
         );
  AND3_X1 U24397 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(ADD_RD1[4]), .ZN(
        n22539) );
  INV_X1 U24398 ( .A(ADD_RD2[0]), .ZN(n19203) );
  NAND2_X1 U24399 ( .A1(DATAIN[0]), .A2(n25562), .ZN(n21252) );
  NAND2_X1 U24400 ( .A1(DATAIN[1]), .A2(n25562), .ZN(n21251) );
  NAND2_X1 U24401 ( .A1(DATAIN[2]), .A2(n25562), .ZN(n21250) );
  NAND2_X1 U24402 ( .A1(DATAIN[4]), .A2(n25562), .ZN(n21248) );
  NAND2_X1 U24403 ( .A1(DATAIN[3]), .A2(n25561), .ZN(n21249) );
  NAND2_X1 U24404 ( .A1(DATAIN[5]), .A2(n25561), .ZN(n21247) );
  NAND2_X1 U24405 ( .A1(DATAIN[6]), .A2(n25561), .ZN(n21246) );
  NAND2_X1 U24406 ( .A1(DATAIN[7]), .A2(n25561), .ZN(n21245) );
  NAND2_X1 U24407 ( .A1(DATAIN[8]), .A2(n25561), .ZN(n21244) );
  NAND2_X1 U24408 ( .A1(DATAIN[9]), .A2(n25561), .ZN(n21243) );
  NAND2_X1 U24409 ( .A1(DATAIN[10]), .A2(n25561), .ZN(n21242) );
  NAND2_X1 U24410 ( .A1(DATAIN[11]), .A2(n25561), .ZN(n21241) );
  NAND2_X1 U24411 ( .A1(DATAIN[12]), .A2(n25561), .ZN(n21240) );
  NAND2_X1 U24412 ( .A1(DATAIN[13]), .A2(n25561), .ZN(n21239) );
  NAND2_X1 U24413 ( .A1(DATAIN[14]), .A2(n25561), .ZN(n21238) );
  NAND2_X1 U24414 ( .A1(DATAIN[15]), .A2(n25560), .ZN(n21237) );
  NAND2_X1 U24415 ( .A1(DATAIN[16]), .A2(n25561), .ZN(n21236) );
  NAND2_X1 U24416 ( .A1(DATAIN[17]), .A2(n25560), .ZN(n21235) );
  NAND2_X1 U24417 ( .A1(DATAIN[18]), .A2(n25560), .ZN(n21234) );
  NAND2_X1 U24418 ( .A1(DATAIN[19]), .A2(n25560), .ZN(n21233) );
  NAND2_X1 U24419 ( .A1(DATAIN[20]), .A2(n25560), .ZN(n21232) );
  NAND2_X1 U24420 ( .A1(DATAIN[21]), .A2(n25560), .ZN(n21231) );
  NAND2_X1 U24421 ( .A1(DATAIN[22]), .A2(n25560), .ZN(n21230) );
  NAND2_X1 U24422 ( .A1(DATAIN[23]), .A2(n25559), .ZN(n21229) );
  NAND2_X1 U24423 ( .A1(DATAIN[24]), .A2(n25560), .ZN(n21228) );
  NAND2_X1 U24424 ( .A1(DATAIN[25]), .A2(n25560), .ZN(n21227) );
  NAND2_X1 U24425 ( .A1(DATAIN[26]), .A2(n25560), .ZN(n21226) );
  NAND2_X1 U24426 ( .A1(DATAIN[27]), .A2(n25560), .ZN(n21225) );
  NAND2_X1 U24427 ( .A1(DATAIN[28]), .A2(n25560), .ZN(n21224) );
  NAND2_X1 U24428 ( .A1(DATAIN[29]), .A2(n25559), .ZN(n21223) );
  NAND2_X1 U24429 ( .A1(DATAIN[30]), .A2(n25559), .ZN(n21222) );
  NAND2_X1 U24430 ( .A1(DATAIN[31]), .A2(n25559), .ZN(n21221) );
  NAND2_X1 U24431 ( .A1(DATAIN[32]), .A2(n25559), .ZN(n21220) );
  NAND2_X1 U24432 ( .A1(DATAIN[33]), .A2(n25559), .ZN(n21219) );
  NAND2_X1 U24433 ( .A1(DATAIN[34]), .A2(n25559), .ZN(n21218) );
  NAND2_X1 U24434 ( .A1(DATAIN[35]), .A2(n25559), .ZN(n21217) );
  NAND2_X1 U24435 ( .A1(DATAIN[36]), .A2(n25559), .ZN(n21216) );
  NAND2_X1 U24436 ( .A1(DATAIN[37]), .A2(n25559), .ZN(n21215) );
  NAND2_X1 U24437 ( .A1(DATAIN[38]), .A2(n25559), .ZN(n21214) );
  NAND2_X1 U24438 ( .A1(DATAIN[39]), .A2(n25559), .ZN(n21213) );
  NAND2_X1 U24439 ( .A1(DATAIN[40]), .A2(n25558), .ZN(n21212) );
  NAND2_X1 U24440 ( .A1(DATAIN[41]), .A2(n25558), .ZN(n21211) );
  NAND2_X1 U24441 ( .A1(DATAIN[42]), .A2(n25558), .ZN(n21210) );
  NAND2_X1 U24442 ( .A1(DATAIN[43]), .A2(n25558), .ZN(n21209) );
  NAND2_X1 U24443 ( .A1(DATAIN[44]), .A2(n25558), .ZN(n21208) );
  NAND2_X1 U24444 ( .A1(DATAIN[45]), .A2(n25558), .ZN(n21207) );
  NAND2_X1 U24445 ( .A1(DATAIN[46]), .A2(n25558), .ZN(n21206) );
  NAND2_X1 U24446 ( .A1(DATAIN[47]), .A2(n25558), .ZN(n21205) );
  NAND2_X1 U24447 ( .A1(DATAIN[48]), .A2(n25558), .ZN(n21204) );
  NAND2_X1 U24448 ( .A1(DATAIN[49]), .A2(n25558), .ZN(n21203) );
  NAND2_X1 U24449 ( .A1(DATAIN[50]), .A2(n25558), .ZN(n21202) );
  NAND2_X1 U24450 ( .A1(DATAIN[51]), .A2(n25558), .ZN(n21201) );
  NAND2_X1 U24451 ( .A1(DATAIN[52]), .A2(n25557), .ZN(n21200) );
  NAND2_X1 U24452 ( .A1(DATAIN[53]), .A2(n25557), .ZN(n21199) );
  NAND2_X1 U24453 ( .A1(DATAIN[54]), .A2(n25557), .ZN(n21198) );
  NAND2_X1 U24454 ( .A1(DATAIN[55]), .A2(n25557), .ZN(n21197) );
  NAND2_X1 U24455 ( .A1(DATAIN[56]), .A2(n25557), .ZN(n21196) );
  NAND2_X1 U24456 ( .A1(DATAIN[57]), .A2(n25557), .ZN(n21195) );
  NAND2_X1 U24457 ( .A1(DATAIN[58]), .A2(n25557), .ZN(n21194) );
  NAND2_X1 U24458 ( .A1(DATAIN[59]), .A2(n25557), .ZN(n21193) );
  NAND2_X1 U24459 ( .A1(DATAIN[60]), .A2(n25557), .ZN(n21192) );
  NAND2_X1 U24460 ( .A1(DATAIN[61]), .A2(n25557), .ZN(n21191) );
  NAND2_X1 U24461 ( .A1(DATAIN[62]), .A2(n25557), .ZN(n21190) );
  NAND2_X1 U24462 ( .A1(DATAIN[63]), .A2(n25557), .ZN(n21188) );
  AND2_X1 U24463 ( .A1(RD1), .A2(ENABLE), .ZN(n21298) );
  INV_X1 U24464 ( .A(ADD_RD1[0]), .ZN(n19198) );
  INV_X1 U24465 ( .A(ADD_RD1[3]), .ZN(n19196) );
  AND2_X1 U24466 ( .A1(WR), .A2(ENABLE), .ZN(n21269) );
  INV_X1 U24467 ( .A(ADD_WR[2]), .ZN(n19193) );
  INV_X1 U24468 ( .A(ADD_WR[0]), .ZN(n19195) );
  INV_X1 U24469 ( .A(ADD_WR[1]), .ZN(n19194) );
  INV_X1 U24470 ( .A(ADD_RD2[2]), .ZN(n19201) );
  INV_X1 U24471 ( .A(DATAIN[40]), .ZN(n19227) );
  INV_X1 U24472 ( .A(DATAIN[41]), .ZN(n19226) );
  INV_X1 U24473 ( .A(DATAIN[42]), .ZN(n19225) );
  INV_X1 U24474 ( .A(DATAIN[43]), .ZN(n19224) );
  INV_X1 U24475 ( .A(DATAIN[44]), .ZN(n19223) );
  INV_X1 U24476 ( .A(DATAIN[45]), .ZN(n19222) );
  INV_X1 U24477 ( .A(DATAIN[46]), .ZN(n19221) );
  INV_X1 U24478 ( .A(DATAIN[47]), .ZN(n19220) );
  INV_X1 U24479 ( .A(DATAIN[48]), .ZN(n19219) );
  INV_X1 U24480 ( .A(DATAIN[49]), .ZN(n19218) );
  INV_X1 U24481 ( .A(DATAIN[50]), .ZN(n19217) );
  INV_X1 U24482 ( .A(DATAIN[51]), .ZN(n19216) );
  INV_X1 U24483 ( .A(DATAIN[52]), .ZN(n19215) );
  INV_X1 U24484 ( .A(DATAIN[53]), .ZN(n19214) );
  INV_X1 U24485 ( .A(DATAIN[54]), .ZN(n19213) );
  INV_X1 U24486 ( .A(DATAIN[55]), .ZN(n19212) );
  INV_X1 U24487 ( .A(DATAIN[56]), .ZN(n19211) );
  INV_X1 U24488 ( .A(DATAIN[57]), .ZN(n19210) );
  INV_X1 U24489 ( .A(DATAIN[58]), .ZN(n19209) );
  INV_X1 U24490 ( .A(DATAIN[59]), .ZN(n19208) );
  INV_X1 U24491 ( .A(DATAIN[60]), .ZN(n19207) );
  INV_X1 U24492 ( .A(DATAIN[61]), .ZN(n19206) );
  INV_X1 U24493 ( .A(DATAIN[62]), .ZN(n19205) );
  INV_X1 U24494 ( .A(DATAIN[63]), .ZN(n19204) );
  INV_X1 U24495 ( .A(DATAIN[0]), .ZN(n19267) );
  INV_X1 U24496 ( .A(DATAIN[1]), .ZN(n19266) );
  INV_X1 U24497 ( .A(DATAIN[2]), .ZN(n19265) );
  INV_X1 U24498 ( .A(DATAIN[3]), .ZN(n19264) );
  INV_X1 U24499 ( .A(DATAIN[4]), .ZN(n19263) );
  INV_X1 U24500 ( .A(DATAIN[5]), .ZN(n19262) );
  INV_X1 U24501 ( .A(DATAIN[6]), .ZN(n19261) );
  INV_X1 U24502 ( .A(DATAIN[7]), .ZN(n19260) );
  INV_X1 U24503 ( .A(DATAIN[8]), .ZN(n19259) );
  INV_X1 U24504 ( .A(DATAIN[9]), .ZN(n19258) );
  INV_X1 U24505 ( .A(DATAIN[10]), .ZN(n19257) );
  INV_X1 U24506 ( .A(DATAIN[11]), .ZN(n19256) );
  INV_X1 U24507 ( .A(DATAIN[12]), .ZN(n19255) );
  INV_X1 U24508 ( .A(DATAIN[13]), .ZN(n19254) );
  INV_X1 U24509 ( .A(DATAIN[14]), .ZN(n19253) );
  INV_X1 U24510 ( .A(DATAIN[15]), .ZN(n19252) );
  INV_X1 U24511 ( .A(DATAIN[16]), .ZN(n19251) );
  INV_X1 U24512 ( .A(DATAIN[17]), .ZN(n19250) );
  INV_X1 U24513 ( .A(DATAIN[18]), .ZN(n19249) );
  INV_X1 U24514 ( .A(DATAIN[19]), .ZN(n19248) );
  INV_X1 U24515 ( .A(DATAIN[20]), .ZN(n19247) );
  INV_X1 U24516 ( .A(DATAIN[21]), .ZN(n19246) );
  INV_X1 U24517 ( .A(DATAIN[22]), .ZN(n19245) );
  INV_X1 U24518 ( .A(DATAIN[23]), .ZN(n19244) );
  INV_X1 U24519 ( .A(DATAIN[24]), .ZN(n19243) );
  INV_X1 U24520 ( .A(DATAIN[25]), .ZN(n19242) );
  INV_X1 U24521 ( .A(DATAIN[26]), .ZN(n19241) );
  INV_X1 U24522 ( .A(DATAIN[27]), .ZN(n19240) );
  INV_X1 U24523 ( .A(DATAIN[28]), .ZN(n19239) );
  INV_X1 U24524 ( .A(DATAIN[29]), .ZN(n19238) );
  INV_X1 U24525 ( .A(DATAIN[30]), .ZN(n19237) );
  INV_X1 U24526 ( .A(DATAIN[31]), .ZN(n19236) );
  INV_X1 U24527 ( .A(DATAIN[32]), .ZN(n19235) );
  INV_X1 U24528 ( .A(DATAIN[33]), .ZN(n19234) );
  INV_X1 U24529 ( .A(DATAIN[34]), .ZN(n19233) );
  INV_X1 U24530 ( .A(DATAIN[35]), .ZN(n19232) );
  INV_X1 U24531 ( .A(DATAIN[36]), .ZN(n19231) );
  INV_X1 U24532 ( .A(DATAIN[37]), .ZN(n19230) );
  INV_X1 U24533 ( .A(DATAIN[38]), .ZN(n19229) );
  INV_X1 U24534 ( .A(DATAIN[39]), .ZN(n19228) );
  INV_X1 U24535 ( .A(ADD_RD2[1]), .ZN(n19202) );
  INV_X1 U24536 ( .A(ADD_RD1[1]), .ZN(n19197) );
  INV_X1 U24537 ( .A(WR), .ZN(n19190) );
  INV_X1 U24538 ( .A(ADD_WR[4]), .ZN(n19191) );
  INV_X1 U24539 ( .A(ADD_WR[3]), .ZN(n19192) );
  INV_X1 U24540 ( .A(RESET), .ZN(n19189) );
  CLKBUF_X1 U24541 ( .A(n22611), .Z(n24401) );
  CLKBUF_X1 U24542 ( .A(n22610), .Z(n24407) );
  CLKBUF_X1 U24543 ( .A(n22608), .Z(n24413) );
  CLKBUF_X1 U24544 ( .A(n22607), .Z(n24419) );
  CLKBUF_X1 U24545 ( .A(n22606), .Z(n24425) );
  CLKBUF_X1 U24546 ( .A(n22605), .Z(n24431) );
  CLKBUF_X1 U24547 ( .A(n22603), .Z(n24437) );
  CLKBUF_X1 U24548 ( .A(n22602), .Z(n24443) );
  CLKBUF_X1 U24549 ( .A(n22601), .Z(n24449) );
  CLKBUF_X1 U24550 ( .A(n22600), .Z(n24455) );
  CLKBUF_X1 U24551 ( .A(n22599), .Z(n24461) );
  CLKBUF_X1 U24552 ( .A(n22598), .Z(n24467) );
  CLKBUF_X1 U24553 ( .A(n22597), .Z(n24473) );
  CLKBUF_X1 U24554 ( .A(n22596), .Z(n24479) );
  CLKBUF_X1 U24555 ( .A(n22595), .Z(n24485) );
  CLKBUF_X1 U24556 ( .A(n22594), .Z(n24491) );
  CLKBUF_X1 U24557 ( .A(n22593), .Z(n24497) );
  CLKBUF_X1 U24558 ( .A(n22588), .Z(n24503) );
  CLKBUF_X1 U24559 ( .A(n22587), .Z(n24509) );
  CLKBUF_X1 U24560 ( .A(n22586), .Z(n24515) );
  CLKBUF_X1 U24561 ( .A(n22584), .Z(n24521) );
  CLKBUF_X1 U24562 ( .A(n22583), .Z(n24527) );
  CLKBUF_X1 U24563 ( .A(n22582), .Z(n24533) );
  CLKBUF_X1 U24564 ( .A(n22581), .Z(n24539) );
  CLKBUF_X1 U24565 ( .A(n22579), .Z(n24545) );
  CLKBUF_X1 U24566 ( .A(n22578), .Z(n24551) );
  CLKBUF_X1 U24567 ( .A(n22577), .Z(n24557) );
  CLKBUF_X1 U24568 ( .A(n22576), .Z(n24563) );
  CLKBUF_X1 U24569 ( .A(n22574), .Z(n24569) );
  CLKBUF_X1 U24570 ( .A(n22573), .Z(n24575) );
  CLKBUF_X1 U24571 ( .A(n22572), .Z(n24581) );
  CLKBUF_X1 U24572 ( .A(n22571), .Z(n24587) );
  CLKBUF_X1 U24573 ( .A(n22569), .Z(n24593) );
  CLKBUF_X1 U24574 ( .A(n22568), .Z(n24599) );
  CLKBUF_X1 U24575 ( .A(n21350), .Z(n24605) );
  CLKBUF_X1 U24576 ( .A(n21349), .Z(n24611) );
  CLKBUF_X1 U24577 ( .A(n21347), .Z(n24617) );
  CLKBUF_X1 U24578 ( .A(n21346), .Z(n24623) );
  CLKBUF_X1 U24579 ( .A(n21345), .Z(n24629) );
  CLKBUF_X1 U24580 ( .A(n21344), .Z(n24635) );
  CLKBUF_X1 U24581 ( .A(n21342), .Z(n24641) );
  CLKBUF_X1 U24582 ( .A(n21341), .Z(n24647) );
  CLKBUF_X1 U24583 ( .A(n21340), .Z(n24653) );
  CLKBUF_X1 U24584 ( .A(n21339), .Z(n24659) );
  CLKBUF_X1 U24585 ( .A(n21337), .Z(n24665) );
  CLKBUF_X1 U24586 ( .A(n21336), .Z(n24671) );
  CLKBUF_X1 U24587 ( .A(n21335), .Z(n24677) );
  CLKBUF_X1 U24588 ( .A(n21334), .Z(n24683) );
  CLKBUF_X1 U24589 ( .A(n21332), .Z(n24689) );
  CLKBUF_X1 U24590 ( .A(n21331), .Z(n24695) );
  CLKBUF_X1 U24591 ( .A(n21326), .Z(n24701) );
  CLKBUF_X1 U24592 ( .A(n21325), .Z(n24707) );
  CLKBUF_X1 U24593 ( .A(n21323), .Z(n24713) );
  CLKBUF_X1 U24594 ( .A(n21322), .Z(n24719) );
  CLKBUF_X1 U24595 ( .A(n21321), .Z(n24725) );
  CLKBUF_X1 U24596 ( .A(n21320), .Z(n24731) );
  CLKBUF_X1 U24597 ( .A(n21318), .Z(n24737) );
  CLKBUF_X1 U24598 ( .A(n21317), .Z(n24743) );
  CLKBUF_X1 U24599 ( .A(n21316), .Z(n24749) );
  CLKBUF_X1 U24600 ( .A(n21315), .Z(n24755) );
  CLKBUF_X1 U24601 ( .A(n21313), .Z(n24761) );
  CLKBUF_X1 U24602 ( .A(n21312), .Z(n24767) );
  CLKBUF_X1 U24603 ( .A(n21311), .Z(n24773) );
  CLKBUF_X1 U24604 ( .A(n21310), .Z(n24779) );
  CLKBUF_X1 U24605 ( .A(n21308), .Z(n24785) );
  CLKBUF_X1 U24606 ( .A(n21307), .Z(n24791) );
  CLKBUF_X1 U24607 ( .A(n21302), .Z(n24797) );
  CLKBUF_X1 U24608 ( .A(n21298), .Z(n24803) );
  CLKBUF_X1 U24609 ( .A(n21297), .Z(n24809) );
  CLKBUF_X1 U24610 ( .A(n19189), .Z(n25554) );
  CLKBUF_X1 U24611 ( .A(n19189), .Z(n25555) );
  CLKBUF_X1 U24612 ( .A(n19189), .Z(n25556) );
endmodule

