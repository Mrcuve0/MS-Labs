package constants is
  
  constant radixN : integer := 4;     -- Radix of the adder
  constant numBit : integer := 32;    -- Number of bits of the adder

end package constants;
