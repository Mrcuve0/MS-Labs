
package constants is

  constant numBitData : integer := 64;
  constant numRegs    : integer := 32;

end package constants;
