

    module controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 ( 
        A, INC_DEC, SUM );
  input [31:0] A;
  output [31:0] SUM;
  input INC_DEC;
  wire   n7, n8, n9;
  wire   [31:0] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(INC_DEC), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(INC_DEC), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(INC_DEC), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(n8), .CI(carry[28]), .CO(carry[29]), .S(SUM[28])
         );
  FA_X1 U1_27 ( .A(A[27]), .B(INC_DEC), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(n8), .CI(carry[26]), .CO(carry[27]), .S(SUM[26])
         );
  FA_X1 U1_25 ( .A(A[25]), .B(INC_DEC), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(n8), .CI(carry[24]), .CO(carry[25]), .S(SUM[24])
         );
  FA_X1 U1_23 ( .A(A[23]), .B(INC_DEC), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(INC_DEC), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(INC_DEC), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(n8), .CI(carry[20]), .CO(carry[21]), .S(SUM[20])
         );
  FA_X1 U1_19 ( .A(A[19]), .B(n8), .CI(carry[19]), .CO(carry[20]), .S(SUM[19])
         );
  FA_X1 U1_18 ( .A(A[18]), .B(n8), .CI(carry[18]), .CO(carry[19]), .S(SUM[18])
         );
  FA_X1 U1_17 ( .A(A[17]), .B(n8), .CI(carry[17]), .CO(carry[18]), .S(SUM[17])
         );
  FA_X1 U1_16 ( .A(A[16]), .B(n8), .CI(carry[16]), .CO(carry[17]), .S(SUM[16])
         );
  FA_X1 U1_15 ( .A(A[15]), .B(n8), .CI(carry[15]), .CO(carry[16]), .S(SUM[15])
         );
  FA_X1 U1_14 ( .A(A[14]), .B(n8), .CI(carry[14]), .CO(carry[15]), .S(SUM[14])
         );
  FA_X1 U1_13 ( .A(A[13]), .B(n8), .CI(carry[13]), .CO(carry[14]), .S(SUM[13])
         );
  FA_X1 U1_12 ( .A(A[12]), .B(n8), .CI(carry[12]), .CO(carry[13]), .S(SUM[12])
         );
  FA_X1 U1_11 ( .A(A[11]), .B(n7), .CI(carry[11]), .CO(carry[12]), .S(SUM[11])
         );
  FA_X1 U1_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(SUM[10])
         );
  FA_X1 U1_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  FA_X1 U1_8 ( .A(A[8]), .B(n7), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(n7), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(n7), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(n7), .CI(n9), .CO(carry[1]) );
  INV_X1 U1 ( .A(n9), .ZN(n7) );
  INV_X1 U2 ( .A(n9), .ZN(n8) );
  INV_X1 U3 ( .A(INC_DEC), .ZN(n9) );
  INV_X1 U4 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 ( clk, 
        reset, enable, cwpOut, swpOut, call, ret, fill, spill, MMUStrobe, 
        dataACK );
  output [3:0] cwpOut;
  output [3:0] swpOut;
  input clk, reset, enable, call, ret, MMUStrobe;
  output fill, spill, dataACK;
  wire   \need_to_fill[0] , \need_to_spill[0] , N436, N437, N438, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, n65, n66, n73, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n4, n6, n8, n9, n192, n205, n214, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n67, n68, n69, n70, n71, n72, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n219, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271;
  wire   [2:0] nextState;
  wire   [3:0] cansaveNext;
  wire   [3:0] canrestoreNext;
  wire   [31:0] actual_round;

  DLH_X1 \cansaveNext_reg[2]  ( .G(N442), .D(N445), .Q(cansaveNext[2]) );
  DLH_X1 \cansaveNext_reg[3]  ( .G(N442), .D(N446), .Q(cansaveNext[3]) );
  DFF_X1 \cansave_reg[3]  ( .D(n227), .CK(clk), .Q(n8), .QN(n244) );
  DLH_X1 \nextState_reg[1]  ( .G(N447), .D(N449), .Q(nextState[1]) );
  DLH_X1 \nextState_reg[0]  ( .G(N447), .D(N448), .Q(nextState[0]) );
  DLH_X1 \nextState_reg[2]  ( .G(N447), .D(N450), .Q(nextState[2]) );
  DLH_X1 \swp_reg[0]  ( .G(N460), .D(N461), .Q(swpOut[0]) );
  DLH_X1 \swp_reg[1]  ( .G(N460), .D(N462), .Q(swpOut[1]) );
  DLH_X1 \actual_round_reg[31]  ( .G(n233), .D(N497), .Q(actual_round[31]) );
  DLH_X1 \actual_round_reg[0]  ( .G(n234), .D(N466), .Q(actual_round[0]) );
  DLH_X1 \actual_round_reg[1]  ( .G(n233), .D(N467), .Q(actual_round[1]) );
  DLH_X1 \actual_round_reg[2]  ( .G(n233), .D(N468), .Q(actual_round[2]) );
  DLH_X1 \actual_round_reg[3]  ( .G(n233), .D(N469), .Q(actual_round[3]) );
  DLH_X1 \actual_round_reg[4]  ( .G(n233), .D(N470), .Q(actual_round[4]) );
  DLH_X1 \actual_round_reg[5]  ( .G(n233), .D(N471), .Q(actual_round[5]) );
  DLH_X1 \actual_round_reg[6]  ( .G(n233), .D(N472), .Q(actual_round[6]) );
  DLH_X1 \actual_round_reg[7]  ( .G(n233), .D(N473), .Q(actual_round[7]) );
  DLH_X1 \actual_round_reg[8]  ( .G(n233), .D(N474), .Q(actual_round[8]) );
  DLH_X1 \actual_round_reg[9]  ( .G(n233), .D(N475), .Q(actual_round[9]) );
  DLH_X1 \actual_round_reg[10]  ( .G(n233), .D(N476), .Q(actual_round[10]) );
  DLH_X1 \actual_round_reg[11]  ( .G(n232), .D(N477), .Q(actual_round[11]) );
  DLH_X1 \actual_round_reg[12]  ( .G(n232), .D(N478), .Q(actual_round[12]) );
  DLH_X1 \actual_round_reg[13]  ( .G(n232), .D(N479), .Q(actual_round[13]) );
  DLH_X1 \actual_round_reg[14]  ( .G(n232), .D(N480), .Q(actual_round[14]) );
  DLH_X1 \actual_round_reg[15]  ( .G(n232), .D(N481), .Q(actual_round[15]) );
  DLH_X1 \actual_round_reg[16]  ( .G(n232), .D(N482), .Q(actual_round[16]) );
  DLH_X1 \actual_round_reg[17]  ( .G(n232), .D(N483), .Q(actual_round[17]) );
  DLH_X1 \actual_round_reg[18]  ( .G(n232), .D(N484), .Q(actual_round[18]) );
  DLH_X1 \actual_round_reg[19]  ( .G(n232), .D(N485), .Q(actual_round[19]) );
  DLH_X1 \actual_round_reg[20]  ( .G(n232), .D(N486), .Q(actual_round[20]) );
  DLH_X1 \actual_round_reg[21]  ( .G(n232), .D(N487), .Q(actual_round[21]) );
  DLH_X1 \actual_round_reg[22]  ( .G(n234), .D(N488), .Q(actual_round[22]) );
  DLH_X1 \actual_round_reg[23]  ( .G(n234), .D(N489), .Q(actual_round[23]) );
  DLH_X1 \actual_round_reg[24]  ( .G(n234), .D(N490), .Q(actual_round[24]) );
  DLH_X1 \actual_round_reg[25]  ( .G(n234), .D(N491), .Q(actual_round[25]) );
  DLH_X1 \actual_round_reg[26]  ( .G(n234), .D(N492), .Q(actual_round[26]) );
  DLH_X1 \actual_round_reg[27]  ( .G(n234), .D(N493), .Q(actual_round[27]) );
  DLH_X1 \actual_round_reg[28]  ( .G(n234), .D(N494), .Q(actual_round[28]) );
  DLH_X1 \actual_round_reg[29]  ( .G(n234), .D(N495), .Q(actual_round[29]) );
  DLH_X1 \actual_round_reg[30]  ( .G(n234), .D(N496), .Q(actual_round[30]) );
  DLH_X1 \swp_reg[2]  ( .G(N460), .D(N463), .Q(swpOut[2]) );
  DLH_X1 \swp_reg[3]  ( .G(N460), .D(N464), .Q(swpOut[3]) );
  DLH_X1 \need_to_spill_reg[0]  ( .G(N438), .D(n157), .Q(\need_to_spill[0] )
         );
  DLH_X1 \canrestoreNext_reg[0]  ( .G(N442), .D(N451), .Q(canrestoreNext[0])
         );
  DFF_X1 \canrestore_reg[0]  ( .D(n223), .CK(clk), .Q(n9), .QN(n259) );
  DLH_X1 \canrestoreNext_reg[2]  ( .G(N442), .D(N453), .Q(canrestoreNext[2])
         );
  DLH_X1 \canrestoreNext_reg[3]  ( .G(N442), .D(N454), .Q(canrestoreNext[3])
         );
  DFF_X1 \canrestore_reg[3]  ( .D(n220), .CK(clk), .Q(n6), .QN(n260) );
  DLH_X1 \need_to_fill_reg[0]  ( .G(N436), .D(N437), .Q(\need_to_fill[0] ) );
  DLH_X1 \canrestoreNext_reg[1]  ( .G(N442), .D(N452), .Q(canrestoreNext[1])
         );
  DLH_X1 spill_reg ( .G(N440), .D(n158), .Q(spill) );
  DLH_X1 fill_reg ( .G(N440), .D(n159), .Q(fill) );
  DLH_X1 dataACK_reg ( .G(N440), .D(N441), .Q(dataACK) );
  DLH_X1 \cwp_reg[3]  ( .G(N455), .D(N459), .Q(cwpOut[3]) );
  DLH_X1 \cwp_reg[0]  ( .G(N455), .D(N456), .Q(cwpOut[0]) );
  DLH_X1 \cwp_reg[1]  ( .G(N455), .D(N457), .Q(cwpOut[1]) );
  DLH_X1 \cansaveNext_reg[1]  ( .G(N442), .D(N444), .Q(cansaveNext[1]) );
  DLH_X1 \cansaveNext_reg[0]  ( .G(N442), .D(N443), .Q(cansaveNext[0]) );
  DLH_X1 \cwp_reg[2]  ( .G(N455), .D(N458), .Q(cwpOut[2]) );
  DFF_X1 \cansave_reg[1]  ( .D(n229), .CK(clk), .Q(n156), .QN(n264) );
  XOR2_X1 U183 ( .A(n88), .B(n89), .Z(n85) );
  XOR2_X1 U184 ( .A(n119), .B(n120), .Z(n118) );
  XOR2_X1 U185 ( .A(n124), .B(n125), .Z(n75) );
  XOR2_X1 U186 ( .A(n127), .B(n134), .Z(n76) );
  XOR2_X1 U187 ( .A(n140), .B(n137), .Z(n77) );
  NAND3_X1 U188 ( .A1(n142), .A2(n253), .A3(n145), .ZN(n79) );
  NAND3_X1 U189 ( .A1(n245), .A2(n111), .A3(n109), .ZN(N442) );
  NAND3_X1 U190 ( .A1(n150), .A2(n107), .A3(call), .ZN(n145) );
  NAND3_X1 U191 ( .A1(n151), .A2(n248), .A3(n152), .ZN(n89) );
  NAND3_X1 U192 ( .A1(n110), .A2(ret), .A3(n100), .ZN(n152) );
  NAND3_X1 U193 ( .A1(n249), .A2(n245), .A3(n74), .ZN(N440) );
  NAND3_X1 U194 ( .A1(n133), .A2(n244), .A3(n192), .ZN(n107) );
  controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 r243 ( 
        .A(actual_round), .INC_DEC(n231), .SUM({N497, N496, N495, N494, N493, 
        N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, 
        N468, N467, N466}) );
  DFF_X1 \canrestore_reg[1]  ( .D(n222), .CK(clk), .QN(n214) );
  DFF_X1 \currentState_reg[1]  ( .D(n225), .CK(clk), .Q(n265), .QN(n65) );
  DFF_X1 \canrestore_reg[2]  ( .D(n221), .CK(clk), .Q(n262), .QN(n4) );
  DFF_X1 \cansave_reg[2]  ( .D(n228), .CK(clk), .QN(n192) );
  DFF_X1 \currentState_reg[2]  ( .D(n224), .CK(clk), .Q(n251), .QN(n205) );
  DFF_X1 \cansave_reg[0]  ( .D(n230), .CK(clk), .Q(n263), .QN(n73) );
  DFF_X1 \currentState_reg[0]  ( .D(n226), .CK(clk), .Q(n261), .QN(n66) );
  NOR3_X1 U3 ( .A1(n205), .A2(n66), .A3(n265), .ZN(n159) );
  NOR3_X1 U4 ( .A1(n261), .A2(n205), .A3(n265), .ZN(n158) );
  INV_X1 U5 ( .A(n130), .ZN(n248) );
  INV_X1 U6 ( .A(n103), .ZN(n249) );
  NAND2_X1 U7 ( .A1(n99), .A2(n248), .ZN(n83) );
  XNOR2_X1 U8 ( .A(n238), .B(n91), .ZN(n94) );
  AND2_X1 U9 ( .A1(n72), .A2(n99), .ZN(n74) );
  INV_X1 U10 ( .A(n122), .ZN(n243) );
  AND2_X1 U11 ( .A1(n99), .A2(n247), .ZN(n117) );
  NOR2_X1 U12 ( .A1(n258), .A2(n250), .ZN(N437) );
  INV_X1 U13 ( .A(n136), .ZN(n240) );
  BUF_X1 U14 ( .A(N465), .Z(n232) );
  BUF_X1 U15 ( .A(N465), .Z(n233) );
  BUF_X1 U16 ( .A(N465), .Z(n234) );
  NAND2_X1 U17 ( .A1(n253), .A2(n245), .ZN(N460) );
  INV_X1 U18 ( .A(n95), .ZN(n247) );
  NOR2_X1 U19 ( .A1(n74), .A2(n76), .ZN(N458) );
  NOR2_X1 U20 ( .A1(n74), .A2(n77), .ZN(N457) );
  INV_X1 U21 ( .A(N441), .ZN(n253) );
  OR2_X1 U22 ( .A1(n235), .A2(n127), .ZN(n126) );
  NOR3_X1 U23 ( .A1(n261), .A2(n251), .A3(n265), .ZN(n103) );
  XNOR2_X1 U24 ( .A(n240), .B(n128), .ZN(n134) );
  XNOR2_X1 U25 ( .A(n78), .B(n136), .ZN(n140) );
  AOI21_X1 U26 ( .B1(n258), .B2(n146), .A(n249), .ZN(n95) );
  OAI21_X1 U27 ( .B1(n252), .B2(n271), .A(n142), .ZN(n136) );
  AOI21_X1 U28 ( .B1(n96), .B2(n89), .A(n87), .ZN(n91) );
  NOR3_X1 U29 ( .A1(n249), .A2(n148), .A3(n269), .ZN(n130) );
  INV_X1 U30 ( .A(n50), .ZN(n266) );
  INV_X1 U31 ( .A(n80), .ZN(n245) );
  NAND2_X1 U32 ( .A1(n267), .A2(n50), .ZN(n43) );
  AOI22_X1 U33 ( .A1(n136), .A2(n137), .B1(n78), .B2(n138), .ZN(n127) );
  OR2_X1 U34 ( .A1(n137), .A2(n136), .ZN(n138) );
  NOR2_X1 U35 ( .A1(n110), .A2(n150), .ZN(n99) );
  NOR2_X1 U36 ( .A1(n246), .A2(n107), .ZN(n157) );
  OAI221_X1 U37 ( .B1(n248), .B2(n78), .C1(n117), .C2(n263), .A(n245), .ZN(
        N443) );
  NOR2_X1 U38 ( .A1(n159), .A2(n158), .ZN(n72) );
  NAND2_X1 U39 ( .A1(n111), .A2(n145), .ZN(n122) );
  INV_X1 U40 ( .A(n159), .ZN(n252) );
  AOI21_X1 U41 ( .B1(n219), .B2(n57), .A(n271), .ZN(N465) );
  NAND2_X1 U42 ( .A1(n158), .A2(n255), .ZN(n57) );
  INV_X1 U43 ( .A(n89), .ZN(n238) );
  INV_X1 U44 ( .A(n110), .ZN(n250) );
  OAI22_X1 U45 ( .A1(n238), .A2(n256), .B1(n97), .B2(n98), .ZN(N452) );
  INV_X1 U46 ( .A(n98), .ZN(n256) );
  NAND2_X1 U47 ( .A1(n257), .A2(n96), .ZN(n98) );
  AOI21_X1 U48 ( .B1(n238), .B2(n83), .A(n95), .ZN(n97) );
  XNOR2_X1 U49 ( .A(N467), .B(n67), .ZN(n64) );
  NOR2_X1 U50 ( .A1(n271), .A2(n72), .ZN(N441) );
  INV_X1 U51 ( .A(n158), .ZN(n254) );
  NAND2_X1 U52 ( .A1(n43), .A2(n50), .ZN(n44) );
  NAND2_X1 U53 ( .A1(n231), .A2(n68), .ZN(n60) );
  INV_X1 U54 ( .A(n148), .ZN(n258) );
  INV_X1 U55 ( .A(n150), .ZN(n246) );
  OAI211_X1 U56 ( .C1(n250), .C2(n149), .A(n249), .B(n155), .ZN(N436) );
  NOR2_X1 U57 ( .A1(N437), .A2(n159), .ZN(n155) );
  OAI211_X1 U58 ( .C1(n231), .C2(n68), .A(n60), .B(n245), .ZN(N463) );
  OAI211_X1 U59 ( .C1(n246), .C2(n268), .A(n249), .B(n154), .ZN(N438) );
  NOR2_X1 U60 ( .A1(n157), .A2(n158), .ZN(n154) );
  INV_X1 U61 ( .A(n63), .ZN(n255) );
  INV_X1 U62 ( .A(n87), .ZN(n257) );
  OAI21_X1 U63 ( .B1(n108), .B2(n268), .A(n109), .ZN(N449) );
  AOI21_X1 U64 ( .B1(n100), .B2(n110), .A(n241), .ZN(n108) );
  INV_X1 U65 ( .A(n111), .ZN(n241) );
  NOR2_X1 U66 ( .A1(n74), .A2(n78), .ZN(N456) );
  OR3_X1 U67 ( .A1(n250), .A2(n148), .A3(n149), .ZN(n142) );
  NOR2_X1 U68 ( .A1(n74), .A2(n75), .ZN(N459) );
  INV_X1 U69 ( .A(n85), .ZN(n236) );
  INV_X1 U70 ( .A(n146), .ZN(n269) );
  AND2_X1 U71 ( .A1(n238), .A2(n145), .ZN(n109) );
  OR2_X1 U72 ( .A1(n79), .A2(n80), .ZN(N455) );
  INV_X1 U73 ( .A(n128), .ZN(n235) );
  OAI211_X1 U74 ( .C1(n73), .C2(n43), .A(n44), .B(n45), .ZN(n230) );
  NAND2_X1 U75 ( .A1(cansaveNext[0]), .A2(n43), .ZN(n45) );
  OAI211_X1 U76 ( .C1(n66), .C2(n43), .A(n44), .B(n49), .ZN(n226) );
  NAND2_X1 U77 ( .A1(nextState[0]), .A2(n43), .ZN(n49) );
  OAI211_X1 U78 ( .C1(n43), .C2(n264), .A(n44), .B(n46), .ZN(n229) );
  NAND2_X1 U79 ( .A1(cansaveNext[1]), .A2(n43), .ZN(n46) );
  OAI21_X1 U80 ( .B1(n205), .B2(n43), .A(n52), .ZN(n224) );
  NAND2_X1 U81 ( .A1(nextState[2]), .A2(n266), .ZN(n52) );
  OAI21_X1 U82 ( .B1(n43), .B2(n260), .A(n56), .ZN(n220) );
  NAND2_X1 U83 ( .A1(canrestoreNext[3]), .A2(n266), .ZN(n56) );
  OAI21_X1 U84 ( .B1(n43), .B2(n259), .A(n53), .ZN(n223) );
  NAND2_X1 U85 ( .A1(canrestoreNext[0]), .A2(n266), .ZN(n53) );
  OAI21_X1 U86 ( .B1(n43), .B2(n244), .A(n48), .ZN(n227) );
  NAND2_X1 U87 ( .A1(cansaveNext[3]), .A2(n266), .ZN(n48) );
  OAI21_X1 U88 ( .B1(n4), .B2(n43), .A(n55), .ZN(n221) );
  NAND2_X1 U89 ( .A1(canrestoreNext[2]), .A2(n266), .ZN(n55) );
  OAI21_X1 U90 ( .B1(n192), .B2(n43), .A(n47), .ZN(n228) );
  NAND2_X1 U91 ( .A1(cansaveNext[2]), .A2(n266), .ZN(n47) );
  OAI21_X1 U92 ( .B1(n65), .B2(n43), .A(n51), .ZN(n225) );
  NAND2_X1 U93 ( .A1(nextState[1]), .A2(n266), .ZN(n51) );
  OAI21_X1 U94 ( .B1(n214), .B2(n43), .A(n54), .ZN(n222) );
  NAND2_X1 U95 ( .A1(canrestoreNext[1]), .A2(n266), .ZN(n54) );
  NOR3_X1 U96 ( .A1(n65), .A2(n66), .A3(n251), .ZN(n110) );
  NOR3_X1 U97 ( .A1(n251), .A2(n66), .A3(n265), .ZN(n80) );
  NOR3_X1 U98 ( .A1(n251), .A2(n65), .A3(n261), .ZN(n150) );
  OAI22_X1 U99 ( .A1(actual_round[0]), .A2(n255), .B1(N466), .B2(n63), .ZN(n67) );
  NOR3_X1 U100 ( .A1(n96), .A2(n6), .A3(n262), .ZN(n148) );
  OAI22_X1 U101 ( .A1(n73), .A2(n264), .B1(n133), .B2(n243), .ZN(n121) );
  XNOR2_X1 U102 ( .A(n240), .B(n129), .ZN(n124) );
  AOI22_X1 U103 ( .A1(n240), .A2(n126), .B1(n235), .B2(n127), .ZN(n125) );
  AOI22_X1 U104 ( .A1(cwpOut[3]), .A2(n79), .B1(n130), .B2(n8), .ZN(n129) );
  OAI21_X1 U105 ( .B1(n89), .B2(n239), .A(n90), .ZN(n88) );
  INV_X1 U106 ( .A(n91), .ZN(n239) );
  OAI21_X1 U107 ( .B1(n91), .B2(n238), .A(n4), .ZN(n90) );
  OAI21_X1 U108 ( .B1(n73), .B2(n248), .A(n147), .ZN(n78) );
  NAND2_X1 U109 ( .A1(cwpOut[0]), .A2(n79), .ZN(n147) );
  NAND4_X1 U110 ( .A1(n146), .A2(n150), .A3(n101), .A4(n107), .ZN(n151) );
  NOR2_X1 U111 ( .A1(n259), .A2(n214), .ZN(n87) );
  AOI22_X1 U112 ( .A1(n159), .A2(swpOut[2]), .B1(n67), .B2(n158), .ZN(n68) );
  NOR2_X1 U113 ( .A1(n270), .A2(call), .ZN(n146) );
  OAI21_X1 U114 ( .B1(n192), .B2(n248), .A(n135), .ZN(n128) );
  NAND2_X1 U115 ( .A1(cwpOut[2]), .A2(n79), .ZN(n135) );
  NAND4_X1 U116 ( .A1(n103), .A2(call), .A3(n107), .A4(n270), .ZN(n111) );
  OAI221_X1 U117 ( .B1(n100), .B2(n250), .C1(n246), .C2(n101), .A(n102), .ZN(
        N450) );
  AOI211_X1 U118 ( .C1(n103), .C2(n104), .A(n157), .B(n105), .ZN(n102) );
  OAI21_X1 U119 ( .B1(n269), .B2(n258), .A(n106), .ZN(n104) );
  NOR3_X1 U120 ( .A1(n265), .A2(n205), .A3(MMUStrobe), .ZN(n105) );
  OAI21_X1 U121 ( .B1(n264), .B2(n248), .A(n141), .ZN(n137) );
  NAND2_X1 U122 ( .A1(cwpOut[1]), .A2(n79), .ZN(n141) );
  OAI221_X1 U123 ( .B1(n112), .B2(n270), .C1(n100), .C2(n250), .A(n113), .ZN(
        N448) );
  NOR2_X1 U124 ( .A1(n114), .A2(n110), .ZN(n112) );
  AOI22_X1 U125 ( .A1(reset), .A2(n80), .B1(n159), .B2(n271), .ZN(n113) );
  AOI21_X1 U126 ( .B1(n249), .B2(n115), .A(call), .ZN(n114) );
  OAI221_X1 U127 ( .B1(n117), .B2(n139), .C1(n248), .C2(n77), .A(n245), .ZN(
        N444) );
  AOI221_X1 U128 ( .B1(n133), .B2(n122), .C1(n143), .C2(n156), .A(n144), .ZN(
        n139) );
  XNOR2_X1 U129 ( .A(n243), .B(n73), .ZN(n143) );
  NOR3_X1 U130 ( .A1(n122), .A2(n156), .A3(n73), .ZN(n144) );
  NAND2_X1 U131 ( .A1(ret), .A2(n107), .ZN(n149) );
  NOR2_X1 U132 ( .A1(n263), .A2(n156), .ZN(n133) );
  NOR3_X1 U133 ( .A1(n247), .A2(n4), .A3(n257), .ZN(n84) );
  NAND4_X1 U134 ( .A1(n66), .A2(n205), .A3(n101), .A4(n107), .ZN(n115) );
  OAI22_X1 U135 ( .A1(n92), .A2(n262), .B1(n4), .B2(n93), .ZN(N453) );
  AOI22_X1 U136 ( .A1(n237), .A2(n83), .B1(n95), .B2(n87), .ZN(n92) );
  AOI22_X1 U137 ( .A1(n94), .A2(n83), .B1(n95), .B2(n257), .ZN(n93) );
  INV_X1 U138 ( .A(n94), .ZN(n237) );
  OAI22_X1 U139 ( .A1(n81), .A2(n260), .B1(n6), .B2(n82), .ZN(N454) );
  AOI21_X1 U140 ( .B1(n85), .B2(n83), .A(n86), .ZN(n81) );
  AOI21_X1 U141 ( .B1(n236), .B2(n83), .A(n84), .ZN(n82) );
  AOI21_X1 U142 ( .B1(n87), .B2(n262), .A(n247), .ZN(n86) );
  OAI22_X1 U143 ( .A1(n75), .A2(n248), .B1(n117), .B2(n118), .ZN(N446) );
  XNOR2_X1 U144 ( .A(n243), .B(n8), .ZN(n120) );
  OAI21_X1 U145 ( .B1(n121), .B2(n122), .A(n123), .ZN(n119) );
  OAI22_X1 U146 ( .A1(n248), .A2(n76), .B1(n117), .B2(n131), .ZN(N445) );
  XNOR2_X1 U147 ( .A(n121), .B(n132), .ZN(n131) );
  XNOR2_X1 U148 ( .A(n192), .B(n122), .ZN(n132) );
  NAND2_X1 U149 ( .A1(enable), .A2(n267), .ZN(n50) );
  NAND2_X1 U150 ( .A1(swpOut[1]), .A2(swpOut[0]), .ZN(n63) );
  INV_X1 U151 ( .A(call), .ZN(n268) );
  INV_X1 U152 ( .A(MMUStrobe), .ZN(n271) );
  NAND4_X1 U153 ( .A1(n74), .A2(call), .A3(n116), .A4(ret), .ZN(N447) );
  NOR2_X1 U154 ( .A1(n80), .A2(n265), .ZN(n116) );
  XNOR2_X1 U155 ( .A(actual_round[1]), .B(n67), .ZN(n62) );
  OAI21_X1 U156 ( .B1(n242), .B2(n243), .A(n192), .ZN(n123) );
  INV_X1 U157 ( .A(n121), .ZN(n242) );
  AND2_X1 U158 ( .A1(n153), .A2(n258), .ZN(n100) );
  NAND2_X1 U159 ( .A1(\need_to_fill[0] ), .A2(n149), .ZN(n153) );
  NAND2_X1 U160 ( .A1(\need_to_spill[0] ), .A2(n268), .ZN(n101) );
  NAND2_X1 U161 ( .A1(n214), .A2(n259), .ZN(n96) );
  AOI21_X1 U162 ( .B1(n99), .B2(n249), .A(n9), .ZN(N451) );
  OAI21_X1 U163 ( .B1(swpOut[0]), .B2(n72), .A(n245), .ZN(N461) );
  INV_X1 U164 ( .A(ret), .ZN(n270) );
  OR3_X1 U165 ( .A1(swpOut[0]), .A2(swpOut[1]), .A3(n252), .ZN(n219) );
  INV_X1 U166 ( .A(reset), .ZN(n267) );
  OR3_X1 U167 ( .A1(n107), .A2(ret), .A3(n268), .ZN(n106) );
  NAND2_X1 U168 ( .A1(n58), .A2(n245), .ZN(N464) );
  XNOR2_X1 U169 ( .A(n59), .B(n60), .ZN(n58) );
  AOI22_X1 U170 ( .A1(n61), .A2(n158), .B1(swpOut[3]), .B2(n159), .ZN(n59) );
  AOI22_X1 U171 ( .A1(n62), .A2(n63), .B1(n255), .B2(n64), .ZN(n61) );
  NAND2_X1 U172 ( .A1(n245), .A2(n69), .ZN(N462) );
  OAI21_X1 U173 ( .B1(n70), .B2(n252), .A(n71), .ZN(n69) );
  OAI21_X1 U174 ( .B1(n70), .B2(n254), .A(n252), .ZN(n71) );
  XNOR2_X1 U175 ( .A(swpOut[1]), .B(swpOut[0]), .ZN(n70) );
  INV_X1 U176 ( .A(n219), .ZN(n231) );
endmodule



    module translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 ( 
        clk, reset, enable, rd1, rd2, wr, add_wr, add_rd1, add_rd2, cwp, 
        add_wr_out, add_rd1_out, add_rd2_out );
  input [4:0] add_wr;
  input [4:0] add_rd1;
  input [4:0] add_rd2;
  input [3:0] cwp;
  output [6:0] add_wr_out;
  output [6:0] add_rd1_out;
  output [6:0] add_rd2_out;
  input clk, reset, enable, rd1, rd2, wr;
  wire   N23, N46, N47, N48, N49, N50, N78, N94, N95, N96, N97, N98, N124,
         N125, N126, N127, N128, N133, N182, N187, N192, \r31/B_AS[4] ,
         \r31/B_AS[3] , \r31/carry[4] , \r31/carry[5] , \r186/B_AS[4] ,
         \r186/B_AS[3] , \r186/carry[4] , \r186/carry[5] , \r32/B_AS[4] ,
         \r32/carry[4] , \r32/carry[5] , n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45;
  assign N23 = add_wr[4];
  assign N46 = add_wr[0];
  assign N47 = add_wr[1];
  assign N48 = add_wr[2];
  assign N78 = add_rd1[4];
  assign N94 = add_rd1[0];
  assign N95 = add_rd1[1];
  assign N96 = add_rd1[2];
  assign N124 = add_rd2[0];
  assign N125 = add_rd2[1];
  assign N126 = add_rd2[2];
  assign N133 = add_rd2[4];
  assign N182 = add_wr[3];
  assign N187 = add_rd1[3];
  assign N192 = add_rd2[3];

  FA_X1 \r31/U1_3  ( .A(N192), .B(\r31/B_AS[3] ), .CI(n38), .CO(\r31/carry[4] ), .S(N127) );
  FA_X1 \r31/U1_4  ( .A(N133), .B(\r31/B_AS[4] ), .CI(\r31/carry[4] ), .CO(
        \r31/carry[5] ), .S(N128) );
  FA_X1 \r186/U1_3  ( .A(N182), .B(\r186/B_AS[3] ), .CI(n39), .CO(
        \r186/carry[4] ), .S(N49) );
  FA_X1 \r186/U1_4  ( .A(N23), .B(\r186/B_AS[4] ), .CI(\r186/carry[4] ), .CO(
        \r186/carry[5] ), .S(N50) );
  FA_X1 \r32/U1_3  ( .A(N187), .B(n37), .CI(n30), .CO(\r32/carry[4] ), .S(N97)
         );
  FA_X1 \r32/U1_4  ( .A(N78), .B(\r32/B_AS[4] ), .CI(\r32/carry[4] ), .CO(
        \r32/carry[5] ), .S(N98) );
  NOR2_X2 U9 ( .A1(n17), .A2(n33), .ZN(add_wr_out[6]) );
  NAND3_X1 U56 ( .A1(n20), .A2(n42), .A3(N23), .ZN(n16) );
  NAND3_X1 U57 ( .A1(n20), .A2(n45), .A3(N133), .ZN(n15) );
  XOR2_X1 U58 ( .A(n27), .B(n30), .Z(n26) );
  NOR2_X1 U3 ( .A1(n22), .A2(n33), .ZN(add_rd2_out[6]) );
  NOR2_X1 U4 ( .A1(n26), .A2(n33), .ZN(add_rd1_out[6]) );
  XNOR2_X1 U5 ( .A(n39), .B(n18), .ZN(n17) );
  NOR2_X1 U6 ( .A1(n19), .A2(n35), .ZN(n18) );
  XNOR2_X1 U7 ( .A(n38), .B(n23), .ZN(n22) );
  NOR2_X1 U8 ( .A1(n24), .A2(n34), .ZN(n23) );
  NAND2_X1 U10 ( .A1(\r32/carry[5] ), .A2(n40), .ZN(n27) );
  NOR2_X1 U11 ( .A1(n33), .A2(n21), .ZN(add_wr_out[5]) );
  XNOR2_X1 U12 ( .A(n35), .B(n19), .ZN(n21) );
  NOR2_X1 U13 ( .A1(n33), .A2(n25), .ZN(add_rd2_out[5]) );
  XNOR2_X1 U14 ( .A(n34), .B(n24), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n33), .A2(n28), .ZN(add_rd1_out[5]) );
  XNOR2_X1 U16 ( .A(\r32/carry[5] ), .B(n40), .ZN(n28) );
  AND2_X1 U17 ( .A1(N50), .A2(enable), .ZN(add_wr_out[4]) );
  AND2_X1 U18 ( .A1(N128), .A2(enable), .ZN(add_rd2_out[4]) );
  AND2_X1 U19 ( .A1(N98), .A2(enable), .ZN(add_rd1_out[4]) );
  AND2_X1 U20 ( .A1(N127), .A2(enable), .ZN(add_rd2_out[3]) );
  AND2_X1 U21 ( .A1(N97), .A2(enable), .ZN(add_rd1_out[3]) );
  AND2_X1 U22 ( .A1(N49), .A2(enable), .ZN(add_wr_out[3]) );
  INV_X1 U23 ( .A(n15), .ZN(n38) );
  INV_X1 U24 ( .A(n16), .ZN(n39) );
  INV_X1 U25 ( .A(\r31/carry[5] ), .ZN(n34) );
  INV_X1 U26 ( .A(\r186/carry[5] ), .ZN(n35) );
  AND2_X1 U27 ( .A1(N94), .A2(enable), .ZN(add_rd1_out[0]) );
  AND2_X1 U28 ( .A1(N125), .A2(enable), .ZN(add_rd2_out[1]) );
  AND2_X1 U29 ( .A1(N95), .A2(enable), .ZN(add_rd1_out[1]) );
  AND2_X1 U30 ( .A1(N126), .A2(enable), .ZN(add_rd2_out[2]) );
  AND2_X1 U31 ( .A1(N96), .A2(enable), .ZN(add_rd1_out[2]) );
  AND2_X1 U32 ( .A1(N124), .A2(enable), .ZN(add_rd2_out[0]) );
  AOI21_X1 U33 ( .B1(N133), .B2(N192), .A(cwp[1]), .ZN(n24) );
  AOI21_X1 U34 ( .B1(N182), .B2(N23), .A(cwp[1]), .ZN(n19) );
  OAI21_X1 U35 ( .B1(n44), .B2(n45), .A(n15), .ZN(\r31/B_AS[3] ) );
  INV_X1 U36 ( .A(N133), .ZN(n44) );
  OAI21_X1 U37 ( .B1(n42), .B2(n41), .A(n16), .ZN(\r186/B_AS[3] ) );
  INV_X1 U38 ( .A(N23), .ZN(n41) );
  NOR2_X1 U39 ( .A1(n37), .A2(n36), .ZN(\r32/B_AS[4] ) );
  AND2_X1 U40 ( .A1(N46), .A2(enable), .ZN(add_wr_out[0]) );
  AND2_X1 U41 ( .A1(N47), .A2(enable), .ZN(add_wr_out[1]) );
  AND3_X1 U42 ( .A1(N78), .A2(n43), .A3(n20), .ZN(n30) );
  INV_X1 U43 ( .A(N187), .ZN(n43) );
  INV_X1 U44 ( .A(cwp[0]), .ZN(n36) );
  NOR2_X1 U45 ( .A1(\r31/B_AS[3] ), .A2(n36), .ZN(\r31/B_AS[4] ) );
  NOR2_X1 U46 ( .A1(\r186/B_AS[3] ), .A2(n36), .ZN(\r186/B_AS[4] ) );
  AND2_X1 U47 ( .A1(N48), .A2(enable), .ZN(add_wr_out[2]) );
  INV_X1 U48 ( .A(n29), .ZN(n40) );
  AOI21_X1 U49 ( .B1(N187), .B2(N78), .A(cwp[1]), .ZN(n29) );
  AND2_X1 U50 ( .A1(cwp[1]), .A2(cwp[0]), .ZN(n20) );
  INV_X1 U51 ( .A(n14), .ZN(n37) );
  AOI21_X1 U52 ( .B1(N187), .B2(N78), .A(n30), .ZN(n14) );
  INV_X1 U53 ( .A(N192), .ZN(n45) );
  INV_X1 U54 ( .A(N182), .ZN(n42) );
  INV_X1 U55 ( .A(enable), .ZN(n33) );
endmodule


module physical_RF_NData32_NRegs72_NAddr7 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [6:0] ADD_WR;
  input [6:0] ADD_RD1;
  input [6:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n97, n98, n99, n578, n580, n582, n584, n586, n588, n590,
         n592, n594, n596, n598, n600, n602, n604, n606, n608, n610, n612,
         n614, n616, n622, n625, n628, n631, n634, n637, n640, n643, n646,
         n649, n652, n653, n655, n656, n658, n659, n661, n662, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n716, n717, n719, n720, n722, n723,
         n725, n726, n728, n729, n731, n732, n734, n735, n737, n738, n740,
         n741, n743, n744, n746, n747, n749, n750, n752, n753, n755, n756,
         n758, n759, n761, n762, n764, n765, n767, n768, n770, n771, n773,
         n774, n776, n777, n779, n780, n782, n783, n785, n786, n788, n789,
         n791, n792, n794, n795, n797, n798, n800, n801, n803, n804, n806,
         n807, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n5383, n5385, n5387, n5393, n5395, n5397, n5403,
         n5405, n5407, n5413, n5415, n5417, n5423, n5425, n5427, n5433, n5435,
         n5437, n5443, n5445, n5447, n5452, n5453, n5455, n5457, n5462, n5463,
         n5465, n5467, n5472, n5473, n5475, n5477, n5482, n5483, n5485, n5487,
         n5492, n5493, n5495, n5497, n5502, n5503, n5505, n5507, n5512, n5513,
         n5515, n5517, n5522, n5523, n5525, n5527, n5532, n5533, n5535, n5537,
         n5542, n5543, n5545, n5547, n5552, n5553, n5555, n5557, n5562, n5563,
         n5565, n5567, n5572, n5573, n5575, n5577, n5582, n5583, n5585, n5587,
         n5592, n5593, n5595, n5597, n5602, n5603, n5605, n5607, n5612, n5613,
         n5615, n5617, n5622, n5623, n5625, n5627, n5632, n5633, n5635, n5637,
         n5642, n5643, n5645, n5647, n5652, n5653, n5655, n5657, n5662, n5663,
         n5665, n5667, n5672, n5673, n5675, n5677, n5682, n5683, n5685, n5687,
         n5692, n5693, n5695, n5697, n5699, n5701, n5703, n5705, n5707, n5709,
         n5711, n5713, n5715, n5717, n5719, n5721, n5723, n5725, n5727, n5729,
         n5731, n5733, n5735, n5737, n5739, n5741, n5743, n5745, n5747, n5749,
         n5751, n5753, n5755, n5757, n5759, n5761, n5763, n5765, n5767, n5769,
         n5771, n5773, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5822, n5824,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6659, n6661, n6663, n6665, n6667, n6669, n6671, n6673,
         n6675, n6677, n6679, n6681, n6683, n6685, n6687, n6689, n6691, n6693,
         n6695, n6697, n6699, n6701, n6703, n6705, n6707, n6709, n6711, n6713,
         n6715, n6717, n6719, n6721, n6723, n6725, n6727, n6729, n6731, n6733,
         n6735, n6737, n6739, n6741, n6743, n6745, n6747, n6749, n6751, n6753,
         n6755, n6757, n6759, n6761, n6763, n6765, n6767, n6769, n6771, n6773,
         n6775, n6777, n6779, n6781, n6783, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5384, n5386, n5388, n5389, n5390,
         n5391, n5392, n5394, n5396, n5398, n5399, n5400, n5401, n5402, n5404,
         n5406, n5408, n5409, n5410, n5411, n5412, n5414, n5416, n5418, n5419,
         n5420, n5421, n5422, n5424, n5426, n5428, n5429, n5430, n5431, n5432,
         n5434, n5436, n5438, n5439, n5440, n5441, n5442, n5444, n5446, n5448,
         n5449, n5450, n5451, n5454, n5456, n5458, n5459, n5460, n5461, n5464,
         n5466, n5468, n5469, n5470, n5471, n5474, n5476, n5478, n5479, n5480,
         n5481, n5484, n5486, n5488, n5489, n5490, n5491, n5494, n5496, n5498,
         n5499, n5500, n5501, n5504, n5506, n5508, n5509, n5510, n5511, n5514,
         n5516, n5518, n5519, n5520, n5521, n5524, n5526, n5528, n5529, n5530,
         n5531, n5534, n5536, n5538, n5539, n5540, n5541, n5544, n5546, n5548,
         n5549, n5550, n5551, n5554, n5556, n5558, n5559, n5560, n5561, n5564,
         n5566, n5568, n5569, n5570, n5571, n5574, n5576, n5578, n5579, n5580,
         n5581, n5584, n5586, n5588, n5589, n5590, n5591, n5594, n5596, n5598,
         n5599, n5600, n5601, n5604, n5606, n5608, n5609, n5610, n5611, n5614,
         n5616, n5618, n5619, n5620, n5621, n5624, n5626, n5628, n5629, n5630,
         n5631, n5634, n5636, n5638, n5639, n5640, n5641, n5644, n5646, n5648,
         n5649, n5650, n5651, n5654, n5656, n5658, n5659, n5660, n5661, n5664,
         n5666, n5668, n5669, n5670, n5671, n5674, n5676, n5678, n5679, n5680,
         n5681, n5684, n5686, n5688, n5689, n5690, n5691, n5694, n5696, n5698,
         n5700, n5702, n5704, n5706, n5708, n5710, n5712, n5714, n5716, n5718,
         n5720, n5722, n5724, n5726, n5728, n5730, n5732, n5734, n5736, n5738,
         n5740, n5742, n5744, n5746, n5748, n5750, n5752, n5754, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107;
  tri   [31:0] OUT1;
  tri   [31:0] OUT2;

  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n9913), .CK(CLK), .Q(n714), .QN(n12648)
         );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n9912), .CK(CLK), .Q(n717), .QN(n12647)
         );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n9911), .CK(CLK), .Q(n720), .QN(n12646)
         );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n9910), .CK(CLK), .Q(n723), .QN(n12645)
         );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n9909), .CK(CLK), .Q(n726), .QN(n12652)
         );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n9908), .CK(CLK), .Q(n729), .QN(n12651)
         );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n9907), .CK(CLK), .Q(n732), .QN(n12650)
         );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n9906), .CK(CLK), .Q(n735), .QN(n12649)
         );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n9905), .CK(CLK), .Q(n738), .QN(n12708)
         );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n9904), .CK(CLK), .Q(n741), .QN(n12706)
         );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n9903), .CK(CLK), .Q(n744), .QN(n12704)
         );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n9902), .CK(CLK), .Q(n747), .QN(n12702)
         );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n9901), .CK(CLK), .Q(n750), .QN(n12700)
         );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n9900), .CK(CLK), .Q(n753), .QN(n12698)
         );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n9899), .CK(CLK), .Q(n756), .QN(n12696)
         );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n9898), .CK(CLK), .Q(n759), .QN(n12694)
         );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n9897), .CK(CLK), .Q(n762), .QN(n12692)
         );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n9896), .CK(CLK), .Q(n765), .QN(n12690)
         );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n9895), .CK(CLK), .Q(n768), .QN(n12688)
         );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n9894), .CK(CLK), .Q(n771), .QN(n12686)
         );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n9893), .CK(CLK), .Q(n774), .QN(n12684)
         );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n9892), .CK(CLK), .Q(n777), .QN(n12682)
         );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n9891), .CK(CLK), .Q(n780), .QN(n12680) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n9890), .CK(CLK), .Q(n783), .QN(n12678) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n9889), .CK(CLK), .Q(n786), .QN(n12676) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n9888), .CK(CLK), .Q(n789), .QN(n12674) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n9887), .CK(CLK), .Q(n792), .QN(n12672) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n9886), .CK(CLK), .Q(n795), .QN(n12670) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n9885), .CK(CLK), .Q(n798), .QN(n12668) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n9884), .CK(CLK), .Q(n801), .QN(n12666) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n9883), .CK(CLK), .Q(n804), .QN(n12664) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n9882), .CK(CLK), .Q(n807), .QN(n12662) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n9785), .CK(CLK), .QN(n14108) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n9784), .CK(CLK), .QN(n14109) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n9783), .CK(CLK), .QN(n14110) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n9782), .CK(CLK), .QN(n14111) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n9781), .CK(CLK), .QN(n14112) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n9780), .CK(CLK), .QN(n14113) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n9779), .CK(CLK), .QN(n14114) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n9778), .CK(CLK), .QN(n14115) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n9777), .CK(CLK), .QN(n14116) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n9776), .CK(CLK), .QN(n14117) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n9775), .CK(CLK), .QN(n14118) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n9774), .CK(CLK), .QN(n14119) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n9773), .CK(CLK), .QN(n14120) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n9772), .CK(CLK), .QN(n14121) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n9771), .CK(CLK), .QN(n14122) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n9770), .CK(CLK), .QN(n14123) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n9769), .CK(CLK), .QN(n14124) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n9768), .CK(CLK), .QN(n14125) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n9767), .CK(CLK), .QN(n14126) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n9766), .CK(CLK), .QN(n14127) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n9765), .CK(CLK), .QN(n14128) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n9764), .CK(CLK), .QN(n14129) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n9763), .CK(CLK), .QN(n14130) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n9762), .CK(CLK), .QN(n14131) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n9761), .CK(CLK), .QN(n14132) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n9760), .CK(CLK), .QN(n14133) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n9759), .CK(CLK), .QN(n14134) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n9758), .CK(CLK), .QN(n14135) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n9757), .CK(CLK), .QN(n14136) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n9756), .CK(CLK), .QN(n14137) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n9755), .CK(CLK), .QN(n14138) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n9754), .CK(CLK), .QN(n14139) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n9753), .CK(CLK), .QN(n14140) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n9752), .CK(CLK), .QN(n14141) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n9751), .CK(CLK), .QN(n14142) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n9750), .CK(CLK), .QN(n14143) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n9749), .CK(CLK), .QN(n14144) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n9748), .CK(CLK), .QN(n14145) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n9747), .CK(CLK), .QN(n14146) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n9746), .CK(CLK), .QN(n14147) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n9745), .CK(CLK), .QN(n14148) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n9744), .CK(CLK), .QN(n14149) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n9743), .CK(CLK), .QN(n14150) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n9742), .CK(CLK), .QN(n14151) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n9741), .CK(CLK), .QN(n14152) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n9740), .CK(CLK), .QN(n14153) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n9739), .CK(CLK), .QN(n14154) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n9738), .CK(CLK), .QN(n14155) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n9737), .CK(CLK), .QN(n14156) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n9736), .CK(CLK), .QN(n14157) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n9735), .CK(CLK), .QN(n14158) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n9734), .CK(CLK), .QN(n14159) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n9733), .CK(CLK), .QN(n14160) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n9732), .CK(CLK), .QN(n14161) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n9731), .CK(CLK), .QN(n14162) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n9730), .CK(CLK), .QN(n14163) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n9729), .CK(CLK), .QN(n14164) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n9728), .CK(CLK), .QN(n14165) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n9727), .CK(CLK), .QN(n14166) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n9726), .CK(CLK), .QN(n14167) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n9725), .CK(CLK), .QN(n14168) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n9724), .CK(CLK), .QN(n14169) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n9723), .CK(CLK), .QN(n14170) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n9722), .CK(CLK), .QN(n14171) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n9721), .CK(CLK), .QN(n14172) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n9720), .CK(CLK), .QN(n14173) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n9719), .CK(CLK), .QN(n14174) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n9718), .CK(CLK), .QN(n14175) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n9717), .CK(CLK), .QN(n14176) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n9716), .CK(CLK), .QN(n14177) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n9715), .CK(CLK), .QN(n14178) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n9714), .CK(CLK), .QN(n14179) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n9713), .CK(CLK), .QN(n14180) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n9712), .CK(CLK), .QN(n14181) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n9711), .CK(CLK), .QN(n14182) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n9710), .CK(CLK), .QN(n14183) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n9709), .CK(CLK), .QN(n14184) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n9708), .CK(CLK), .QN(n14185) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n9707), .CK(CLK), .QN(n14186) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n9706), .CK(CLK), .QN(n14187) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n9705), .CK(CLK), .QN(n14188) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n9704), .CK(CLK), .QN(n14189) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n9703), .CK(CLK), .QN(n14190) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n9702), .CK(CLK), .QN(n14191) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n9701), .CK(CLK), .QN(n14192) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n9700), .CK(CLK), .QN(n14193) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n9699), .CK(CLK), .QN(n14194) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n9698), .CK(CLK), .QN(n14195) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n9697), .CK(CLK), .QN(n14196) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n9696), .CK(CLK), .QN(n14197) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n9695), .CK(CLK), .QN(n14198) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n9694), .CK(CLK), .QN(n14199) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n9693), .CK(CLK), .QN(n14200) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n9692), .CK(CLK), .QN(n14201) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n9691), .CK(CLK), .QN(n14202) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n9690), .CK(CLK), .QN(n14203) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n9625), .CK(CLK), .Q(n713), .QN(n12656)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n9624), .CK(CLK), .Q(n716), .QN(n12655)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n9623), .CK(CLK), .Q(n719), .QN(n12654)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n9622), .CK(CLK), .Q(n722), .QN(n12653)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n9621), .CK(CLK), .Q(n725), .QN(n12660)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n9620), .CK(CLK), .Q(n728), .QN(n12659)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n9619), .CK(CLK), .Q(n731), .QN(n12658)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n9618), .CK(CLK), .Q(n734), .QN(n12657)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n9617), .CK(CLK), .Q(n737), .QN(n12707)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n9616), .CK(CLK), .Q(n740), .QN(n12705)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n9615), .CK(CLK), .Q(n743), .QN(n12703)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n9614), .CK(CLK), .Q(n746), .QN(n12701)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n9613), .CK(CLK), .Q(n749), .QN(n12699)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n9612), .CK(CLK), .Q(n752), .QN(n12697)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n9611), .CK(CLK), .Q(n755), .QN(n12695)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n9610), .CK(CLK), .Q(n758), .QN(n12693)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n9609), .CK(CLK), .Q(n761), .QN(n12691)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n9608), .CK(CLK), .Q(n764), .QN(n12689)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n9607), .CK(CLK), .Q(n767), .QN(n12687)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n9606), .CK(CLK), .Q(n770), .QN(n12685)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n9605), .CK(CLK), .Q(n773), .QN(n12683)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n9604), .CK(CLK), .Q(n776), .QN(n12681)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n9603), .CK(CLK), .Q(n779), .QN(n12679)
         );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n9602), .CK(CLK), .Q(n782), .QN(n12677)
         );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n9601), .CK(CLK), .Q(n785), .QN(n12675)
         );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n9600), .CK(CLK), .Q(n788), .QN(n12673)
         );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n9599), .CK(CLK), .Q(n791), .QN(n12671)
         );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n9598), .CK(CLK), .Q(n794), .QN(n12669)
         );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n9597), .CK(CLK), .Q(n797), .QN(n12667)
         );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n9596), .CK(CLK), .Q(n800), .QN(n12665)
         );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n9595), .CK(CLK), .Q(n803), .QN(n12663)
         );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n9594), .CK(CLK), .Q(n806), .QN(n12661)
         );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n9497), .CK(CLK), .QN(n14280) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n9496), .CK(CLK), .QN(n14281) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n9495), .CK(CLK), .QN(n14282) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n9494), .CK(CLK), .QN(n14283) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n9493), .CK(CLK), .QN(n14284) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n9492), .CK(CLK), .QN(n14285) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n9491), .CK(CLK), .QN(n14286) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n9490), .CK(CLK), .QN(n14287) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n9489), .CK(CLK), .QN(n14288) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n9488), .CK(CLK), .QN(n14289) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n9487), .CK(CLK), .QN(n14290) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n9486), .CK(CLK), .QN(n14291) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n9485), .CK(CLK), .QN(n14292) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n9484), .CK(CLK), .QN(n14293) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n9483), .CK(CLK), .QN(n14294) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n9482), .CK(CLK), .QN(n14295) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n9481), .CK(CLK), .QN(n14296) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n9480), .CK(CLK), .QN(n14297) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n9479), .CK(CLK), .QN(n14298) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n9478), .CK(CLK), .QN(n14299) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n9477), .CK(CLK), .QN(n14300) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n9476), .CK(CLK), .QN(n14301) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n9475), .CK(CLK), .QN(n14302) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n9474), .CK(CLK), .QN(n14303) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n9473), .CK(CLK), .QN(n14304) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n9472), .CK(CLK), .QN(n14305) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n9471), .CK(CLK), .QN(n14306) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n9470), .CK(CLK), .QN(n14307) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n9469), .CK(CLK), .QN(n14308) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n9468), .CK(CLK), .QN(n14309) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n9467), .CK(CLK), .QN(n14310) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n9466), .CK(CLK), .QN(n14311) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n9465), .CK(CLK), .QN(n14312) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n9464), .CK(CLK), .QN(n14313) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n9463), .CK(CLK), .QN(n14314) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n9462), .CK(CLK), .QN(n14315) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n9461), .CK(CLK), .QN(n14316) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n9460), .CK(CLK), .QN(n14317) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n9459), .CK(CLK), .QN(n14318) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n9458), .CK(CLK), .QN(n14319) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n9457), .CK(CLK), .QN(n14320) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n9456), .CK(CLK), .QN(n14321) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n9455), .CK(CLK), .QN(n14322) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n9454), .CK(CLK), .QN(n14323) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n9453), .CK(CLK), .QN(n14324) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n9452), .CK(CLK), .QN(n14325) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n9451), .CK(CLK), .QN(n14326) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n9450), .CK(CLK), .QN(n14327) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n9449), .CK(CLK), .QN(n14328) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n9448), .CK(CLK), .QN(n14329) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n9447), .CK(CLK), .QN(n14330) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n9446), .CK(CLK), .QN(n14331) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n9445), .CK(CLK), .QN(n14332) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n9444), .CK(CLK), .QN(n14333) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n9443), .CK(CLK), .QN(n14334) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n9442), .CK(CLK), .QN(n14335) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n9441), .CK(CLK), .QN(n14336) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n9440), .CK(CLK), .QN(n14337) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n9439), .CK(CLK), .QN(n14338) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n9438), .CK(CLK), .QN(n14339) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n9437), .CK(CLK), .QN(n14340) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n9436), .CK(CLK), .QN(n14341) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n9435), .CK(CLK), .QN(n14342) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n9434), .CK(CLK), .QN(n14343) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n9433), .CK(CLK), .QN(n14344) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n9432), .CK(CLK), .QN(n14345) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n9431), .CK(CLK), .QN(n14346) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n9430), .CK(CLK), .QN(n14347) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n9429), .CK(CLK), .QN(n14348) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n9428), .CK(CLK), .QN(n14349) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n9427), .CK(CLK), .QN(n14350) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n9426), .CK(CLK), .QN(n14351) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n9425), .CK(CLK), .QN(n14352) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n9424), .CK(CLK), .QN(n14353) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n9423), .CK(CLK), .QN(n14354) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n9422), .CK(CLK), .QN(n14355) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n9421), .CK(CLK), .QN(n14356) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n9420), .CK(CLK), .QN(n14357) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n9419), .CK(CLK), .QN(n14358) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n9418), .CK(CLK), .QN(n14359) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n9417), .CK(CLK), .QN(n14360) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n9416), .CK(CLK), .QN(n14361) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n9415), .CK(CLK), .QN(n14362) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n9414), .CK(CLK), .QN(n14363) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n9413), .CK(CLK), .QN(n14364) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n9412), .CK(CLK), .QN(n14365) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n9411), .CK(CLK), .QN(n14366) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n9410), .CK(CLK), .QN(n14367) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n9409), .CK(CLK), .QN(n14368) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n9408), .CK(CLK), .QN(n14369) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n9407), .CK(CLK), .QN(n14370) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n9406), .CK(CLK), .QN(n14371) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n9405), .CK(CLK), .QN(n14372) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n9404), .CK(CLK), .QN(n14373) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n9403), .CK(CLK), .QN(n14374) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n9402), .CK(CLK), .QN(n14375) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n9401), .CK(CLK), .QN(n14376) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n9400), .CK(CLK), .QN(n14377) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n9399), .CK(CLK), .QN(n14378) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n9398), .CK(CLK), .QN(n14379) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n9397), .CK(CLK), .QN(n14380) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n9396), .CK(CLK), .QN(n14381) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n9395), .CK(CLK), .QN(n14382) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n9394), .CK(CLK), .QN(n14383) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n9393), .CK(CLK), .QN(n14384) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n9392), .CK(CLK), .QN(n14385) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n9391), .CK(CLK), .QN(n14386) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n9390), .CK(CLK), .QN(n14387) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n9389), .CK(CLK), .QN(n14388) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n9388), .CK(CLK), .QN(n14389) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n9387), .CK(CLK), .QN(n14390) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n9386), .CK(CLK), .QN(n14391) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n9385), .CK(CLK), .QN(n14392) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n9384), .CK(CLK), .QN(n14393) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n9383), .CK(CLK), .QN(n14394) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n9382), .CK(CLK), .QN(n14395) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n9381), .CK(CLK), .QN(n14396) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n9380), .CK(CLK), .QN(n14397) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n9379), .CK(CLK), .QN(n14398) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n9378), .CK(CLK), .QN(n14399) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n9377), .CK(CLK), .QN(n14400) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n9376), .CK(CLK), .QN(n14401) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n9375), .CK(CLK), .QN(n14402) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n9374), .CK(CLK), .QN(n14403) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n9373), .CK(CLK), .QN(n14404) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n9372), .CK(CLK), .QN(n14405) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n9371), .CK(CLK), .QN(n14406) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n9370), .CK(CLK), .QN(n14407) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n9369), .CK(CLK), .QN(n14408) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n9368), .CK(CLK), .QN(n14409) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n9367), .CK(CLK), .QN(n14410) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n9366), .CK(CLK), .QN(n14411) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n9365), .CK(CLK), .QN(n14412) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n9364), .CK(CLK), .QN(n14413) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n9363), .CK(CLK), .QN(n14414) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n9362), .CK(CLK), .QN(n14415) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n9361), .CK(CLK), .QN(n14416) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n9360), .CK(CLK), .QN(n14417) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n9359), .CK(CLK), .QN(n14418) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n9358), .CK(CLK), .QN(n14419) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n9357), .CK(CLK), .QN(n14420) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n9356), .CK(CLK), .QN(n14421) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n9355), .CK(CLK), .QN(n14422) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n9354), .CK(CLK), .QN(n14423) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n9353), .CK(CLK), .QN(n14424) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n9352), .CK(CLK), .QN(n14425) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n9351), .CK(CLK), .QN(n14426) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n9350), .CK(CLK), .QN(n14427) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n9349), .CK(CLK), .QN(n14428) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n9348), .CK(CLK), .QN(n14429) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n9347), .CK(CLK), .QN(n14430) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n9346), .CK(CLK), .QN(n14431) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n9345), .CK(CLK), .QN(n14432) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n9344), .CK(CLK), .QN(n14433) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n9343), .CK(CLK), .QN(n14434) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n9342), .CK(CLK), .QN(n14435) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n9341), .CK(CLK), .QN(n14436) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n9340), .CK(CLK), .QN(n14437) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n9339), .CK(CLK), .QN(n14438) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n9338), .CK(CLK), .QN(n14439) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n9305), .CK(CLK), .Q(n97), .QN(n14459)
         );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n9304), .CK(CLK), .Q(n99), .QN(n14460)
         );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n9209), .CK(CLK), .QN(n14493) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n9208), .CK(CLK), .QN(n14494) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n9207), .CK(CLK), .QN(n14495) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n9206), .CK(CLK), .QN(n14496) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n9205), .CK(CLK), .QN(n14497) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n9204), .CK(CLK), .QN(n14498) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n9203), .CK(CLK), .QN(n14499) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n9202), .CK(CLK), .QN(n14500) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n9201), .CK(CLK), .QN(n14501) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n9200), .CK(CLK), .QN(n14502) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n9199), .CK(CLK), .QN(n14503) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n9198), .CK(CLK), .QN(n14504) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n9197), .CK(CLK), .QN(n14505) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n9196), .CK(CLK), .QN(n14506) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n9195), .CK(CLK), .QN(n14507) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n9194), .CK(CLK), .QN(n14508) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n9193), .CK(CLK), .QN(n14509) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n9192), .CK(CLK), .QN(n14510) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n9191), .CK(CLK), .QN(n14511) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n9190), .CK(CLK), .QN(n14512) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n9189), .CK(CLK), .QN(n14513) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n9188), .CK(CLK), .QN(n14514) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n9187), .CK(CLK), .QN(n14515) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n9186), .CK(CLK), .QN(n14516) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n9185), .CK(CLK), .QN(n14517) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n9184), .CK(CLK), .QN(n14518) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n9183), .CK(CLK), .QN(n14519) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n9182), .CK(CLK), .QN(n14520) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n9181), .CK(CLK), .QN(n14521) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n9180), .CK(CLK), .QN(n14522) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n9179), .CK(CLK), .QN(n14523) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n9178), .CK(CLK), .QN(n14524) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n9177), .CK(CLK), .QN(n14525) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n9176), .CK(CLK), .QN(n14526) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n9175), .CK(CLK), .QN(n14527) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n9174), .CK(CLK), .QN(n14528) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n9173), .CK(CLK), .QN(n14529) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n9172), .CK(CLK), .QN(n14530) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n9171), .CK(CLK), .QN(n14531) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n9170), .CK(CLK), .QN(n14532) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n9169), .CK(CLK), .QN(n14533) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n9168), .CK(CLK), .QN(n14534) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n9167), .CK(CLK), .QN(n14535) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n9166), .CK(CLK), .QN(n14536) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n9165), .CK(CLK), .QN(n14537) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n9164), .CK(CLK), .QN(n14538) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n9163), .CK(CLK), .QN(n14539) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n9162), .CK(CLK), .QN(n14540) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n9161), .CK(CLK), .QN(n14541) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n9160), .CK(CLK), .QN(n14542) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n9159), .CK(CLK), .QN(n14543) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n9158), .CK(CLK), .QN(n14544) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n9157), .CK(CLK), .QN(n14545) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n9156), .CK(CLK), .QN(n14546) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n9155), .CK(CLK), .QN(n14547) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n9154), .CK(CLK), .QN(n14548) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n9153), .CK(CLK), .QN(n14549) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n9152), .CK(CLK), .QN(n14550) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n9151), .CK(CLK), .QN(n14551) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n9150), .CK(CLK), .QN(n14552) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n9149), .CK(CLK), .QN(n14553) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n9148), .CK(CLK), .QN(n14554) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n9147), .CK(CLK), .QN(n14555) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n9146), .CK(CLK), .QN(n14556) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n9145), .CK(CLK), .QN(n14557) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n9144), .CK(CLK), .QN(n14558) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n9143), .CK(CLK), .QN(n14559) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n9142), .CK(CLK), .QN(n14560) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n9141), .CK(CLK), .QN(n14561) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n9140), .CK(CLK), .QN(n14562) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n9139), .CK(CLK), .QN(n14563) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n9138), .CK(CLK), .QN(n14564) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n9137), .CK(CLK), .QN(n14565) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n9136), .CK(CLK), .QN(n14566) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n9135), .CK(CLK), .QN(n14567) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n9134), .CK(CLK), .QN(n14568) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n9133), .CK(CLK), .QN(n14569) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n9132), .CK(CLK), .QN(n14570) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n9131), .CK(CLK), .QN(n14571) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n9130), .CK(CLK), .QN(n14572) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n9129), .CK(CLK), .QN(n14573) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n9128), .CK(CLK), .QN(n14574) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n9127), .CK(CLK), .QN(n14575) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n9126), .CK(CLK), .QN(n14576) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n9125), .CK(CLK), .QN(n14577) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n9124), .CK(CLK), .QN(n14578) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n9123), .CK(CLK), .QN(n14579) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n9122), .CK(CLK), .QN(n14580) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n9121), .CK(CLK), .QN(n14581) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n9120), .CK(CLK), .QN(n14582) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n9119), .CK(CLK), .QN(n14583) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n9118), .CK(CLK), .QN(n14584) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n9117), .CK(CLK), .QN(n14585) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n9116), .CK(CLK), .QN(n14586) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n9115), .CK(CLK), .QN(n14587) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n9114), .CK(CLK), .QN(n14588) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n9113), .CK(CLK), .QN(n14589) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n9112), .CK(CLK), .QN(n14590) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n9111), .CK(CLK), .QN(n14591) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n9110), .CK(CLK), .QN(n14592) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n9109), .CK(CLK), .QN(n14593) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n9108), .CK(CLK), .QN(n14594) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n9107), .CK(CLK), .QN(n14595) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n9106), .CK(CLK), .QN(n14596) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n9105), .CK(CLK), .QN(n14597) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n9104), .CK(CLK), .QN(n14598) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n9103), .CK(CLK), .QN(n14599) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n9102), .CK(CLK), .QN(n14600) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n9101), .CK(CLK), .QN(n14601) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n9100), .CK(CLK), .QN(n14602) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n9099), .CK(CLK), .QN(n14603) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n9098), .CK(CLK), .QN(n14604) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n9097), .CK(CLK), .QN(n14605) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n9096), .CK(CLK), .QN(n14606) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n9095), .CK(CLK), .QN(n14607) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n9094), .CK(CLK), .QN(n14608) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n9093), .CK(CLK), .QN(n14609) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n9092), .CK(CLK), .QN(n14610) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n9091), .CK(CLK), .QN(n14611) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n9090), .CK(CLK), .QN(n14612) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n9089), .CK(CLK), .QN(n14613) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n9088), .CK(CLK), .QN(n14614) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n9087), .CK(CLK), .QN(n14615) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n9086), .CK(CLK), .QN(n14616) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n9085), .CK(CLK), .QN(n14617) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n9084), .CK(CLK), .QN(n14618) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n9083), .CK(CLK), .QN(n14619) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n9082), .CK(CLK), .QN(n14620) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n9081), .CK(CLK), .QN(n14621) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n9080), .CK(CLK), .QN(n14622) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n9079), .CK(CLK), .QN(n14623) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n9078), .CK(CLK), .QN(n14624) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n9077), .CK(CLK), .QN(n14625) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n9076), .CK(CLK), .QN(n14626) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n9075), .CK(CLK), .QN(n14627) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n9074), .CK(CLK), .QN(n14628) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n9073), .CK(CLK), .QN(n14629) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n9072), .CK(CLK), .QN(n14630) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n9071), .CK(CLK), .QN(n14631) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n9070), .CK(CLK), .QN(n14632) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n9069), .CK(CLK), .QN(n14633) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n9068), .CK(CLK), .QN(n14634) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n9067), .CK(CLK), .QN(n14635) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n9066), .CK(CLK), .QN(n14636) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n9065), .CK(CLK), .QN(n14637) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n9064), .CK(CLK), .QN(n14638) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n9063), .CK(CLK), .QN(n14639) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n9062), .CK(CLK), .QN(n14640) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n9061), .CK(CLK), .QN(n14641) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n9060), .CK(CLK), .QN(n14642) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n9059), .CK(CLK), .QN(n14643) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n9058), .CK(CLK), .QN(n14644) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n9057), .CK(CLK), .QN(n14645) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n9056), .CK(CLK), .QN(n14646) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n9055), .CK(CLK), .QN(n14647) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n9054), .CK(CLK), .QN(n14648) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n9053), .CK(CLK), .QN(n14649) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n9052), .CK(CLK), .QN(n14650) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n9051), .CK(CLK), .QN(n14651) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n9050), .CK(CLK), .QN(n14652) );
  DFF_X1 \REGISTERS_reg[33][31]  ( .D(n8921), .CK(CLK), .QN(n14692) );
  DFF_X1 \REGISTERS_reg[33][30]  ( .D(n8920), .CK(CLK), .QN(n14693) );
  DFF_X1 \REGISTERS_reg[33][29]  ( .D(n8919), .CK(CLK), .QN(n14694) );
  DFF_X1 \REGISTERS_reg[33][28]  ( .D(n8918), .CK(CLK), .QN(n14695) );
  DFF_X1 \REGISTERS_reg[33][27]  ( .D(n8917), .CK(CLK), .QN(n14696) );
  DFF_X1 \REGISTERS_reg[33][26]  ( .D(n8916), .CK(CLK), .QN(n14697) );
  DFF_X1 \REGISTERS_reg[33][25]  ( .D(n8915), .CK(CLK), .QN(n14698) );
  DFF_X1 \REGISTERS_reg[33][24]  ( .D(n8914), .CK(CLK), .QN(n14699) );
  DFF_X1 \REGISTERS_reg[33][23]  ( .D(n8913), .CK(CLK), .QN(n14700) );
  DFF_X1 \REGISTERS_reg[33][22]  ( .D(n8912), .CK(CLK), .QN(n14701) );
  DFF_X1 \REGISTERS_reg[33][21]  ( .D(n8911), .CK(CLK), .QN(n14702) );
  DFF_X1 \REGISTERS_reg[33][20]  ( .D(n8910), .CK(CLK), .QN(n14703) );
  DFF_X1 \REGISTERS_reg[33][19]  ( .D(n8909), .CK(CLK), .QN(n14704) );
  DFF_X1 \REGISTERS_reg[33][18]  ( .D(n8908), .CK(CLK), .QN(n14705) );
  DFF_X1 \REGISTERS_reg[33][17]  ( .D(n8907), .CK(CLK), .QN(n14706) );
  DFF_X1 \REGISTERS_reg[33][16]  ( .D(n8906), .CK(CLK), .QN(n14707) );
  DFF_X1 \REGISTERS_reg[33][15]  ( .D(n8905), .CK(CLK), .QN(n14708) );
  DFF_X1 \REGISTERS_reg[33][14]  ( .D(n8904), .CK(CLK), .QN(n14709) );
  DFF_X1 \REGISTERS_reg[33][13]  ( .D(n8903), .CK(CLK), .QN(n14710) );
  DFF_X1 \REGISTERS_reg[33][12]  ( .D(n8902), .CK(CLK), .QN(n14711) );
  DFF_X1 \REGISTERS_reg[33][11]  ( .D(n8901), .CK(CLK), .QN(n14712) );
  DFF_X1 \REGISTERS_reg[33][10]  ( .D(n8900), .CK(CLK), .QN(n14713) );
  DFF_X1 \REGISTERS_reg[33][9]  ( .D(n8899), .CK(CLK), .QN(n14714) );
  DFF_X1 \REGISTERS_reg[33][8]  ( .D(n8898), .CK(CLK), .QN(n14715) );
  DFF_X1 \REGISTERS_reg[33][7]  ( .D(n8897), .CK(CLK), .QN(n14716) );
  DFF_X1 \REGISTERS_reg[33][6]  ( .D(n8896), .CK(CLK), .QN(n14717) );
  DFF_X1 \REGISTERS_reg[33][5]  ( .D(n8895), .CK(CLK), .QN(n14718) );
  DFF_X1 \REGISTERS_reg[33][4]  ( .D(n8894), .CK(CLK), .QN(n14719) );
  DFF_X1 \REGISTERS_reg[33][3]  ( .D(n8893), .CK(CLK), .QN(n14720) );
  DFF_X1 \REGISTERS_reg[33][2]  ( .D(n8892), .CK(CLK), .QN(n14721) );
  DFF_X1 \REGISTERS_reg[33][1]  ( .D(n8891), .CK(CLK), .QN(n14722) );
  DFF_X1 \REGISTERS_reg[33][0]  ( .D(n8890), .CK(CLK), .QN(n14723) );
  DFF_X1 \REGISTERS_reg[34][31]  ( .D(n8889), .CK(CLK), .QN(n14724) );
  DFF_X1 \REGISTERS_reg[34][30]  ( .D(n8888), .CK(CLK), .QN(n14725) );
  DFF_X1 \REGISTERS_reg[34][29]  ( .D(n8887), .CK(CLK), .QN(n14726) );
  DFF_X1 \REGISTERS_reg[34][28]  ( .D(n8886), .CK(CLK), .QN(n14727) );
  DFF_X1 \REGISTERS_reg[34][27]  ( .D(n8885), .CK(CLK), .QN(n14728) );
  DFF_X1 \REGISTERS_reg[34][26]  ( .D(n8884), .CK(CLK), .QN(n14729) );
  DFF_X1 \REGISTERS_reg[34][25]  ( .D(n8883), .CK(CLK), .QN(n14730) );
  DFF_X1 \REGISTERS_reg[34][24]  ( .D(n8882), .CK(CLK), .QN(n14731) );
  DFF_X1 \REGISTERS_reg[34][23]  ( .D(n8881), .CK(CLK), .QN(n14732) );
  DFF_X1 \REGISTERS_reg[34][22]  ( .D(n8880), .CK(CLK), .QN(n14733) );
  DFF_X1 \REGISTERS_reg[34][21]  ( .D(n8879), .CK(CLK), .QN(n14734) );
  DFF_X1 \REGISTERS_reg[34][20]  ( .D(n8878), .CK(CLK), .QN(n14735) );
  DFF_X1 \REGISTERS_reg[34][19]  ( .D(n8877), .CK(CLK), .QN(n14736) );
  DFF_X1 \REGISTERS_reg[34][18]  ( .D(n8876), .CK(CLK), .QN(n14737) );
  DFF_X1 \REGISTERS_reg[34][17]  ( .D(n8875), .CK(CLK), .QN(n14738) );
  DFF_X1 \REGISTERS_reg[34][16]  ( .D(n8874), .CK(CLK), .QN(n14739) );
  DFF_X1 \REGISTERS_reg[34][15]  ( .D(n8873), .CK(CLK), .QN(n14740) );
  DFF_X1 \REGISTERS_reg[34][14]  ( .D(n8872), .CK(CLK), .QN(n14741) );
  DFF_X1 \REGISTERS_reg[34][13]  ( .D(n8871), .CK(CLK), .QN(n14742) );
  DFF_X1 \REGISTERS_reg[34][12]  ( .D(n8870), .CK(CLK), .QN(n14743) );
  DFF_X1 \REGISTERS_reg[34][11]  ( .D(n8869), .CK(CLK), .QN(n14744) );
  DFF_X1 \REGISTERS_reg[34][10]  ( .D(n8868), .CK(CLK), .QN(n14745) );
  DFF_X1 \REGISTERS_reg[34][9]  ( .D(n8867), .CK(CLK), .QN(n14746) );
  DFF_X1 \REGISTERS_reg[34][8]  ( .D(n8866), .CK(CLK), .QN(n14747) );
  DFF_X1 \REGISTERS_reg[34][7]  ( .D(n8865), .CK(CLK), .QN(n14748) );
  DFF_X1 \REGISTERS_reg[34][6]  ( .D(n8864), .CK(CLK), .QN(n14749) );
  DFF_X1 \REGISTERS_reg[34][5]  ( .D(n8863), .CK(CLK), .QN(n14750) );
  DFF_X1 \REGISTERS_reg[34][4]  ( .D(n8862), .CK(CLK), .QN(n14751) );
  DFF_X1 \REGISTERS_reg[34][3]  ( .D(n8861), .CK(CLK), .QN(n14752) );
  DFF_X1 \REGISTERS_reg[34][2]  ( .D(n8860), .CK(CLK), .QN(n14753) );
  DFF_X1 \REGISTERS_reg[34][1]  ( .D(n8859), .CK(CLK), .QN(n14754) );
  DFF_X1 \REGISTERS_reg[34][0]  ( .D(n8858), .CK(CLK), .QN(n14755) );
  DFF_X1 \REGISTERS_reg[35][31]  ( .D(n8857), .CK(CLK), .QN(n14756) );
  DFF_X1 \REGISTERS_reg[35][30]  ( .D(n8856), .CK(CLK), .QN(n14757) );
  DFF_X1 \REGISTERS_reg[35][29]  ( .D(n8855), .CK(CLK), .QN(n14758) );
  DFF_X1 \REGISTERS_reg[35][28]  ( .D(n8854), .CK(CLK), .QN(n14759) );
  DFF_X1 \REGISTERS_reg[35][27]  ( .D(n8853), .CK(CLK), .QN(n14760) );
  DFF_X1 \REGISTERS_reg[35][26]  ( .D(n8852), .CK(CLK), .QN(n14761) );
  DFF_X1 \REGISTERS_reg[35][25]  ( .D(n8851), .CK(CLK), .QN(n14762) );
  DFF_X1 \REGISTERS_reg[35][24]  ( .D(n8850), .CK(CLK), .QN(n14763) );
  DFF_X1 \REGISTERS_reg[35][23]  ( .D(n8849), .CK(CLK), .QN(n14764) );
  DFF_X1 \REGISTERS_reg[35][22]  ( .D(n8848), .CK(CLK), .QN(n14765) );
  DFF_X1 \REGISTERS_reg[35][21]  ( .D(n8847), .CK(CLK), .QN(n14766) );
  DFF_X1 \REGISTERS_reg[35][20]  ( .D(n8846), .CK(CLK), .QN(n14767) );
  DFF_X1 \REGISTERS_reg[35][19]  ( .D(n8845), .CK(CLK), .QN(n14768) );
  DFF_X1 \REGISTERS_reg[35][18]  ( .D(n8844), .CK(CLK), .QN(n14769) );
  DFF_X1 \REGISTERS_reg[35][17]  ( .D(n8843), .CK(CLK), .QN(n14770) );
  DFF_X1 \REGISTERS_reg[35][16]  ( .D(n8842), .CK(CLK), .QN(n14771) );
  DFF_X1 \REGISTERS_reg[35][15]  ( .D(n8841), .CK(CLK), .QN(n14772) );
  DFF_X1 \REGISTERS_reg[35][14]  ( .D(n8840), .CK(CLK), .QN(n14773) );
  DFF_X1 \REGISTERS_reg[35][13]  ( .D(n8839), .CK(CLK), .QN(n14774) );
  DFF_X1 \REGISTERS_reg[35][12]  ( .D(n8838), .CK(CLK), .QN(n14775) );
  DFF_X1 \REGISTERS_reg[35][11]  ( .D(n8837), .CK(CLK), .QN(n14776) );
  DFF_X1 \REGISTERS_reg[35][10]  ( .D(n8836), .CK(CLK), .QN(n14777) );
  DFF_X1 \REGISTERS_reg[35][9]  ( .D(n8835), .CK(CLK), .QN(n14778) );
  DFF_X1 \REGISTERS_reg[35][8]  ( .D(n8834), .CK(CLK), .QN(n14779) );
  DFF_X1 \REGISTERS_reg[35][7]  ( .D(n8833), .CK(CLK), .QN(n14780) );
  DFF_X1 \REGISTERS_reg[35][6]  ( .D(n8832), .CK(CLK), .QN(n14781) );
  DFF_X1 \REGISTERS_reg[35][5]  ( .D(n8831), .CK(CLK), .QN(n14782) );
  DFF_X1 \REGISTERS_reg[35][4]  ( .D(n8830), .CK(CLK), .QN(n14783) );
  DFF_X1 \REGISTERS_reg[35][3]  ( .D(n8829), .CK(CLK), .QN(n14784) );
  DFF_X1 \REGISTERS_reg[35][2]  ( .D(n8828), .CK(CLK), .QN(n14785) );
  DFF_X1 \REGISTERS_reg[35][1]  ( .D(n8827), .CK(CLK), .QN(n14786) );
  DFF_X1 \REGISTERS_reg[35][0]  ( .D(n8826), .CK(CLK), .QN(n14787) );
  DFF_X1 \REGISTERS_reg[36][31]  ( .D(n8825), .CK(CLK), .QN(n14788) );
  DFF_X1 \REGISTERS_reg[36][30]  ( .D(n8824), .CK(CLK), .QN(n14789) );
  DFF_X1 \REGISTERS_reg[36][29]  ( .D(n8823), .CK(CLK), .QN(n14790) );
  DFF_X1 \REGISTERS_reg[36][28]  ( .D(n8822), .CK(CLK), .QN(n14791) );
  DFF_X1 \REGISTERS_reg[36][27]  ( .D(n8821), .CK(CLK), .QN(n14792) );
  DFF_X1 \REGISTERS_reg[36][26]  ( .D(n8820), .CK(CLK), .QN(n14793) );
  DFF_X1 \REGISTERS_reg[36][25]  ( .D(n8819), .CK(CLK), .QN(n14794) );
  DFF_X1 \REGISTERS_reg[36][24]  ( .D(n8818), .CK(CLK), .QN(n14795) );
  DFF_X1 \REGISTERS_reg[36][23]  ( .D(n8817), .CK(CLK), .QN(n14796) );
  DFF_X1 \REGISTERS_reg[36][22]  ( .D(n8816), .CK(CLK), .QN(n14797) );
  DFF_X1 \REGISTERS_reg[36][21]  ( .D(n8815), .CK(CLK), .QN(n14798) );
  DFF_X1 \REGISTERS_reg[36][20]  ( .D(n8814), .CK(CLK), .QN(n14799) );
  DFF_X1 \REGISTERS_reg[36][19]  ( .D(n8813), .CK(CLK), .QN(n14800) );
  DFF_X1 \REGISTERS_reg[36][18]  ( .D(n8812), .CK(CLK), .QN(n14801) );
  DFF_X1 \REGISTERS_reg[36][17]  ( .D(n8811), .CK(CLK), .QN(n14802) );
  DFF_X1 \REGISTERS_reg[36][16]  ( .D(n8810), .CK(CLK), .QN(n14803) );
  DFF_X1 \REGISTERS_reg[36][15]  ( .D(n8809), .CK(CLK), .QN(n14804) );
  DFF_X1 \REGISTERS_reg[36][14]  ( .D(n8808), .CK(CLK), .QN(n14805) );
  DFF_X1 \REGISTERS_reg[36][13]  ( .D(n8807), .CK(CLK), .QN(n14806) );
  DFF_X1 \REGISTERS_reg[36][12]  ( .D(n8806), .CK(CLK), .QN(n14807) );
  DFF_X1 \REGISTERS_reg[36][11]  ( .D(n8805), .CK(CLK), .QN(n14808) );
  DFF_X1 \REGISTERS_reg[36][10]  ( .D(n8804), .CK(CLK), .QN(n14809) );
  DFF_X1 \REGISTERS_reg[36][9]  ( .D(n8803), .CK(CLK), .QN(n14810) );
  DFF_X1 \REGISTERS_reg[36][8]  ( .D(n8802), .CK(CLK), .QN(n14811) );
  DFF_X1 \REGISTERS_reg[36][7]  ( .D(n8801), .CK(CLK), .QN(n14812) );
  DFF_X1 \REGISTERS_reg[36][6]  ( .D(n8800), .CK(CLK), .QN(n14813) );
  DFF_X1 \REGISTERS_reg[36][5]  ( .D(n8799), .CK(CLK), .QN(n14814) );
  DFF_X1 \REGISTERS_reg[36][4]  ( .D(n8798), .CK(CLK), .QN(n14815) );
  DFF_X1 \REGISTERS_reg[36][3]  ( .D(n8797), .CK(CLK), .QN(n14816) );
  DFF_X1 \REGISTERS_reg[36][2]  ( .D(n8796), .CK(CLK), .QN(n14817) );
  DFF_X1 \REGISTERS_reg[36][1]  ( .D(n8795), .CK(CLK), .QN(n14818) );
  DFF_X1 \REGISTERS_reg[36][0]  ( .D(n8794), .CK(CLK), .QN(n14819) );
  DFF_X1 \REGISTERS_reg[37][31]  ( .D(n8793), .CK(CLK), .QN(n14820) );
  DFF_X1 \REGISTERS_reg[37][30]  ( .D(n8792), .CK(CLK), .QN(n14821) );
  DFF_X1 \REGISTERS_reg[37][29]  ( .D(n8791), .CK(CLK), .QN(n14822) );
  DFF_X1 \REGISTERS_reg[37][28]  ( .D(n8790), .CK(CLK), .QN(n14823) );
  DFF_X1 \REGISTERS_reg[37][27]  ( .D(n8789), .CK(CLK), .QN(n14824) );
  DFF_X1 \REGISTERS_reg[37][26]  ( .D(n8788), .CK(CLK), .QN(n14825) );
  DFF_X1 \REGISTERS_reg[37][25]  ( .D(n8787), .CK(CLK), .QN(n14826) );
  DFF_X1 \REGISTERS_reg[37][24]  ( .D(n8786), .CK(CLK), .QN(n14827) );
  DFF_X1 \REGISTERS_reg[37][23]  ( .D(n8785), .CK(CLK), .QN(n14828) );
  DFF_X1 \REGISTERS_reg[37][22]  ( .D(n8784), .CK(CLK), .QN(n14829) );
  DFF_X1 \REGISTERS_reg[37][21]  ( .D(n8783), .CK(CLK), .QN(n14830) );
  DFF_X1 \REGISTERS_reg[37][20]  ( .D(n8782), .CK(CLK), .QN(n14831) );
  DFF_X1 \REGISTERS_reg[37][19]  ( .D(n8781), .CK(CLK), .QN(n14832) );
  DFF_X1 \REGISTERS_reg[37][18]  ( .D(n8780), .CK(CLK), .QN(n14833) );
  DFF_X1 \REGISTERS_reg[37][17]  ( .D(n8779), .CK(CLK), .QN(n14834) );
  DFF_X1 \REGISTERS_reg[37][16]  ( .D(n8778), .CK(CLK), .QN(n14835) );
  DFF_X1 \REGISTERS_reg[37][15]  ( .D(n8777), .CK(CLK), .QN(n14836) );
  DFF_X1 \REGISTERS_reg[37][14]  ( .D(n8776), .CK(CLK), .QN(n14837) );
  DFF_X1 \REGISTERS_reg[37][13]  ( .D(n8775), .CK(CLK), .QN(n14838) );
  DFF_X1 \REGISTERS_reg[37][12]  ( .D(n8774), .CK(CLK), .QN(n14839) );
  DFF_X1 \REGISTERS_reg[37][11]  ( .D(n8773), .CK(CLK), .QN(n14840) );
  DFF_X1 \REGISTERS_reg[37][10]  ( .D(n8772), .CK(CLK), .QN(n14841) );
  DFF_X1 \REGISTERS_reg[37][9]  ( .D(n8771), .CK(CLK), .QN(n14842) );
  DFF_X1 \REGISTERS_reg[37][8]  ( .D(n8770), .CK(CLK), .QN(n14843) );
  DFF_X1 \REGISTERS_reg[37][7]  ( .D(n8769), .CK(CLK), .QN(n14844) );
  DFF_X1 \REGISTERS_reg[37][6]  ( .D(n8768), .CK(CLK), .QN(n14845) );
  DFF_X1 \REGISTERS_reg[37][5]  ( .D(n8767), .CK(CLK), .QN(n14846) );
  DFF_X1 \REGISTERS_reg[37][4]  ( .D(n8766), .CK(CLK), .QN(n14847) );
  DFF_X1 \REGISTERS_reg[37][3]  ( .D(n8765), .CK(CLK), .QN(n14848) );
  DFF_X1 \REGISTERS_reg[37][2]  ( .D(n8764), .CK(CLK), .QN(n14849) );
  DFF_X1 \REGISTERS_reg[37][1]  ( .D(n8763), .CK(CLK), .QN(n14850) );
  DFF_X1 \REGISTERS_reg[37][0]  ( .D(n8762), .CK(CLK), .QN(n14851) );
  DFF_X1 \REGISTERS_reg[38][19]  ( .D(n8749), .CK(CLK), .Q(n578), .QN(n12921)
         );
  DFF_X1 \REGISTERS_reg[38][18]  ( .D(n8748), .CK(CLK), .Q(n580), .QN(n12920)
         );
  DFF_X1 \REGISTERS_reg[38][17]  ( .D(n8747), .CK(CLK), .Q(n582), .QN(n12919)
         );
  DFF_X1 \REGISTERS_reg[38][16]  ( .D(n8746), .CK(CLK), .Q(n584), .QN(n12918)
         );
  DFF_X1 \REGISTERS_reg[38][15]  ( .D(n8745), .CK(CLK), .Q(n586), .QN(n12917)
         );
  DFF_X1 \REGISTERS_reg[38][14]  ( .D(n8744), .CK(CLK), .Q(n588), .QN(n12916)
         );
  DFF_X1 \REGISTERS_reg[38][13]  ( .D(n8743), .CK(CLK), .Q(n590), .QN(n12915)
         );
  DFF_X1 \REGISTERS_reg[38][12]  ( .D(n8742), .CK(CLK), .Q(n592), .QN(n12914)
         );
  DFF_X1 \REGISTERS_reg[38][11]  ( .D(n8741), .CK(CLK), .Q(n594), .QN(n12913)
         );
  DFF_X1 \REGISTERS_reg[38][10]  ( .D(n8740), .CK(CLK), .Q(n596), .QN(n12912)
         );
  DFF_X1 \REGISTERS_reg[38][9]  ( .D(n8739), .CK(CLK), .Q(n598), .QN(n12911)
         );
  DFF_X1 \REGISTERS_reg[38][8]  ( .D(n8738), .CK(CLK), .Q(n600), .QN(n12910)
         );
  DFF_X1 \REGISTERS_reg[38][7]  ( .D(n8737), .CK(CLK), .Q(n602), .QN(n12909)
         );
  DFF_X1 \REGISTERS_reg[38][6]  ( .D(n8736), .CK(CLK), .Q(n604), .QN(n12908)
         );
  DFF_X1 \REGISTERS_reg[38][5]  ( .D(n8735), .CK(CLK), .Q(n606), .QN(n12907)
         );
  DFF_X1 \REGISTERS_reg[38][4]  ( .D(n8734), .CK(CLK), .Q(n608), .QN(n12906)
         );
  DFF_X1 \REGISTERS_reg[38][3]  ( .D(n8733), .CK(CLK), .Q(n610), .QN(n12905)
         );
  DFF_X1 \REGISTERS_reg[38][2]  ( .D(n8732), .CK(CLK), .Q(n612), .QN(n12904)
         );
  DFF_X1 \REGISTERS_reg[38][1]  ( .D(n8731), .CK(CLK), .Q(n614), .QN(n12903)
         );
  DFF_X1 \REGISTERS_reg[38][0]  ( .D(n8730), .CK(CLK), .Q(n616), .QN(n12902)
         );
  DFF_X1 \REGISTERS_reg[39][31]  ( .D(n8729), .CK(CLK), .Q(n98), .QN(n12709)
         );
  DFF_X1 \REGISTERS_reg[41][31]  ( .D(n8665), .CK(CLK), .Q(n6241), .QN(n12901)
         );
  DFF_X1 \REGISTERS_reg[41][30]  ( .D(n8664), .CK(CLK), .Q(n6240), .QN(n12900)
         );
  DFF_X1 \REGISTERS_reg[41][29]  ( .D(n8663), .CK(CLK), .Q(n6239), .QN(n12899)
         );
  DFF_X1 \REGISTERS_reg[41][28]  ( .D(n8662), .CK(CLK), .Q(n6238), .QN(n12898)
         );
  DFF_X1 \REGISTERS_reg[41][27]  ( .D(n8661), .CK(CLK), .Q(n6237), .QN(n12897)
         );
  DFF_X1 \REGISTERS_reg[41][26]  ( .D(n8660), .CK(CLK), .Q(n6236), .QN(n12896)
         );
  DFF_X1 \REGISTERS_reg[41][25]  ( .D(n8659), .CK(CLK), .Q(n6235), .QN(n12895)
         );
  DFF_X1 \REGISTERS_reg[41][24]  ( .D(n8658), .CK(CLK), .Q(n6234), .QN(n12894)
         );
  DFF_X1 \REGISTERS_reg[41][23]  ( .D(n8657), .CK(CLK), .Q(n6233), .QN(n12893)
         );
  DFF_X1 \REGISTERS_reg[41][22]  ( .D(n8656), .CK(CLK), .Q(n6232), .QN(n12892)
         );
  DFF_X1 \REGISTERS_reg[41][21]  ( .D(n8655), .CK(CLK), .Q(n6231), .QN(n12891)
         );
  DFF_X1 \REGISTERS_reg[41][20]  ( .D(n8654), .CK(CLK), .Q(n6230), .QN(n12890)
         );
  DFF_X1 \REGISTERS_reg[41][19]  ( .D(n8653), .CK(CLK), .Q(n6229), .QN(n12889)
         );
  DFF_X1 \REGISTERS_reg[41][18]  ( .D(n8652), .CK(CLK), .Q(n6228), .QN(n12888)
         );
  DFF_X1 \REGISTERS_reg[41][17]  ( .D(n8651), .CK(CLK), .Q(n6227), .QN(n12887)
         );
  DFF_X1 \REGISTERS_reg[41][16]  ( .D(n8650), .CK(CLK), .Q(n6226), .QN(n12886)
         );
  DFF_X1 \REGISTERS_reg[41][15]  ( .D(n8649), .CK(CLK), .Q(n6225), .QN(n12885)
         );
  DFF_X1 \REGISTERS_reg[41][14]  ( .D(n8648), .CK(CLK), .Q(n6224), .QN(n12884)
         );
  DFF_X1 \REGISTERS_reg[41][13]  ( .D(n8647), .CK(CLK), .Q(n6223), .QN(n12883)
         );
  DFF_X1 \REGISTERS_reg[41][12]  ( .D(n8646), .CK(CLK), .Q(n6222), .QN(n12882)
         );
  DFF_X1 \REGISTERS_reg[41][11]  ( .D(n8645), .CK(CLK), .Q(n6221), .QN(n12881)
         );
  DFF_X1 \REGISTERS_reg[41][10]  ( .D(n8644), .CK(CLK), .Q(n6220), .QN(n12880)
         );
  DFF_X1 \REGISTERS_reg[41][9]  ( .D(n8643), .CK(CLK), .Q(n6219), .QN(n12879)
         );
  DFF_X1 \REGISTERS_reg[41][8]  ( .D(n8642), .CK(CLK), .Q(n6218), .QN(n12878)
         );
  DFF_X1 \REGISTERS_reg[41][7]  ( .D(n8641), .CK(CLK), .Q(n6217), .QN(n12877)
         );
  DFF_X1 \REGISTERS_reg[41][6]  ( .D(n8640), .CK(CLK), .Q(n6216), .QN(n12876)
         );
  DFF_X1 \REGISTERS_reg[41][5]  ( .D(n8639), .CK(CLK), .Q(n6215), .QN(n12875)
         );
  DFF_X1 \REGISTERS_reg[41][4]  ( .D(n8638), .CK(CLK), .Q(n6214), .QN(n12874)
         );
  DFF_X1 \REGISTERS_reg[41][3]  ( .D(n8637), .CK(CLK), .Q(n6213), .QN(n12873)
         );
  DFF_X1 \REGISTERS_reg[41][2]  ( .D(n8636), .CK(CLK), .Q(n6212), .QN(n12872)
         );
  DFF_X1 \REGISTERS_reg[41][1]  ( .D(n8635), .CK(CLK), .Q(n6211), .QN(n12871)
         );
  DFF_X1 \REGISTERS_reg[41][0]  ( .D(n8634), .CK(CLK), .Q(n6210), .QN(n12870)
         );
  DFF_X1 \REGISTERS_reg[42][31]  ( .D(n8633), .CK(CLK), .QN(n14852) );
  DFF_X1 \REGISTERS_reg[42][30]  ( .D(n8632), .CK(CLK), .QN(n14853) );
  DFF_X1 \REGISTERS_reg[42][29]  ( .D(n8631), .CK(CLK), .QN(n14854) );
  DFF_X1 \REGISTERS_reg[42][28]  ( .D(n8630), .CK(CLK), .QN(n14855) );
  DFF_X1 \REGISTERS_reg[42][27]  ( .D(n8629), .CK(CLK), .QN(n14856) );
  DFF_X1 \REGISTERS_reg[42][26]  ( .D(n8628), .CK(CLK), .QN(n14857) );
  DFF_X1 \REGISTERS_reg[42][25]  ( .D(n8627), .CK(CLK), .QN(n14858) );
  DFF_X1 \REGISTERS_reg[42][24]  ( .D(n8626), .CK(CLK), .QN(n14859) );
  DFF_X1 \REGISTERS_reg[42][23]  ( .D(n8625), .CK(CLK), .QN(n14860) );
  DFF_X1 \REGISTERS_reg[42][22]  ( .D(n8624), .CK(CLK), .QN(n14861) );
  DFF_X1 \REGISTERS_reg[42][21]  ( .D(n8623), .CK(CLK), .QN(n14862) );
  DFF_X1 \REGISTERS_reg[42][20]  ( .D(n8622), .CK(CLK), .QN(n14863) );
  DFF_X1 \REGISTERS_reg[42][19]  ( .D(n8621), .CK(CLK), .QN(n14864) );
  DFF_X1 \REGISTERS_reg[42][18]  ( .D(n8620), .CK(CLK), .QN(n14865) );
  DFF_X1 \REGISTERS_reg[42][17]  ( .D(n8619), .CK(CLK), .QN(n14866) );
  DFF_X1 \REGISTERS_reg[42][16]  ( .D(n8618), .CK(CLK), .QN(n14867) );
  DFF_X1 \REGISTERS_reg[42][15]  ( .D(n8617), .CK(CLK), .QN(n14868) );
  DFF_X1 \REGISTERS_reg[42][14]  ( .D(n8616), .CK(CLK), .QN(n14869) );
  DFF_X1 \REGISTERS_reg[42][13]  ( .D(n8615), .CK(CLK), .QN(n14870) );
  DFF_X1 \REGISTERS_reg[42][12]  ( .D(n8614), .CK(CLK), .QN(n14871) );
  DFF_X1 \REGISTERS_reg[42][11]  ( .D(n8613), .CK(CLK), .QN(n14872) );
  DFF_X1 \REGISTERS_reg[42][10]  ( .D(n8612), .CK(CLK), .QN(n14873) );
  DFF_X1 \REGISTERS_reg[42][9]  ( .D(n8611), .CK(CLK), .QN(n14874) );
  DFF_X1 \REGISTERS_reg[42][8]  ( .D(n8610), .CK(CLK), .QN(n14875) );
  DFF_X1 \REGISTERS_reg[42][7]  ( .D(n8609), .CK(CLK), .QN(n14876) );
  DFF_X1 \REGISTERS_reg[42][6]  ( .D(n8608), .CK(CLK), .QN(n14877) );
  DFF_X1 \REGISTERS_reg[42][5]  ( .D(n8607), .CK(CLK), .QN(n14878) );
  DFF_X1 \REGISTERS_reg[42][4]  ( .D(n8606), .CK(CLK), .QN(n14879) );
  DFF_X1 \REGISTERS_reg[42][3]  ( .D(n8605), .CK(CLK), .QN(n14880) );
  DFF_X1 \REGISTERS_reg[42][2]  ( .D(n8604), .CK(CLK), .QN(n14881) );
  DFF_X1 \REGISTERS_reg[42][1]  ( .D(n8603), .CK(CLK), .QN(n14882) );
  DFF_X1 \REGISTERS_reg[42][0]  ( .D(n8602), .CK(CLK), .QN(n14883) );
  DFF_X1 \REGISTERS_reg[43][31]  ( .D(n8601), .CK(CLK), .QN(n14884) );
  DFF_X1 \REGISTERS_reg[43][30]  ( .D(n8600), .CK(CLK), .QN(n14885) );
  DFF_X1 \REGISTERS_reg[43][29]  ( .D(n8599), .CK(CLK), .QN(n14886) );
  DFF_X1 \REGISTERS_reg[43][28]  ( .D(n8598), .CK(CLK), .QN(n14887) );
  DFF_X1 \REGISTERS_reg[43][27]  ( .D(n8597), .CK(CLK), .QN(n14888) );
  DFF_X1 \REGISTERS_reg[43][26]  ( .D(n8596), .CK(CLK), .QN(n14889) );
  DFF_X1 \REGISTERS_reg[43][25]  ( .D(n8595), .CK(CLK), .QN(n14890) );
  DFF_X1 \REGISTERS_reg[43][24]  ( .D(n8594), .CK(CLK), .QN(n14891) );
  DFF_X1 \REGISTERS_reg[43][23]  ( .D(n8593), .CK(CLK), .QN(n14892) );
  DFF_X1 \REGISTERS_reg[43][22]  ( .D(n8592), .CK(CLK), .QN(n14893) );
  DFF_X1 \REGISTERS_reg[43][21]  ( .D(n8591), .CK(CLK), .QN(n14894) );
  DFF_X1 \REGISTERS_reg[43][20]  ( .D(n8590), .CK(CLK), .QN(n14895) );
  DFF_X1 \REGISTERS_reg[43][19]  ( .D(n8589), .CK(CLK), .QN(n14896) );
  DFF_X1 \REGISTERS_reg[43][18]  ( .D(n8588), .CK(CLK), .QN(n14897) );
  DFF_X1 \REGISTERS_reg[43][17]  ( .D(n8587), .CK(CLK), .QN(n14898) );
  DFF_X1 \REGISTERS_reg[43][16]  ( .D(n8586), .CK(CLK), .QN(n14899) );
  DFF_X1 \REGISTERS_reg[43][15]  ( .D(n8585), .CK(CLK), .QN(n14900) );
  DFF_X1 \REGISTERS_reg[43][14]  ( .D(n8584), .CK(CLK), .QN(n14901) );
  DFF_X1 \REGISTERS_reg[43][13]  ( .D(n8583), .CK(CLK), .QN(n14902) );
  DFF_X1 \REGISTERS_reg[43][12]  ( .D(n8582), .CK(CLK), .QN(n14903) );
  DFF_X1 \REGISTERS_reg[43][11]  ( .D(n8581), .CK(CLK), .QN(n14904) );
  DFF_X1 \REGISTERS_reg[43][10]  ( .D(n8580), .CK(CLK), .QN(n14905) );
  DFF_X1 \REGISTERS_reg[43][9]  ( .D(n8579), .CK(CLK), .QN(n14906) );
  DFF_X1 \REGISTERS_reg[43][8]  ( .D(n8578), .CK(CLK), .QN(n14907) );
  DFF_X1 \REGISTERS_reg[43][7]  ( .D(n8577), .CK(CLK), .QN(n14908) );
  DFF_X1 \REGISTERS_reg[43][6]  ( .D(n8576), .CK(CLK), .QN(n14909) );
  DFF_X1 \REGISTERS_reg[43][5]  ( .D(n8575), .CK(CLK), .QN(n14910) );
  DFF_X1 \REGISTERS_reg[43][4]  ( .D(n8574), .CK(CLK), .QN(n14911) );
  DFF_X1 \REGISTERS_reg[43][3]  ( .D(n8573), .CK(CLK), .QN(n14912) );
  DFF_X1 \REGISTERS_reg[43][2]  ( .D(n8572), .CK(CLK), .QN(n14913) );
  DFF_X1 \REGISTERS_reg[43][1]  ( .D(n8571), .CK(CLK), .QN(n14914) );
  DFF_X1 \REGISTERS_reg[43][0]  ( .D(n8570), .CK(CLK), .QN(n14915) );
  DFF_X1 \REGISTERS_reg[44][31]  ( .D(n8569), .CK(CLK), .QN(n14916) );
  DFF_X1 \REGISTERS_reg[44][30]  ( .D(n8568), .CK(CLK), .QN(n14917) );
  DFF_X1 \REGISTERS_reg[44][29]  ( .D(n8567), .CK(CLK), .QN(n14918) );
  DFF_X1 \REGISTERS_reg[44][28]  ( .D(n8566), .CK(CLK), .QN(n14919) );
  DFF_X1 \REGISTERS_reg[44][27]  ( .D(n8565), .CK(CLK), .QN(n14920) );
  DFF_X1 \REGISTERS_reg[44][26]  ( .D(n8564), .CK(CLK), .QN(n14921) );
  DFF_X1 \REGISTERS_reg[44][25]  ( .D(n8563), .CK(CLK), .QN(n14922) );
  DFF_X1 \REGISTERS_reg[44][24]  ( .D(n8562), .CK(CLK), .QN(n14923) );
  DFF_X1 \REGISTERS_reg[44][23]  ( .D(n8561), .CK(CLK), .QN(n14924) );
  DFF_X1 \REGISTERS_reg[44][22]  ( .D(n8560), .CK(CLK), .QN(n14925) );
  DFF_X1 \REGISTERS_reg[44][21]  ( .D(n8559), .CK(CLK), .QN(n14926) );
  DFF_X1 \REGISTERS_reg[44][20]  ( .D(n8558), .CK(CLK), .QN(n14927) );
  DFF_X1 \REGISTERS_reg[44][19]  ( .D(n8557), .CK(CLK), .QN(n14928) );
  DFF_X1 \REGISTERS_reg[44][18]  ( .D(n8556), .CK(CLK), .QN(n14929) );
  DFF_X1 \REGISTERS_reg[44][17]  ( .D(n8555), .CK(CLK), .QN(n14930) );
  DFF_X1 \REGISTERS_reg[44][16]  ( .D(n8554), .CK(CLK), .QN(n14931) );
  DFF_X1 \REGISTERS_reg[44][15]  ( .D(n8553), .CK(CLK), .QN(n14932) );
  DFF_X1 \REGISTERS_reg[44][14]  ( .D(n8552), .CK(CLK), .QN(n14933) );
  DFF_X1 \REGISTERS_reg[44][13]  ( .D(n8551), .CK(CLK), .QN(n14934) );
  DFF_X1 \REGISTERS_reg[44][12]  ( .D(n8550), .CK(CLK), .QN(n14935) );
  DFF_X1 \REGISTERS_reg[44][11]  ( .D(n8549), .CK(CLK), .QN(n14936) );
  DFF_X1 \REGISTERS_reg[44][10]  ( .D(n8548), .CK(CLK), .QN(n14937) );
  DFF_X1 \REGISTERS_reg[44][9]  ( .D(n8547), .CK(CLK), .QN(n14938) );
  DFF_X1 \REGISTERS_reg[44][8]  ( .D(n8546), .CK(CLK), .QN(n14939) );
  DFF_X1 \REGISTERS_reg[44][7]  ( .D(n8545), .CK(CLK), .QN(n14940) );
  DFF_X1 \REGISTERS_reg[44][6]  ( .D(n8544), .CK(CLK), .QN(n14941) );
  DFF_X1 \REGISTERS_reg[44][5]  ( .D(n8543), .CK(CLK), .QN(n14942) );
  DFF_X1 \REGISTERS_reg[44][4]  ( .D(n8542), .CK(CLK), .QN(n14943) );
  DFF_X1 \REGISTERS_reg[44][3]  ( .D(n8541), .CK(CLK), .QN(n14944) );
  DFF_X1 \REGISTERS_reg[44][2]  ( .D(n8540), .CK(CLK), .QN(n14945) );
  DFF_X1 \REGISTERS_reg[44][1]  ( .D(n8539), .CK(CLK), .QN(n14946) );
  DFF_X1 \REGISTERS_reg[44][0]  ( .D(n8538), .CK(CLK), .QN(n14947) );
  DFF_X1 \REGISTERS_reg[46][31]  ( .D(n8505), .CK(CLK), .Q(n6177), .QN(n12869)
         );
  DFF_X1 \REGISTERS_reg[46][30]  ( .D(n8504), .CK(CLK), .Q(n6176), .QN(n12868)
         );
  DFF_X1 \REGISTERS_reg[46][29]  ( .D(n8503), .CK(CLK), .Q(n6175), .QN(n12867)
         );
  DFF_X1 \REGISTERS_reg[46][28]  ( .D(n8502), .CK(CLK), .Q(n6174), .QN(n12866)
         );
  DFF_X1 \REGISTERS_reg[46][27]  ( .D(n8501), .CK(CLK), .Q(n6173), .QN(n12865)
         );
  DFF_X1 \REGISTERS_reg[46][26]  ( .D(n8500), .CK(CLK), .Q(n6172), .QN(n12864)
         );
  DFF_X1 \REGISTERS_reg[46][25]  ( .D(n8499), .CK(CLK), .Q(n6171), .QN(n12863)
         );
  DFF_X1 \REGISTERS_reg[46][24]  ( .D(n8498), .CK(CLK), .Q(n6170), .QN(n12862)
         );
  DFF_X1 \REGISTERS_reg[46][23]  ( .D(n8497), .CK(CLK), .Q(n6169), .QN(n12861)
         );
  DFF_X1 \REGISTERS_reg[46][22]  ( .D(n8496), .CK(CLK), .Q(n6168), .QN(n12860)
         );
  DFF_X1 \REGISTERS_reg[46][21]  ( .D(n8495), .CK(CLK), .Q(n6167), .QN(n12859)
         );
  DFF_X1 \REGISTERS_reg[46][20]  ( .D(n8494), .CK(CLK), .Q(n6166), .QN(n12858)
         );
  DFF_X1 \REGISTERS_reg[46][19]  ( .D(n8493), .CK(CLK), .Q(n6165), .QN(n12857)
         );
  DFF_X1 \REGISTERS_reg[46][18]  ( .D(n8492), .CK(CLK), .Q(n6164), .QN(n12856)
         );
  DFF_X1 \REGISTERS_reg[46][17]  ( .D(n8491), .CK(CLK), .Q(n6163), .QN(n12855)
         );
  DFF_X1 \REGISTERS_reg[46][16]  ( .D(n8490), .CK(CLK), .Q(n6162), .QN(n12854)
         );
  DFF_X1 \REGISTERS_reg[46][15]  ( .D(n8489), .CK(CLK), .Q(n6161), .QN(n12853)
         );
  DFF_X1 \REGISTERS_reg[46][14]  ( .D(n8488), .CK(CLK), .Q(n6160), .QN(n12852)
         );
  DFF_X1 \REGISTERS_reg[46][13]  ( .D(n8487), .CK(CLK), .Q(n6159), .QN(n12851)
         );
  DFF_X1 \REGISTERS_reg[46][12]  ( .D(n8486), .CK(CLK), .Q(n6158), .QN(n12850)
         );
  DFF_X1 \REGISTERS_reg[46][11]  ( .D(n8485), .CK(CLK), .Q(n6157), .QN(n12849)
         );
  DFF_X1 \REGISTERS_reg[46][10]  ( .D(n8484), .CK(CLK), .Q(n6156), .QN(n12848)
         );
  DFF_X1 \REGISTERS_reg[46][9]  ( .D(n8483), .CK(CLK), .Q(n6155), .QN(n12847)
         );
  DFF_X1 \REGISTERS_reg[46][8]  ( .D(n8482), .CK(CLK), .Q(n6154), .QN(n12846)
         );
  DFF_X1 \REGISTERS_reg[46][7]  ( .D(n8481), .CK(CLK), .Q(n6153), .QN(n12845)
         );
  DFF_X1 \REGISTERS_reg[46][6]  ( .D(n8480), .CK(CLK), .Q(n6152), .QN(n12844)
         );
  DFF_X1 \REGISTERS_reg[46][5]  ( .D(n8479), .CK(CLK), .Q(n6151), .QN(n12843)
         );
  DFF_X1 \REGISTERS_reg[46][4]  ( .D(n8478), .CK(CLK), .Q(n6150), .QN(n12842)
         );
  DFF_X1 \REGISTERS_reg[46][3]  ( .D(n8477), .CK(CLK), .Q(n6149), .QN(n12841)
         );
  DFF_X1 \REGISTERS_reg[46][2]  ( .D(n8476), .CK(CLK), .Q(n6148), .QN(n12840)
         );
  DFF_X1 \REGISTERS_reg[46][1]  ( .D(n8475), .CK(CLK), .Q(n6147), .QN(n12839)
         );
  DFF_X1 \REGISTERS_reg[46][0]  ( .D(n8474), .CK(CLK), .Q(n6146), .QN(n12838)
         );
  DFF_X1 \REGISTERS_reg[47][31]  ( .D(n8473), .CK(CLK), .QN(n14949) );
  DFF_X1 \REGISTERS_reg[47][30]  ( .D(n8472), .CK(CLK), .QN(n14950) );
  DFF_X1 \REGISTERS_reg[47][29]  ( .D(n8471), .CK(CLK), .QN(n14951) );
  DFF_X1 \REGISTERS_reg[47][28]  ( .D(n8470), .CK(CLK), .QN(n14952) );
  DFF_X1 \REGISTERS_reg[47][27]  ( .D(n8469), .CK(CLK), .QN(n14953) );
  DFF_X1 \REGISTERS_reg[47][26]  ( .D(n8468), .CK(CLK), .QN(n14954) );
  DFF_X1 \REGISTERS_reg[47][25]  ( .D(n8467), .CK(CLK), .QN(n14955) );
  DFF_X1 \REGISTERS_reg[47][24]  ( .D(n8466), .CK(CLK), .QN(n14956) );
  DFF_X1 \REGISTERS_reg[47][23]  ( .D(n8465), .CK(CLK), .QN(n14957) );
  DFF_X1 \REGISTERS_reg[47][22]  ( .D(n8464), .CK(CLK), .QN(n14958) );
  DFF_X1 \REGISTERS_reg[47][21]  ( .D(n8463), .CK(CLK), .QN(n14959) );
  DFF_X1 \REGISTERS_reg[47][20]  ( .D(n8462), .CK(CLK), .QN(n14960) );
  DFF_X1 \REGISTERS_reg[47][19]  ( .D(n8461), .CK(CLK), .QN(n14961) );
  DFF_X1 \REGISTERS_reg[47][18]  ( .D(n8460), .CK(CLK), .QN(n14962) );
  DFF_X1 \REGISTERS_reg[47][17]  ( .D(n8459), .CK(CLK), .QN(n14963) );
  DFF_X1 \REGISTERS_reg[47][16]  ( .D(n8458), .CK(CLK), .QN(n14964) );
  DFF_X1 \REGISTERS_reg[47][15]  ( .D(n8457), .CK(CLK), .QN(n14965) );
  DFF_X1 \REGISTERS_reg[47][14]  ( .D(n8456), .CK(CLK), .QN(n14966) );
  DFF_X1 \REGISTERS_reg[47][13]  ( .D(n8455), .CK(CLK), .QN(n14967) );
  DFF_X1 \REGISTERS_reg[47][12]  ( .D(n8454), .CK(CLK), .QN(n14968) );
  DFF_X1 \REGISTERS_reg[47][11]  ( .D(n8453), .CK(CLK), .QN(n14969) );
  DFF_X1 \REGISTERS_reg[47][10]  ( .D(n8452), .CK(CLK), .QN(n14970) );
  DFF_X1 \REGISTERS_reg[47][9]  ( .D(n8451), .CK(CLK), .QN(n14971) );
  DFF_X1 \REGISTERS_reg[47][8]  ( .D(n8450), .CK(CLK), .QN(n14972) );
  DFF_X1 \REGISTERS_reg[47][7]  ( .D(n8449), .CK(CLK), .QN(n14973) );
  DFF_X1 \REGISTERS_reg[47][6]  ( .D(n8448), .CK(CLK), .QN(n14974) );
  DFF_X1 \REGISTERS_reg[47][5]  ( .D(n8447), .CK(CLK), .QN(n14975) );
  DFF_X1 \REGISTERS_reg[47][4]  ( .D(n8446), .CK(CLK), .QN(n14976) );
  DFF_X1 \REGISTERS_reg[47][3]  ( .D(n8445), .CK(CLK), .QN(n14977) );
  DFF_X1 \REGISTERS_reg[47][2]  ( .D(n8444), .CK(CLK), .QN(n14978) );
  DFF_X1 \REGISTERS_reg[47][1]  ( .D(n8443), .CK(CLK), .QN(n14979) );
  DFF_X1 \REGISTERS_reg[47][0]  ( .D(n8442), .CK(CLK), .QN(n14980) );
  DFF_X1 \REGISTERS_reg[51][31]  ( .D(n8345), .CK(CLK), .QN(n15014) );
  DFF_X1 \REGISTERS_reg[51][30]  ( .D(n8344), .CK(CLK), .QN(n15015) );
  DFF_X1 \REGISTERS_reg[51][29]  ( .D(n8343), .CK(CLK), .QN(n15016) );
  DFF_X1 \REGISTERS_reg[51][28]  ( .D(n8342), .CK(CLK), .QN(n15017) );
  DFF_X1 \REGISTERS_reg[51][27]  ( .D(n8341), .CK(CLK), .QN(n15018) );
  DFF_X1 \REGISTERS_reg[51][26]  ( .D(n8340), .CK(CLK), .QN(n15019) );
  DFF_X1 \REGISTERS_reg[51][25]  ( .D(n8339), .CK(CLK), .QN(n15020) );
  DFF_X1 \REGISTERS_reg[51][24]  ( .D(n8338), .CK(CLK), .QN(n15021) );
  DFF_X1 \REGISTERS_reg[51][23]  ( .D(n8337), .CK(CLK), .QN(n15022) );
  DFF_X1 \REGISTERS_reg[51][22]  ( .D(n8336), .CK(CLK), .QN(n15023) );
  DFF_X1 \REGISTERS_reg[51][21]  ( .D(n8335), .CK(CLK), .QN(n15024) );
  DFF_X1 \REGISTERS_reg[51][20]  ( .D(n8334), .CK(CLK), .QN(n15025) );
  DFF_X1 \REGISTERS_reg[51][19]  ( .D(n8333), .CK(CLK), .QN(n15026) );
  DFF_X1 \REGISTERS_reg[51][18]  ( .D(n8332), .CK(CLK), .QN(n15027) );
  DFF_X1 \REGISTERS_reg[51][17]  ( .D(n8331), .CK(CLK), .QN(n15028) );
  DFF_X1 \REGISTERS_reg[51][16]  ( .D(n8330), .CK(CLK), .QN(n15029) );
  DFF_X1 \REGISTERS_reg[51][15]  ( .D(n8329), .CK(CLK), .QN(n15030) );
  DFF_X1 \REGISTERS_reg[51][14]  ( .D(n8328), .CK(CLK), .QN(n15031) );
  DFF_X1 \REGISTERS_reg[51][13]  ( .D(n8327), .CK(CLK), .QN(n15032) );
  DFF_X1 \REGISTERS_reg[51][12]  ( .D(n8326), .CK(CLK), .QN(n15033) );
  DFF_X1 \REGISTERS_reg[51][11]  ( .D(n8325), .CK(CLK), .QN(n15034) );
  DFF_X1 \REGISTERS_reg[51][10]  ( .D(n8324), .CK(CLK), .QN(n15035) );
  DFF_X1 \REGISTERS_reg[51][9]  ( .D(n8323), .CK(CLK), .QN(n15036) );
  DFF_X1 \REGISTERS_reg[51][8]  ( .D(n8322), .CK(CLK), .QN(n15037) );
  DFF_X1 \REGISTERS_reg[51][7]  ( .D(n8321), .CK(CLK), .QN(n15038) );
  DFF_X1 \REGISTERS_reg[51][6]  ( .D(n8320), .CK(CLK), .QN(n15039) );
  DFF_X1 \REGISTERS_reg[51][5]  ( .D(n8319), .CK(CLK), .QN(n15040) );
  DFF_X1 \REGISTERS_reg[51][4]  ( .D(n8318), .CK(CLK), .QN(n15041) );
  DFF_X1 \REGISTERS_reg[51][3]  ( .D(n8317), .CK(CLK), .QN(n15042) );
  DFF_X1 \REGISTERS_reg[51][2]  ( .D(n8316), .CK(CLK), .QN(n15043) );
  DFF_X1 \REGISTERS_reg[51][1]  ( .D(n8315), .CK(CLK), .QN(n15044) );
  DFF_X1 \REGISTERS_reg[51][0]  ( .D(n8314), .CK(CLK), .QN(n15045) );
  DFF_X1 \REGISTERS_reg[52][31]  ( .D(n8313), .CK(CLK), .QN(n15046) );
  DFF_X1 \REGISTERS_reg[52][30]  ( .D(n8312), .CK(CLK), .QN(n15047) );
  DFF_X1 \REGISTERS_reg[52][29]  ( .D(n8311), .CK(CLK), .QN(n15048) );
  DFF_X1 \REGISTERS_reg[52][28]  ( .D(n8310), .CK(CLK), .QN(n15049) );
  DFF_X1 \REGISTERS_reg[52][27]  ( .D(n8309), .CK(CLK), .QN(n15050) );
  DFF_X1 \REGISTERS_reg[52][26]  ( .D(n8308), .CK(CLK), .QN(n15051) );
  DFF_X1 \REGISTERS_reg[52][25]  ( .D(n8307), .CK(CLK), .QN(n15052) );
  DFF_X1 \REGISTERS_reg[52][24]  ( .D(n8306), .CK(CLK), .QN(n15053) );
  DFF_X1 \REGISTERS_reg[52][23]  ( .D(n8305), .CK(CLK), .QN(n15054) );
  DFF_X1 \REGISTERS_reg[52][22]  ( .D(n8304), .CK(CLK), .QN(n15055) );
  DFF_X1 \REGISTERS_reg[52][21]  ( .D(n8303), .CK(CLK), .QN(n15056) );
  DFF_X1 \REGISTERS_reg[52][20]  ( .D(n8302), .CK(CLK), .QN(n15057) );
  DFF_X1 \REGISTERS_reg[52][19]  ( .D(n8301), .CK(CLK), .QN(n15058) );
  DFF_X1 \REGISTERS_reg[52][18]  ( .D(n8300), .CK(CLK), .QN(n15059) );
  DFF_X1 \REGISTERS_reg[52][17]  ( .D(n8299), .CK(CLK), .QN(n15060) );
  DFF_X1 \REGISTERS_reg[52][16]  ( .D(n8298), .CK(CLK), .QN(n15061) );
  DFF_X1 \REGISTERS_reg[52][15]  ( .D(n8297), .CK(CLK), .QN(n15062) );
  DFF_X1 \REGISTERS_reg[52][14]  ( .D(n8296), .CK(CLK), .QN(n15063) );
  DFF_X1 \REGISTERS_reg[52][13]  ( .D(n8295), .CK(CLK), .QN(n15064) );
  DFF_X1 \REGISTERS_reg[52][12]  ( .D(n8294), .CK(CLK), .QN(n15065) );
  DFF_X1 \REGISTERS_reg[52][11]  ( .D(n8293), .CK(CLK), .QN(n15066) );
  DFF_X1 \REGISTERS_reg[52][10]  ( .D(n8292), .CK(CLK), .QN(n15067) );
  DFF_X1 \REGISTERS_reg[52][9]  ( .D(n8291), .CK(CLK), .QN(n15068) );
  DFF_X1 \REGISTERS_reg[52][8]  ( .D(n8290), .CK(CLK), .QN(n15069) );
  DFF_X1 \REGISTERS_reg[52][7]  ( .D(n8289), .CK(CLK), .QN(n15070) );
  DFF_X1 \REGISTERS_reg[52][6]  ( .D(n8288), .CK(CLK), .QN(n15071) );
  DFF_X1 \REGISTERS_reg[52][5]  ( .D(n8287), .CK(CLK), .QN(n15072) );
  DFF_X1 \REGISTERS_reg[52][4]  ( .D(n8286), .CK(CLK), .QN(n15073) );
  DFF_X1 \REGISTERS_reg[52][3]  ( .D(n8285), .CK(CLK), .QN(n15074) );
  DFF_X1 \REGISTERS_reg[52][2]  ( .D(n8284), .CK(CLK), .QN(n15075) );
  DFF_X1 \REGISTERS_reg[52][1]  ( .D(n8283), .CK(CLK), .QN(n15076) );
  DFF_X1 \REGISTERS_reg[52][0]  ( .D(n8282), .CK(CLK), .QN(n15077) );
  DFF_X1 \REGISTERS_reg[53][31]  ( .D(n8281), .CK(CLK), .QN(n15078) );
  DFF_X1 \REGISTERS_reg[53][30]  ( .D(n8280), .CK(CLK), .QN(n15079) );
  DFF_X1 \REGISTERS_reg[53][29]  ( .D(n8279), .CK(CLK), .QN(n15080) );
  DFF_X1 \REGISTERS_reg[53][28]  ( .D(n8278), .CK(CLK), .QN(n15081) );
  DFF_X1 \REGISTERS_reg[53][27]  ( .D(n8277), .CK(CLK), .QN(n15082) );
  DFF_X1 \REGISTERS_reg[53][26]  ( .D(n8276), .CK(CLK), .QN(n15083) );
  DFF_X1 \REGISTERS_reg[53][25]  ( .D(n8275), .CK(CLK), .QN(n15084) );
  DFF_X1 \REGISTERS_reg[53][24]  ( .D(n8274), .CK(CLK), .QN(n15085) );
  DFF_X1 \REGISTERS_reg[53][23]  ( .D(n8273), .CK(CLK), .QN(n15086) );
  DFF_X1 \REGISTERS_reg[53][22]  ( .D(n8272), .CK(CLK), .QN(n15087) );
  DFF_X1 \REGISTERS_reg[53][21]  ( .D(n8271), .CK(CLK), .QN(n15088) );
  DFF_X1 \REGISTERS_reg[53][20]  ( .D(n8270), .CK(CLK), .QN(n15089) );
  DFF_X1 \REGISTERS_reg[53][19]  ( .D(n8269), .CK(CLK), .QN(n15090) );
  DFF_X1 \REGISTERS_reg[53][18]  ( .D(n8268), .CK(CLK), .QN(n15091) );
  DFF_X1 \REGISTERS_reg[53][17]  ( .D(n8267), .CK(CLK), .QN(n15092) );
  DFF_X1 \REGISTERS_reg[53][16]  ( .D(n8266), .CK(CLK), .QN(n15093) );
  DFF_X1 \REGISTERS_reg[53][15]  ( .D(n8265), .CK(CLK), .QN(n15094) );
  DFF_X1 \REGISTERS_reg[53][14]  ( .D(n8264), .CK(CLK), .QN(n15095) );
  DFF_X1 \REGISTERS_reg[53][13]  ( .D(n8263), .CK(CLK), .QN(n15096) );
  DFF_X1 \REGISTERS_reg[53][12]  ( .D(n8262), .CK(CLK), .QN(n15097) );
  DFF_X1 \REGISTERS_reg[53][11]  ( .D(n8261), .CK(CLK), .QN(n15098) );
  DFF_X1 \REGISTERS_reg[53][10]  ( .D(n8260), .CK(CLK), .QN(n15099) );
  DFF_X1 \REGISTERS_reg[53][9]  ( .D(n8259), .CK(CLK), .QN(n15100) );
  DFF_X1 \REGISTERS_reg[53][8]  ( .D(n8258), .CK(CLK), .QN(n15101) );
  DFF_X1 \REGISTERS_reg[53][7]  ( .D(n8257), .CK(CLK), .QN(n15102) );
  DFF_X1 \REGISTERS_reg[53][6]  ( .D(n8256), .CK(CLK), .QN(n15103) );
  DFF_X1 \REGISTERS_reg[53][5]  ( .D(n8255), .CK(CLK), .QN(n15104) );
  DFF_X1 \REGISTERS_reg[53][4]  ( .D(n8254), .CK(CLK), .QN(n15105) );
  DFF_X1 \REGISTERS_reg[53][3]  ( .D(n8253), .CK(CLK), .QN(n15106) );
  DFF_X1 \REGISTERS_reg[53][2]  ( .D(n8252), .CK(CLK), .QN(n15107) );
  DFF_X1 \REGISTERS_reg[53][1]  ( .D(n8251), .CK(CLK), .QN(n15108) );
  DFF_X1 \REGISTERS_reg[53][0]  ( .D(n8250), .CK(CLK), .QN(n15109) );
  DFF_X1 \REGISTERS_reg[54][31]  ( .D(n8249), .CK(CLK), .QN(n15110) );
  DFF_X1 \REGISTERS_reg[54][30]  ( .D(n8248), .CK(CLK), .QN(n15111) );
  DFF_X1 \REGISTERS_reg[54][29]  ( .D(n8247), .CK(CLK), .QN(n15112) );
  DFF_X1 \REGISTERS_reg[54][28]  ( .D(n8246), .CK(CLK), .QN(n15113) );
  DFF_X1 \REGISTERS_reg[54][27]  ( .D(n8245), .CK(CLK), .QN(n15114) );
  DFF_X1 \REGISTERS_reg[54][26]  ( .D(n8244), .CK(CLK), .QN(n15115) );
  DFF_X1 \REGISTERS_reg[54][25]  ( .D(n8243), .CK(CLK), .QN(n15116) );
  DFF_X1 \REGISTERS_reg[54][24]  ( .D(n8242), .CK(CLK), .QN(n15117) );
  DFF_X1 \REGISTERS_reg[54][23]  ( .D(n8241), .CK(CLK), .QN(n15118) );
  DFF_X1 \REGISTERS_reg[54][22]  ( .D(n8240), .CK(CLK), .QN(n15119) );
  DFF_X1 \REGISTERS_reg[54][21]  ( .D(n8239), .CK(CLK), .QN(n15120) );
  DFF_X1 \REGISTERS_reg[54][20]  ( .D(n8238), .CK(CLK), .QN(n15121) );
  DFF_X1 \REGISTERS_reg[54][19]  ( .D(n8237), .CK(CLK), .QN(n15122) );
  DFF_X1 \REGISTERS_reg[54][18]  ( .D(n8236), .CK(CLK), .QN(n15123) );
  DFF_X1 \REGISTERS_reg[54][17]  ( .D(n8235), .CK(CLK), .QN(n15124) );
  DFF_X1 \REGISTERS_reg[54][16]  ( .D(n8234), .CK(CLK), .QN(n15125) );
  DFF_X1 \REGISTERS_reg[54][15]  ( .D(n8233), .CK(CLK), .QN(n15126) );
  DFF_X1 \REGISTERS_reg[54][14]  ( .D(n8232), .CK(CLK), .QN(n15127) );
  DFF_X1 \REGISTERS_reg[54][13]  ( .D(n8231), .CK(CLK), .QN(n15128) );
  DFF_X1 \REGISTERS_reg[54][12]  ( .D(n8230), .CK(CLK), .QN(n15129) );
  DFF_X1 \REGISTERS_reg[54][11]  ( .D(n8229), .CK(CLK), .QN(n15130) );
  DFF_X1 \REGISTERS_reg[54][10]  ( .D(n8228), .CK(CLK), .QN(n15131) );
  DFF_X1 \REGISTERS_reg[54][9]  ( .D(n8227), .CK(CLK), .QN(n15132) );
  DFF_X1 \REGISTERS_reg[54][8]  ( .D(n8226), .CK(CLK), .QN(n15133) );
  DFF_X1 \REGISTERS_reg[54][7]  ( .D(n8225), .CK(CLK), .QN(n15134) );
  DFF_X1 \REGISTERS_reg[54][6]  ( .D(n8224), .CK(CLK), .QN(n15135) );
  DFF_X1 \REGISTERS_reg[54][5]  ( .D(n8223), .CK(CLK), .QN(n15136) );
  DFF_X1 \REGISTERS_reg[54][4]  ( .D(n8222), .CK(CLK), .QN(n15137) );
  DFF_X1 \REGISTERS_reg[54][3]  ( .D(n8221), .CK(CLK), .QN(n15138) );
  DFF_X1 \REGISTERS_reg[54][2]  ( .D(n8220), .CK(CLK), .QN(n15139) );
  DFF_X1 \REGISTERS_reg[54][1]  ( .D(n8219), .CK(CLK), .QN(n15140) );
  DFF_X1 \REGISTERS_reg[54][0]  ( .D(n8218), .CK(CLK), .QN(n15141) );
  DFF_X1 \REGISTERS_reg[55][31]  ( .D(n8217), .CK(CLK), .QN(n15142) );
  DFF_X1 \REGISTERS_reg[55][30]  ( .D(n8216), .CK(CLK), .QN(n15143) );
  DFF_X1 \REGISTERS_reg[55][29]  ( .D(n8215), .CK(CLK), .QN(n15144) );
  DFF_X1 \REGISTERS_reg[55][28]  ( .D(n8214), .CK(CLK), .QN(n15145) );
  DFF_X1 \REGISTERS_reg[55][27]  ( .D(n8213), .CK(CLK), .QN(n15146) );
  DFF_X1 \REGISTERS_reg[55][26]  ( .D(n8212), .CK(CLK), .QN(n15147) );
  DFF_X1 \REGISTERS_reg[55][25]  ( .D(n8211), .CK(CLK), .QN(n15148) );
  DFF_X1 \REGISTERS_reg[55][24]  ( .D(n8210), .CK(CLK), .QN(n15149) );
  DFF_X1 \REGISTERS_reg[55][23]  ( .D(n8209), .CK(CLK), .QN(n15150) );
  DFF_X1 \REGISTERS_reg[55][22]  ( .D(n8208), .CK(CLK), .QN(n15151) );
  DFF_X1 \REGISTERS_reg[55][21]  ( .D(n8207), .CK(CLK), .QN(n15152) );
  DFF_X1 \REGISTERS_reg[55][20]  ( .D(n8206), .CK(CLK), .QN(n15153) );
  DFF_X1 \REGISTERS_reg[55][19]  ( .D(n8205), .CK(CLK), .QN(n15154) );
  DFF_X1 \REGISTERS_reg[55][18]  ( .D(n8204), .CK(CLK), .QN(n15155) );
  DFF_X1 \REGISTERS_reg[55][17]  ( .D(n8203), .CK(CLK), .QN(n15156) );
  DFF_X1 \REGISTERS_reg[55][16]  ( .D(n8202), .CK(CLK), .QN(n15157) );
  DFF_X1 \REGISTERS_reg[55][15]  ( .D(n8201), .CK(CLK), .QN(n15158) );
  DFF_X1 \REGISTERS_reg[55][14]  ( .D(n8200), .CK(CLK), .QN(n15159) );
  DFF_X1 \REGISTERS_reg[55][13]  ( .D(n8199), .CK(CLK), .QN(n15160) );
  DFF_X1 \REGISTERS_reg[55][12]  ( .D(n8198), .CK(CLK), .QN(n15161) );
  DFF_X1 \REGISTERS_reg[55][11]  ( .D(n8197), .CK(CLK), .QN(n15162) );
  DFF_X1 \REGISTERS_reg[55][10]  ( .D(n8196), .CK(CLK), .QN(n15163) );
  DFF_X1 \REGISTERS_reg[55][9]  ( .D(n8195), .CK(CLK), .QN(n15164) );
  DFF_X1 \REGISTERS_reg[55][8]  ( .D(n8194), .CK(CLK), .QN(n15165) );
  DFF_X1 \REGISTERS_reg[55][7]  ( .D(n8193), .CK(CLK), .QN(n15166) );
  DFF_X1 \REGISTERS_reg[55][6]  ( .D(n8192), .CK(CLK), .QN(n15167) );
  DFF_X1 \REGISTERS_reg[55][5]  ( .D(n8191), .CK(CLK), .QN(n15168) );
  DFF_X1 \REGISTERS_reg[55][4]  ( .D(n8190), .CK(CLK), .QN(n15169) );
  DFF_X1 \REGISTERS_reg[55][3]  ( .D(n8189), .CK(CLK), .QN(n15170) );
  DFF_X1 \REGISTERS_reg[55][2]  ( .D(n8188), .CK(CLK), .QN(n15171) );
  DFF_X1 \REGISTERS_reg[55][1]  ( .D(n8187), .CK(CLK), .QN(n15172) );
  DFF_X1 \REGISTERS_reg[55][0]  ( .D(n8186), .CK(CLK), .QN(n15173) );
  DFF_X1 \REGISTERS_reg[56][31]  ( .D(n8185), .CK(CLK), .Q(n6081), .QN(n12725)
         );
  DFF_X1 \REGISTERS_reg[56][30]  ( .D(n8184), .CK(CLK), .Q(n6080), .QN(n12724)
         );
  DFF_X1 \REGISTERS_reg[56][29]  ( .D(n8183), .CK(CLK), .Q(n6079), .QN(n12723)
         );
  DFF_X1 \REGISTERS_reg[56][28]  ( .D(n8182), .CK(CLK), .Q(n6078), .QN(n12722)
         );
  DFF_X1 \REGISTERS_reg[56][27]  ( .D(n8181), .CK(CLK), .Q(n6077), .QN(n12721)
         );
  DFF_X1 \REGISTERS_reg[56][26]  ( .D(n8180), .CK(CLK), .Q(n6076), .QN(n12720)
         );
  DFF_X1 \REGISTERS_reg[56][25]  ( .D(n8179), .CK(CLK), .Q(n6075), .QN(n12719)
         );
  DFF_X1 \REGISTERS_reg[56][24]  ( .D(n8178), .CK(CLK), .Q(n6074), .QN(n12718)
         );
  DFF_X1 \REGISTERS_reg[56][23]  ( .D(n8177), .CK(CLK), .Q(n6073), .QN(n12773)
         );
  DFF_X1 \REGISTERS_reg[56][22]  ( .D(n8176), .CK(CLK), .Q(n6072), .QN(n12772)
         );
  DFF_X1 \REGISTERS_reg[56][21]  ( .D(n8175), .CK(CLK), .Q(n6071), .QN(n12771)
         );
  DFF_X1 \REGISTERS_reg[56][20]  ( .D(n8174), .CK(CLK), .Q(n6070), .QN(n12770)
         );
  DFF_X1 \REGISTERS_reg[56][19]  ( .D(n8173), .CK(CLK), .Q(n6069), .QN(n12769)
         );
  DFF_X1 \REGISTERS_reg[56][18]  ( .D(n8172), .CK(CLK), .Q(n6068), .QN(n12768)
         );
  DFF_X1 \REGISTERS_reg[56][17]  ( .D(n8171), .CK(CLK), .Q(n6067), .QN(n12767)
         );
  DFF_X1 \REGISTERS_reg[56][16]  ( .D(n8170), .CK(CLK), .Q(n6066), .QN(n12766)
         );
  DFF_X1 \REGISTERS_reg[56][15]  ( .D(n8169), .CK(CLK), .Q(n6065), .QN(n12765)
         );
  DFF_X1 \REGISTERS_reg[56][14]  ( .D(n8168), .CK(CLK), .Q(n6064), .QN(n12764)
         );
  DFF_X1 \REGISTERS_reg[56][13]  ( .D(n8167), .CK(CLK), .Q(n6063), .QN(n12763)
         );
  DFF_X1 \REGISTERS_reg[56][12]  ( .D(n8166), .CK(CLK), .Q(n6062), .QN(n12762)
         );
  DFF_X1 \REGISTERS_reg[56][11]  ( .D(n8165), .CK(CLK), .Q(n6061), .QN(n12761)
         );
  DFF_X1 \REGISTERS_reg[56][10]  ( .D(n8164), .CK(CLK), .Q(n6060), .QN(n12760)
         );
  DFF_X1 \REGISTERS_reg[56][9]  ( .D(n8163), .CK(CLK), .Q(n6059), .QN(n12759)
         );
  DFF_X1 \REGISTERS_reg[56][8]  ( .D(n8162), .CK(CLK), .Q(n6058), .QN(n12758)
         );
  DFF_X1 \REGISTERS_reg[56][7]  ( .D(n8161), .CK(CLK), .Q(n6057), .QN(n12757)
         );
  DFF_X1 \REGISTERS_reg[56][6]  ( .D(n8160), .CK(CLK), .Q(n6056), .QN(n12756)
         );
  DFF_X1 \REGISTERS_reg[56][5]  ( .D(n8159), .CK(CLK), .Q(n6055), .QN(n12755)
         );
  DFF_X1 \REGISTERS_reg[56][4]  ( .D(n8158), .CK(CLK), .Q(n6054), .QN(n12754)
         );
  DFF_X1 \REGISTERS_reg[56][3]  ( .D(n8157), .CK(CLK), .Q(n6053), .QN(n12753)
         );
  DFF_X1 \REGISTERS_reg[56][2]  ( .D(n8156), .CK(CLK), .Q(n6052), .QN(n12752)
         );
  DFF_X1 \REGISTERS_reg[56][1]  ( .D(n8155), .CK(CLK), .Q(n6051), .QN(n12751)
         );
  DFF_X1 \REGISTERS_reg[56][0]  ( .D(n8154), .CK(CLK), .Q(n6050), .QN(n12750)
         );
  DFF_X1 \REGISTERS_reg[57][31]  ( .D(n8153), .CK(CLK), .Q(n6049), .QN(n12717)
         );
  DFF_X1 \REGISTERS_reg[57][30]  ( .D(n8152), .CK(CLK), .Q(n6048), .QN(n12716)
         );
  DFF_X1 \REGISTERS_reg[57][29]  ( .D(n8151), .CK(CLK), .Q(n6047), .QN(n12715)
         );
  DFF_X1 \REGISTERS_reg[57][28]  ( .D(n8150), .CK(CLK), .Q(n6046), .QN(n12714)
         );
  DFF_X1 \REGISTERS_reg[57][27]  ( .D(n8149), .CK(CLK), .Q(n6045), .QN(n12713)
         );
  DFF_X1 \REGISTERS_reg[57][26]  ( .D(n8148), .CK(CLK), .Q(n6044), .QN(n12712)
         );
  DFF_X1 \REGISTERS_reg[57][25]  ( .D(n8147), .CK(CLK), .Q(n6043), .QN(n12711)
         );
  DFF_X1 \REGISTERS_reg[57][24]  ( .D(n8146), .CK(CLK), .Q(n6042), .QN(n12710)
         );
  DFF_X1 \REGISTERS_reg[57][23]  ( .D(n8145), .CK(CLK), .Q(n6041), .QN(n12749)
         );
  DFF_X1 \REGISTERS_reg[57][22]  ( .D(n8144), .CK(CLK), .Q(n6040), .QN(n12748)
         );
  DFF_X1 \REGISTERS_reg[57][21]  ( .D(n8143), .CK(CLK), .Q(n6039), .QN(n12747)
         );
  DFF_X1 \REGISTERS_reg[57][20]  ( .D(n8142), .CK(CLK), .Q(n6038), .QN(n12746)
         );
  DFF_X1 \REGISTERS_reg[57][19]  ( .D(n8141), .CK(CLK), .Q(n6037), .QN(n12745)
         );
  DFF_X1 \REGISTERS_reg[57][18]  ( .D(n8140), .CK(CLK), .Q(n6036), .QN(n12744)
         );
  DFF_X1 \REGISTERS_reg[57][17]  ( .D(n8139), .CK(CLK), .Q(n6035), .QN(n12743)
         );
  DFF_X1 \REGISTERS_reg[57][16]  ( .D(n8138), .CK(CLK), .Q(n6034), .QN(n12742)
         );
  DFF_X1 \REGISTERS_reg[57][15]  ( .D(n8137), .CK(CLK), .Q(n6033), .QN(n12741)
         );
  DFF_X1 \REGISTERS_reg[57][14]  ( .D(n8136), .CK(CLK), .Q(n6032), .QN(n12740)
         );
  DFF_X1 \REGISTERS_reg[57][13]  ( .D(n8135), .CK(CLK), .Q(n6031), .QN(n12739)
         );
  DFF_X1 \REGISTERS_reg[57][12]  ( .D(n8134), .CK(CLK), .Q(n6030), .QN(n12738)
         );
  DFF_X1 \REGISTERS_reg[57][11]  ( .D(n8133), .CK(CLK), .Q(n6029), .QN(n12737)
         );
  DFF_X1 \REGISTERS_reg[57][10]  ( .D(n8132), .CK(CLK), .Q(n6028), .QN(n12736)
         );
  DFF_X1 \REGISTERS_reg[57][9]  ( .D(n8131), .CK(CLK), .Q(n6027), .QN(n12735)
         );
  DFF_X1 \REGISTERS_reg[57][8]  ( .D(n8130), .CK(CLK), .Q(n6026), .QN(n12734)
         );
  DFF_X1 \REGISTERS_reg[57][7]  ( .D(n8129), .CK(CLK), .Q(n6025), .QN(n12733)
         );
  DFF_X1 \REGISTERS_reg[57][6]  ( .D(n8128), .CK(CLK), .Q(n6024), .QN(n12732)
         );
  DFF_X1 \REGISTERS_reg[57][5]  ( .D(n8127), .CK(CLK), .Q(n6023), .QN(n12731)
         );
  DFF_X1 \REGISTERS_reg[57][4]  ( .D(n8126), .CK(CLK), .Q(n6022), .QN(n12730)
         );
  DFF_X1 \REGISTERS_reg[57][3]  ( .D(n8125), .CK(CLK), .Q(n6021), .QN(n12729)
         );
  DFF_X1 \REGISTERS_reg[57][2]  ( .D(n8124), .CK(CLK), .Q(n6020), .QN(n12728)
         );
  DFF_X1 \REGISTERS_reg[57][1]  ( .D(n8123), .CK(CLK), .Q(n6019), .QN(n12727)
         );
  DFF_X1 \REGISTERS_reg[57][0]  ( .D(n8122), .CK(CLK), .Q(n6018), .QN(n12726)
         );
  DFF_X1 \REGISTERS_reg[59][31]  ( .D(n8089), .CK(CLK), .Q(n5985), .QN(n12837)
         );
  DFF_X1 \REGISTERS_reg[59][30]  ( .D(n8088), .CK(CLK), .Q(n5984), .QN(n12836)
         );
  DFF_X1 \REGISTERS_reg[59][29]  ( .D(n8087), .CK(CLK), .Q(n5983), .QN(n12835)
         );
  DFF_X1 \REGISTERS_reg[59][28]  ( .D(n8086), .CK(CLK), .Q(n5982), .QN(n12834)
         );
  DFF_X1 \REGISTERS_reg[59][27]  ( .D(n8085), .CK(CLK), .Q(n5981), .QN(n12833)
         );
  DFF_X1 \REGISTERS_reg[59][26]  ( .D(n8084), .CK(CLK), .Q(n5980), .QN(n12832)
         );
  DFF_X1 \REGISTERS_reg[59][25]  ( .D(n8083), .CK(CLK), .Q(n5979), .QN(n12831)
         );
  DFF_X1 \REGISTERS_reg[59][24]  ( .D(n8082), .CK(CLK), .Q(n5978), .QN(n12830)
         );
  DFF_X1 \REGISTERS_reg[59][23]  ( .D(n8081), .CK(CLK), .Q(n5977), .QN(n12829)
         );
  DFF_X1 \REGISTERS_reg[59][22]  ( .D(n8080), .CK(CLK), .Q(n5976), .QN(n12828)
         );
  DFF_X1 \REGISTERS_reg[59][21]  ( .D(n8079), .CK(CLK), .Q(n5975), .QN(n12827)
         );
  DFF_X1 \REGISTERS_reg[59][20]  ( .D(n8078), .CK(CLK), .Q(n5974), .QN(n12826)
         );
  DFF_X1 \REGISTERS_reg[59][19]  ( .D(n8077), .CK(CLK), .Q(n5973), .QN(n12825)
         );
  DFF_X1 \REGISTERS_reg[59][18]  ( .D(n8076), .CK(CLK), .Q(n5972), .QN(n12824)
         );
  DFF_X1 \REGISTERS_reg[59][17]  ( .D(n8075), .CK(CLK), .Q(n5971), .QN(n12823)
         );
  DFF_X1 \REGISTERS_reg[59][16]  ( .D(n8074), .CK(CLK), .Q(n5970), .QN(n12822)
         );
  DFF_X1 \REGISTERS_reg[59][15]  ( .D(n8073), .CK(CLK), .Q(n5969), .QN(n12821)
         );
  DFF_X1 \REGISTERS_reg[59][14]  ( .D(n8072), .CK(CLK), .Q(n5968), .QN(n12820)
         );
  DFF_X1 \REGISTERS_reg[59][13]  ( .D(n8071), .CK(CLK), .Q(n5967), .QN(n12819)
         );
  DFF_X1 \REGISTERS_reg[59][12]  ( .D(n8070), .CK(CLK), .Q(n5966), .QN(n12818)
         );
  DFF_X1 \REGISTERS_reg[59][11]  ( .D(n8069), .CK(CLK), .Q(n5965), .QN(n12817)
         );
  DFF_X1 \REGISTERS_reg[59][10]  ( .D(n8068), .CK(CLK), .Q(n5964), .QN(n12816)
         );
  DFF_X1 \REGISTERS_reg[59][9]  ( .D(n8067), .CK(CLK), .Q(n5963), .QN(n12815)
         );
  DFF_X1 \REGISTERS_reg[59][8]  ( .D(n8066), .CK(CLK), .Q(n5962), .QN(n12814)
         );
  DFF_X1 \REGISTERS_reg[59][7]  ( .D(n8065), .CK(CLK), .Q(n5961), .QN(n12813)
         );
  DFF_X1 \REGISTERS_reg[59][6]  ( .D(n8064), .CK(CLK), .Q(n5960), .QN(n12812)
         );
  DFF_X1 \REGISTERS_reg[59][5]  ( .D(n8063), .CK(CLK), .Q(n5959), .QN(n12811)
         );
  DFF_X1 \REGISTERS_reg[59][4]  ( .D(n8062), .CK(CLK), .Q(n5958), .QN(n12810)
         );
  DFF_X1 \REGISTERS_reg[59][3]  ( .D(n8061), .CK(CLK), .Q(n5957), .QN(n12809)
         );
  DFF_X1 \REGISTERS_reg[59][2]  ( .D(n8060), .CK(CLK), .Q(n5956), .QN(n12808)
         );
  DFF_X1 \REGISTERS_reg[59][1]  ( .D(n8059), .CK(CLK), .Q(n5955), .QN(n12807)
         );
  DFF_X1 \REGISTERS_reg[59][0]  ( .D(n8058), .CK(CLK), .Q(n5954), .QN(n12806)
         );
  DFF_X1 \REGISTERS_reg[60][31]  ( .D(n8057), .CK(CLK), .QN(n15206) );
  DFF_X1 \REGISTERS_reg[60][30]  ( .D(n8056), .CK(CLK), .QN(n15207) );
  DFF_X1 \REGISTERS_reg[60][29]  ( .D(n8055), .CK(CLK), .QN(n15208) );
  DFF_X1 \REGISTERS_reg[60][28]  ( .D(n8054), .CK(CLK), .QN(n15209) );
  DFF_X1 \REGISTERS_reg[60][27]  ( .D(n8053), .CK(CLK), .QN(n15210) );
  DFF_X1 \REGISTERS_reg[60][26]  ( .D(n8052), .CK(CLK), .QN(n15211) );
  DFF_X1 \REGISTERS_reg[60][25]  ( .D(n8051), .CK(CLK), .QN(n15212) );
  DFF_X1 \REGISTERS_reg[60][24]  ( .D(n8050), .CK(CLK), .QN(n15213) );
  DFF_X1 \REGISTERS_reg[60][23]  ( .D(n8049), .CK(CLK), .QN(n15214) );
  DFF_X1 \REGISTERS_reg[60][22]  ( .D(n8048), .CK(CLK), .QN(n15215) );
  DFF_X1 \REGISTERS_reg[60][21]  ( .D(n8047), .CK(CLK), .QN(n15216) );
  DFF_X1 \REGISTERS_reg[60][20]  ( .D(n8046), .CK(CLK), .QN(n15217) );
  DFF_X1 \REGISTERS_reg[60][19]  ( .D(n8045), .CK(CLK), .QN(n15218) );
  DFF_X1 \REGISTERS_reg[60][18]  ( .D(n8044), .CK(CLK), .QN(n15219) );
  DFF_X1 \REGISTERS_reg[60][17]  ( .D(n8043), .CK(CLK), .QN(n15220) );
  DFF_X1 \REGISTERS_reg[60][16]  ( .D(n8042), .CK(CLK), .QN(n15221) );
  DFF_X1 \REGISTERS_reg[60][15]  ( .D(n8041), .CK(CLK), .QN(n15222) );
  DFF_X1 \REGISTERS_reg[60][14]  ( .D(n8040), .CK(CLK), .QN(n15223) );
  DFF_X1 \REGISTERS_reg[60][13]  ( .D(n8039), .CK(CLK), .QN(n15224) );
  DFF_X1 \REGISTERS_reg[60][12]  ( .D(n8038), .CK(CLK), .QN(n15225) );
  DFF_X1 \REGISTERS_reg[60][11]  ( .D(n8037), .CK(CLK), .QN(n15226) );
  DFF_X1 \REGISTERS_reg[60][10]  ( .D(n8036), .CK(CLK), .QN(n15227) );
  DFF_X1 \REGISTERS_reg[60][9]  ( .D(n8035), .CK(CLK), .QN(n15228) );
  DFF_X1 \REGISTERS_reg[60][8]  ( .D(n8034), .CK(CLK), .QN(n15229) );
  DFF_X1 \REGISTERS_reg[60][7]  ( .D(n8033), .CK(CLK), .QN(n15230) );
  DFF_X1 \REGISTERS_reg[60][6]  ( .D(n8032), .CK(CLK), .QN(n15231) );
  DFF_X1 \REGISTERS_reg[60][5]  ( .D(n8031), .CK(CLK), .QN(n15232) );
  DFF_X1 \REGISTERS_reg[60][4]  ( .D(n8030), .CK(CLK), .QN(n15233) );
  DFF_X1 \REGISTERS_reg[60][3]  ( .D(n8029), .CK(CLK), .QN(n15234) );
  DFF_X1 \REGISTERS_reg[60][2]  ( .D(n8028), .CK(CLK), .QN(n15235) );
  DFF_X1 \REGISTERS_reg[60][1]  ( .D(n8027), .CK(CLK), .QN(n15236) );
  DFF_X1 \REGISTERS_reg[60][0]  ( .D(n8026), .CK(CLK), .QN(n15237) );
  DFF_X1 \REGISTERS_reg[61][31]  ( .D(n8025), .CK(CLK), .QN(n15238) );
  DFF_X1 \REGISTERS_reg[61][30]  ( .D(n8024), .CK(CLK), .QN(n15239) );
  DFF_X1 \REGISTERS_reg[61][29]  ( .D(n8023), .CK(CLK), .QN(n15240) );
  DFF_X1 \REGISTERS_reg[61][28]  ( .D(n8022), .CK(CLK), .QN(n15241) );
  DFF_X1 \REGISTERS_reg[61][27]  ( .D(n8021), .CK(CLK), .QN(n15242) );
  DFF_X1 \REGISTERS_reg[61][26]  ( .D(n8020), .CK(CLK), .QN(n15243) );
  DFF_X1 \REGISTERS_reg[61][25]  ( .D(n8019), .CK(CLK), .QN(n15244) );
  DFF_X1 \REGISTERS_reg[61][24]  ( .D(n8018), .CK(CLK), .QN(n15245) );
  DFF_X1 \REGISTERS_reg[61][23]  ( .D(n8017), .CK(CLK), .QN(n15246) );
  DFF_X1 \REGISTERS_reg[61][22]  ( .D(n8016), .CK(CLK), .QN(n15247) );
  DFF_X1 \REGISTERS_reg[61][21]  ( .D(n8015), .CK(CLK), .QN(n15248) );
  DFF_X1 \REGISTERS_reg[61][20]  ( .D(n8014), .CK(CLK), .QN(n15249) );
  DFF_X1 \REGISTERS_reg[61][19]  ( .D(n8013), .CK(CLK), .QN(n15250) );
  DFF_X1 \REGISTERS_reg[61][18]  ( .D(n8012), .CK(CLK), .QN(n15251) );
  DFF_X1 \REGISTERS_reg[61][17]  ( .D(n8011), .CK(CLK), .QN(n15252) );
  DFF_X1 \REGISTERS_reg[61][16]  ( .D(n8010), .CK(CLK), .QN(n15253) );
  DFF_X1 \REGISTERS_reg[61][15]  ( .D(n8009), .CK(CLK), .QN(n15254) );
  DFF_X1 \REGISTERS_reg[61][14]  ( .D(n8008), .CK(CLK), .QN(n15255) );
  DFF_X1 \REGISTERS_reg[61][13]  ( .D(n8007), .CK(CLK), .QN(n15256) );
  DFF_X1 \REGISTERS_reg[61][12]  ( .D(n8006), .CK(CLK), .QN(n15257) );
  DFF_X1 \REGISTERS_reg[61][11]  ( .D(n8005), .CK(CLK), .QN(n15258) );
  DFF_X1 \REGISTERS_reg[61][10]  ( .D(n8004), .CK(CLK), .QN(n15259) );
  DFF_X1 \REGISTERS_reg[61][9]  ( .D(n8003), .CK(CLK), .QN(n15260) );
  DFF_X1 \REGISTERS_reg[61][8]  ( .D(n8002), .CK(CLK), .QN(n15261) );
  DFF_X1 \REGISTERS_reg[61][7]  ( .D(n8001), .CK(CLK), .QN(n15262) );
  DFF_X1 \REGISTERS_reg[61][6]  ( .D(n8000), .CK(CLK), .QN(n15263) );
  DFF_X1 \REGISTERS_reg[61][5]  ( .D(n7999), .CK(CLK), .QN(n15264) );
  DFF_X1 \REGISTERS_reg[61][4]  ( .D(n7998), .CK(CLK), .QN(n15265) );
  DFF_X1 \REGISTERS_reg[61][3]  ( .D(n7997), .CK(CLK), .QN(n15266) );
  DFF_X1 \REGISTERS_reg[61][2]  ( .D(n7996), .CK(CLK), .QN(n15267) );
  DFF_X1 \REGISTERS_reg[61][1]  ( .D(n7995), .CK(CLK), .QN(n15268) );
  DFF_X1 \REGISTERS_reg[61][0]  ( .D(n7994), .CK(CLK), .QN(n15269) );
  DFF_X1 \REGISTERS_reg[62][31]  ( .D(n7993), .CK(CLK), .QN(n15270) );
  DFF_X1 \REGISTERS_reg[62][30]  ( .D(n7992), .CK(CLK), .QN(n15271) );
  DFF_X1 \REGISTERS_reg[62][29]  ( .D(n7991), .CK(CLK), .QN(n15272) );
  DFF_X1 \REGISTERS_reg[62][28]  ( .D(n7990), .CK(CLK), .QN(n15273) );
  DFF_X1 \REGISTERS_reg[62][27]  ( .D(n7989), .CK(CLK), .QN(n15274) );
  DFF_X1 \REGISTERS_reg[62][26]  ( .D(n7988), .CK(CLK), .QN(n15275) );
  DFF_X1 \REGISTERS_reg[62][25]  ( .D(n7987), .CK(CLK), .QN(n15276) );
  DFF_X1 \REGISTERS_reg[62][24]  ( .D(n7986), .CK(CLK), .QN(n15277) );
  DFF_X1 \REGISTERS_reg[62][23]  ( .D(n7985), .CK(CLK), .QN(n15278) );
  DFF_X1 \REGISTERS_reg[62][22]  ( .D(n7984), .CK(CLK), .QN(n15279) );
  DFF_X1 \REGISTERS_reg[62][21]  ( .D(n7983), .CK(CLK), .QN(n15280) );
  DFF_X1 \REGISTERS_reg[62][20]  ( .D(n7982), .CK(CLK), .QN(n15281) );
  DFF_X1 \REGISTERS_reg[62][19]  ( .D(n7981), .CK(CLK), .QN(n15282) );
  DFF_X1 \REGISTERS_reg[62][18]  ( .D(n7980), .CK(CLK), .QN(n15283) );
  DFF_X1 \REGISTERS_reg[62][17]  ( .D(n7979), .CK(CLK), .QN(n15284) );
  DFF_X1 \REGISTERS_reg[62][16]  ( .D(n7978), .CK(CLK), .QN(n15285) );
  DFF_X1 \REGISTERS_reg[62][15]  ( .D(n7977), .CK(CLK), .QN(n15286) );
  DFF_X1 \REGISTERS_reg[62][14]  ( .D(n7976), .CK(CLK), .QN(n15287) );
  DFF_X1 \REGISTERS_reg[62][13]  ( .D(n7975), .CK(CLK), .QN(n15288) );
  DFF_X1 \REGISTERS_reg[62][12]  ( .D(n7974), .CK(CLK), .QN(n15289) );
  DFF_X1 \REGISTERS_reg[62][11]  ( .D(n7973), .CK(CLK), .QN(n15290) );
  DFF_X1 \REGISTERS_reg[62][10]  ( .D(n7972), .CK(CLK), .QN(n15291) );
  DFF_X1 \REGISTERS_reg[62][9]  ( .D(n7971), .CK(CLK), .QN(n15292) );
  DFF_X1 \REGISTERS_reg[62][8]  ( .D(n7970), .CK(CLK), .QN(n15293) );
  DFF_X1 \REGISTERS_reg[62][7]  ( .D(n7969), .CK(CLK), .QN(n15294) );
  DFF_X1 \REGISTERS_reg[62][6]  ( .D(n7968), .CK(CLK), .QN(n15295) );
  DFF_X1 \REGISTERS_reg[62][5]  ( .D(n7967), .CK(CLK), .QN(n15296) );
  DFF_X1 \REGISTERS_reg[62][4]  ( .D(n7966), .CK(CLK), .QN(n15297) );
  DFF_X1 \REGISTERS_reg[62][3]  ( .D(n7965), .CK(CLK), .QN(n15298) );
  DFF_X1 \REGISTERS_reg[62][2]  ( .D(n7964), .CK(CLK), .QN(n15299) );
  DFF_X1 \REGISTERS_reg[62][1]  ( .D(n7963), .CK(CLK), .QN(n15300) );
  DFF_X1 \REGISTERS_reg[62][0]  ( .D(n7962), .CK(CLK), .QN(n15301) );
  DFF_X1 \REGISTERS_reg[64][31]  ( .D(n7929), .CK(CLK), .Q(n5921), .QN(n12805)
         );
  DFF_X1 \REGISTERS_reg[64][30]  ( .D(n7928), .CK(CLK), .Q(n5920), .QN(n12804)
         );
  DFF_X1 \REGISTERS_reg[64][29]  ( .D(n7927), .CK(CLK), .Q(n5919), .QN(n12803)
         );
  DFF_X1 \REGISTERS_reg[64][28]  ( .D(n7926), .CK(CLK), .Q(n5918), .QN(n12802)
         );
  DFF_X1 \REGISTERS_reg[64][27]  ( .D(n7925), .CK(CLK), .Q(n5917), .QN(n12801)
         );
  DFF_X1 \REGISTERS_reg[64][26]  ( .D(n7924), .CK(CLK), .Q(n5916), .QN(n12800)
         );
  DFF_X1 \REGISTERS_reg[64][25]  ( .D(n7923), .CK(CLK), .Q(n5915), .QN(n12799)
         );
  DFF_X1 \REGISTERS_reg[64][24]  ( .D(n7922), .CK(CLK), .Q(n5914), .QN(n12798)
         );
  DFF_X1 \REGISTERS_reg[64][23]  ( .D(n7921), .CK(CLK), .Q(n5913), .QN(n12797)
         );
  DFF_X1 \REGISTERS_reg[64][22]  ( .D(n7920), .CK(CLK), .Q(n5912), .QN(n12796)
         );
  DFF_X1 \REGISTERS_reg[64][21]  ( .D(n7919), .CK(CLK), .Q(n5911), .QN(n12795)
         );
  DFF_X1 \REGISTERS_reg[64][20]  ( .D(n7918), .CK(CLK), .Q(n5910), .QN(n12794)
         );
  DFF_X1 \REGISTERS_reg[64][19]  ( .D(n7917), .CK(CLK), .Q(n5909), .QN(n12793)
         );
  DFF_X1 \REGISTERS_reg[64][18]  ( .D(n7916), .CK(CLK), .Q(n5908), .QN(n12792)
         );
  DFF_X1 \REGISTERS_reg[64][17]  ( .D(n7915), .CK(CLK), .Q(n5907), .QN(n12791)
         );
  DFF_X1 \REGISTERS_reg[64][16]  ( .D(n7914), .CK(CLK), .Q(n5906), .QN(n12790)
         );
  DFF_X1 \REGISTERS_reg[64][15]  ( .D(n7913), .CK(CLK), .Q(n5905), .QN(n12789)
         );
  DFF_X1 \REGISTERS_reg[64][14]  ( .D(n7912), .CK(CLK), .Q(n5904), .QN(n12788)
         );
  DFF_X1 \REGISTERS_reg[64][13]  ( .D(n7911), .CK(CLK), .Q(n5903), .QN(n12787)
         );
  DFF_X1 \REGISTERS_reg[64][12]  ( .D(n7910), .CK(CLK), .Q(n5902), .QN(n12786)
         );
  DFF_X1 \REGISTERS_reg[64][11]  ( .D(n7909), .CK(CLK), .Q(n5901), .QN(n12785)
         );
  DFF_X1 \REGISTERS_reg[64][10]  ( .D(n7908), .CK(CLK), .Q(n5900), .QN(n12784)
         );
  DFF_X1 \REGISTERS_reg[64][9]  ( .D(n7907), .CK(CLK), .Q(n5899), .QN(n12783)
         );
  DFF_X1 \REGISTERS_reg[64][8]  ( .D(n7906), .CK(CLK), .Q(n5898), .QN(n12782)
         );
  DFF_X1 \REGISTERS_reg[64][7]  ( .D(n7905), .CK(CLK), .Q(n5897), .QN(n12781)
         );
  DFF_X1 \REGISTERS_reg[64][6]  ( .D(n7904), .CK(CLK), .Q(n5896), .QN(n12780)
         );
  DFF_X1 \REGISTERS_reg[64][5]  ( .D(n7903), .CK(CLK), .Q(n5895), .QN(n12779)
         );
  DFF_X1 \REGISTERS_reg[64][4]  ( .D(n7902), .CK(CLK), .Q(n5894), .QN(n12778)
         );
  DFF_X1 \REGISTERS_reg[64][3]  ( .D(n7901), .CK(CLK), .Q(n5893), .QN(n12777)
         );
  DFF_X1 \REGISTERS_reg[64][2]  ( .D(n7900), .CK(CLK), .Q(n5892), .QN(n12776)
         );
  DFF_X1 \REGISTERS_reg[64][1]  ( .D(n7899), .CK(CLK), .Q(n5891), .QN(n12775)
         );
  DFF_X1 \REGISTERS_reg[64][0]  ( .D(n7898), .CK(CLK), .Q(n5890), .QN(n12774)
         );
  DFF_X1 \REGISTERS_reg[65][31]  ( .D(n7897), .CK(CLK), .QN(n15334) );
  DFF_X1 \REGISTERS_reg[65][30]  ( .D(n7896), .CK(CLK), .QN(n15335) );
  DFF_X1 \REGISTERS_reg[65][29]  ( .D(n7895), .CK(CLK), .QN(n15336) );
  DFF_X1 \REGISTERS_reg[65][28]  ( .D(n7894), .CK(CLK), .QN(n15337) );
  DFF_X1 \REGISTERS_reg[65][27]  ( .D(n7893), .CK(CLK), .QN(n15338) );
  DFF_X1 \REGISTERS_reg[65][26]  ( .D(n7892), .CK(CLK), .QN(n15339) );
  DFF_X1 \REGISTERS_reg[65][25]  ( .D(n7891), .CK(CLK), .QN(n15340) );
  DFF_X1 \REGISTERS_reg[65][24]  ( .D(n7890), .CK(CLK), .QN(n15341) );
  DFF_X1 \REGISTERS_reg[65][23]  ( .D(n7889), .CK(CLK), .QN(n15342) );
  DFF_X1 \REGISTERS_reg[65][22]  ( .D(n7888), .CK(CLK), .QN(n15343) );
  DFF_X1 \REGISTERS_reg[65][21]  ( .D(n7887), .CK(CLK), .QN(n15344) );
  DFF_X1 \REGISTERS_reg[65][20]  ( .D(n7886), .CK(CLK), .QN(n15345) );
  DFF_X1 \REGISTERS_reg[65][19]  ( .D(n7885), .CK(CLK), .QN(n15346) );
  DFF_X1 \REGISTERS_reg[65][18]  ( .D(n7884), .CK(CLK), .QN(n15347) );
  DFF_X1 \REGISTERS_reg[65][17]  ( .D(n7883), .CK(CLK), .QN(n15348) );
  DFF_X1 \REGISTERS_reg[65][16]  ( .D(n7882), .CK(CLK), .QN(n15349) );
  DFF_X1 \REGISTERS_reg[65][15]  ( .D(n7881), .CK(CLK), .QN(n15350) );
  DFF_X1 \REGISTERS_reg[65][14]  ( .D(n7880), .CK(CLK), .QN(n15351) );
  DFF_X1 \REGISTERS_reg[65][13]  ( .D(n7879), .CK(CLK), .QN(n15352) );
  DFF_X1 \REGISTERS_reg[65][12]  ( .D(n7878), .CK(CLK), .QN(n15353) );
  DFF_X1 \REGISTERS_reg[65][11]  ( .D(n7877), .CK(CLK), .QN(n15354) );
  DFF_X1 \REGISTERS_reg[65][10]  ( .D(n7876), .CK(CLK), .QN(n15355) );
  DFF_X1 \REGISTERS_reg[65][9]  ( .D(n7875), .CK(CLK), .QN(n15356) );
  DFF_X1 \REGISTERS_reg[65][8]  ( .D(n7874), .CK(CLK), .QN(n15357) );
  DFF_X1 \REGISTERS_reg[65][7]  ( .D(n7873), .CK(CLK), .QN(n15358) );
  DFF_X1 \REGISTERS_reg[65][6]  ( .D(n7872), .CK(CLK), .QN(n15359) );
  DFF_X1 \REGISTERS_reg[65][5]  ( .D(n7871), .CK(CLK), .QN(n15360) );
  DFF_X1 \REGISTERS_reg[65][4]  ( .D(n7870), .CK(CLK), .QN(n15361) );
  DFF_X1 \REGISTERS_reg[65][3]  ( .D(n7869), .CK(CLK), .QN(n15362) );
  DFF_X1 \REGISTERS_reg[65][2]  ( .D(n7868), .CK(CLK), .QN(n15363) );
  DFF_X1 \REGISTERS_reg[65][1]  ( .D(n7867), .CK(CLK), .QN(n15364) );
  DFF_X1 \REGISTERS_reg[65][0]  ( .D(n7866), .CK(CLK), .QN(n15365) );
  DFF_X1 \REGISTERS_reg[66][31]  ( .D(n7865), .CK(CLK), .QN(n15366) );
  DFF_X1 \REGISTERS_reg[66][30]  ( .D(n7864), .CK(CLK), .QN(n15367) );
  DFF_X1 \REGISTERS_reg[66][29]  ( .D(n7863), .CK(CLK), .QN(n15368) );
  DFF_X1 \REGISTERS_reg[66][28]  ( .D(n7862), .CK(CLK), .QN(n15369) );
  DFF_X1 \REGISTERS_reg[66][27]  ( .D(n7861), .CK(CLK), .QN(n15370) );
  DFF_X1 \REGISTERS_reg[66][26]  ( .D(n7860), .CK(CLK), .QN(n15371) );
  DFF_X1 \REGISTERS_reg[66][25]  ( .D(n7859), .CK(CLK), .QN(n15372) );
  DFF_X1 \REGISTERS_reg[66][24]  ( .D(n7858), .CK(CLK), .QN(n15373) );
  DFF_X1 \REGISTERS_reg[66][23]  ( .D(n7857), .CK(CLK), .QN(n15374) );
  DFF_X1 \REGISTERS_reg[66][22]  ( .D(n7856), .CK(CLK), .QN(n15375) );
  DFF_X1 \REGISTERS_reg[66][21]  ( .D(n7855), .CK(CLK), .QN(n15376) );
  DFF_X1 \REGISTERS_reg[66][20]  ( .D(n7854), .CK(CLK), .QN(n15377) );
  DFF_X1 \REGISTERS_reg[66][19]  ( .D(n7853), .CK(CLK), .QN(n15378) );
  DFF_X1 \REGISTERS_reg[66][18]  ( .D(n7852), .CK(CLK), .QN(n15379) );
  DFF_X1 \REGISTERS_reg[66][17]  ( .D(n7851), .CK(CLK), .QN(n15380) );
  DFF_X1 \REGISTERS_reg[66][16]  ( .D(n7850), .CK(CLK), .QN(n15381) );
  DFF_X1 \REGISTERS_reg[66][15]  ( .D(n7849), .CK(CLK), .QN(n15382) );
  DFF_X1 \REGISTERS_reg[66][14]  ( .D(n7848), .CK(CLK), .QN(n15383) );
  DFF_X1 \REGISTERS_reg[66][13]  ( .D(n7847), .CK(CLK), .QN(n15384) );
  DFF_X1 \REGISTERS_reg[66][12]  ( .D(n7846), .CK(CLK), .QN(n15385) );
  DFF_X1 \REGISTERS_reg[66][11]  ( .D(n7845), .CK(CLK), .QN(n15386) );
  DFF_X1 \REGISTERS_reg[66][10]  ( .D(n7844), .CK(CLK), .QN(n15387) );
  DFF_X1 \REGISTERS_reg[66][9]  ( .D(n7843), .CK(CLK), .QN(n15388) );
  DFF_X1 \REGISTERS_reg[66][8]  ( .D(n7842), .CK(CLK), .QN(n15389) );
  DFF_X1 \REGISTERS_reg[66][7]  ( .D(n7841), .CK(CLK), .QN(n15390) );
  DFF_X1 \REGISTERS_reg[66][6]  ( .D(n7840), .CK(CLK), .QN(n15391) );
  DFF_X1 \REGISTERS_reg[66][5]  ( .D(n7839), .CK(CLK), .QN(n15392) );
  DFF_X1 \REGISTERS_reg[66][4]  ( .D(n7838), .CK(CLK), .QN(n15393) );
  DFF_X1 \REGISTERS_reg[66][3]  ( .D(n7837), .CK(CLK), .QN(n15394) );
  DFF_X1 \REGISTERS_reg[66][2]  ( .D(n7836), .CK(CLK), .QN(n15395) );
  DFF_X1 \REGISTERS_reg[66][1]  ( .D(n7835), .CK(CLK), .QN(n15396) );
  DFF_X1 \REGISTERS_reg[66][0]  ( .D(n7834), .CK(CLK), .QN(n15397) );
  DFF_X1 \REGISTERS_reg[69][31]  ( .D(n7769), .CK(CLK), .QN(n15462) );
  DFF_X1 \REGISTERS_reg[69][30]  ( .D(n7768), .CK(CLK), .QN(n15463) );
  DFF_X1 \REGISTERS_reg[69][29]  ( .D(n7767), .CK(CLK), .QN(n15464) );
  DFF_X1 \REGISTERS_reg[69][28]  ( .D(n7766), .CK(CLK), .QN(n15465) );
  DFF_X1 \REGISTERS_reg[69][27]  ( .D(n7765), .CK(CLK), .QN(n15466) );
  DFF_X1 \REGISTERS_reg[69][26]  ( .D(n7764), .CK(CLK), .QN(n15467) );
  DFF_X1 \REGISTERS_reg[69][25]  ( .D(n7763), .CK(CLK), .QN(n15468) );
  DFF_X1 \REGISTERS_reg[69][24]  ( .D(n7762), .CK(CLK), .QN(n15469) );
  DFF_X1 \REGISTERS_reg[69][23]  ( .D(n7761), .CK(CLK), .QN(n15470) );
  DFF_X1 \REGISTERS_reg[69][22]  ( .D(n7760), .CK(CLK), .QN(n15471) );
  DFF_X1 \REGISTERS_reg[69][21]  ( .D(n7759), .CK(CLK), .QN(n15472) );
  DFF_X1 \REGISTERS_reg[69][20]  ( .D(n7758), .CK(CLK), .QN(n15473) );
  DFF_X1 \REGISTERS_reg[69][19]  ( .D(n7757), .CK(CLK), .QN(n15474) );
  DFF_X1 \REGISTERS_reg[69][18]  ( .D(n7756), .CK(CLK), .QN(n15475) );
  DFF_X1 \REGISTERS_reg[69][17]  ( .D(n7755), .CK(CLK), .QN(n15476) );
  DFF_X1 \REGISTERS_reg[69][16]  ( .D(n7754), .CK(CLK), .QN(n15477) );
  DFF_X1 \REGISTERS_reg[69][15]  ( .D(n7753), .CK(CLK), .QN(n15478) );
  DFF_X1 \REGISTERS_reg[69][14]  ( .D(n7752), .CK(CLK), .QN(n15479) );
  DFF_X1 \REGISTERS_reg[69][13]  ( .D(n7751), .CK(CLK), .QN(n15480) );
  DFF_X1 \REGISTERS_reg[69][12]  ( .D(n7750), .CK(CLK), .QN(n15481) );
  DFF_X1 \REGISTERS_reg[69][11]  ( .D(n7749), .CK(CLK), .QN(n15482) );
  DFF_X1 \REGISTERS_reg[69][10]  ( .D(n7748), .CK(CLK), .QN(n15483) );
  DFF_X1 \REGISTERS_reg[69][9]  ( .D(n7747), .CK(CLK), .QN(n15484) );
  DFF_X1 \REGISTERS_reg[69][8]  ( .D(n7746), .CK(CLK), .QN(n15485) );
  DFF_X1 \REGISTERS_reg[69][7]  ( .D(n7745), .CK(CLK), .QN(n15486) );
  DFF_X1 \REGISTERS_reg[69][6]  ( .D(n7744), .CK(CLK), .QN(n15487) );
  DFF_X1 \REGISTERS_reg[69][5]  ( .D(n7743), .CK(CLK), .QN(n15488) );
  DFF_X1 \REGISTERS_reg[69][4]  ( .D(n7742), .CK(CLK), .QN(n15489) );
  DFF_X1 \REGISTERS_reg[69][3]  ( .D(n7741), .CK(CLK), .QN(n15490) );
  DFF_X1 \REGISTERS_reg[69][2]  ( .D(n7740), .CK(CLK), .QN(n15491) );
  DFF_X1 \REGISTERS_reg[69][1]  ( .D(n7739), .CK(CLK), .QN(n15492) );
  DFF_X1 \REGISTERS_reg[69][0]  ( .D(n7738), .CK(CLK), .QN(n15493) );
  DFF_X1 \REGISTERS_reg[70][31]  ( .D(n7737), .CK(CLK), .QN(n15494) );
  DFF_X1 \REGISTERS_reg[70][30]  ( .D(n7736), .CK(CLK), .QN(n15495) );
  DFF_X1 \REGISTERS_reg[70][29]  ( .D(n7735), .CK(CLK), .QN(n15496) );
  DFF_X1 \REGISTERS_reg[70][28]  ( .D(n7734), .CK(CLK), .QN(n15497) );
  DFF_X1 \REGISTERS_reg[70][27]  ( .D(n7733), .CK(CLK), .QN(n15498) );
  DFF_X1 \REGISTERS_reg[70][26]  ( .D(n7732), .CK(CLK), .QN(n15499) );
  DFF_X1 \REGISTERS_reg[70][25]  ( .D(n7731), .CK(CLK), .QN(n15500) );
  DFF_X1 \REGISTERS_reg[70][24]  ( .D(n7730), .CK(CLK), .QN(n15501) );
  DFF_X1 \REGISTERS_reg[70][23]  ( .D(n7729), .CK(CLK), .QN(n15502) );
  DFF_X1 \REGISTERS_reg[70][22]  ( .D(n7728), .CK(CLK), .QN(n15503) );
  DFF_X1 \REGISTERS_reg[70][21]  ( .D(n7727), .CK(CLK), .QN(n15504) );
  DFF_X1 \REGISTERS_reg[70][20]  ( .D(n7726), .CK(CLK), .QN(n15505) );
  DFF_X1 \REGISTERS_reg[70][19]  ( .D(n7725), .CK(CLK), .QN(n15506) );
  DFF_X1 \REGISTERS_reg[70][18]  ( .D(n7724), .CK(CLK), .QN(n15507) );
  DFF_X1 \REGISTERS_reg[70][17]  ( .D(n7723), .CK(CLK), .QN(n15508) );
  DFF_X1 \REGISTERS_reg[70][16]  ( .D(n7722), .CK(CLK), .QN(n15509) );
  DFF_X1 \REGISTERS_reg[70][15]  ( .D(n7721), .CK(CLK), .QN(n15510) );
  DFF_X1 \REGISTERS_reg[70][14]  ( .D(n7720), .CK(CLK), .QN(n15511) );
  DFF_X1 \REGISTERS_reg[70][13]  ( .D(n7719), .CK(CLK), .QN(n15512) );
  DFF_X1 \REGISTERS_reg[70][12]  ( .D(n7718), .CK(CLK), .QN(n15513) );
  DFF_X1 \REGISTERS_reg[70][11]  ( .D(n7717), .CK(CLK), .QN(n15514) );
  DFF_X1 \REGISTERS_reg[70][10]  ( .D(n7716), .CK(CLK), .QN(n15515) );
  DFF_X1 \REGISTERS_reg[70][9]  ( .D(n7715), .CK(CLK), .QN(n15516) );
  DFF_X1 \REGISTERS_reg[70][8]  ( .D(n7714), .CK(CLK), .QN(n15517) );
  DFF_X1 \REGISTERS_reg[70][7]  ( .D(n7713), .CK(CLK), .QN(n15518) );
  DFF_X1 \REGISTERS_reg[70][6]  ( .D(n7712), .CK(CLK), .QN(n15519) );
  DFF_X1 \REGISTERS_reg[70][5]  ( .D(n7711), .CK(CLK), .QN(n15520) );
  DFF_X1 \REGISTERS_reg[70][4]  ( .D(n7710), .CK(CLK), .QN(n15521) );
  DFF_X1 \REGISTERS_reg[70][3]  ( .D(n7709), .CK(CLK), .QN(n15522) );
  DFF_X1 \REGISTERS_reg[70][2]  ( .D(n7708), .CK(CLK), .QN(n15523) );
  DFF_X1 \REGISTERS_reg[70][1]  ( .D(n7707), .CK(CLK), .QN(n15524) );
  DFF_X1 \REGISTERS_reg[70][0]  ( .D(n7706), .CK(CLK), .QN(n15525) );
  DFF_X1 \REGISTERS_reg[71][31]  ( .D(n7705), .CK(CLK), .QN(n15526) );
  DFF_X1 \REGISTERS_reg[71][30]  ( .D(n7704), .CK(CLK), .QN(n15527) );
  DFF_X1 \REGISTERS_reg[71][29]  ( .D(n7703), .CK(CLK), .QN(n15528) );
  DFF_X1 \REGISTERS_reg[71][28]  ( .D(n7702), .CK(CLK), .QN(n15529) );
  DFF_X1 \REGISTERS_reg[71][27]  ( .D(n7701), .CK(CLK), .QN(n15530) );
  DFF_X1 \REGISTERS_reg[71][26]  ( .D(n7700), .CK(CLK), .QN(n15531) );
  DFF_X1 \REGISTERS_reg[71][25]  ( .D(n7699), .CK(CLK), .QN(n15532) );
  DFF_X1 \REGISTERS_reg[71][24]  ( .D(n7698), .CK(CLK), .QN(n15533) );
  DFF_X1 \REGISTERS_reg[71][23]  ( .D(n7697), .CK(CLK), .QN(n15534) );
  DFF_X1 \REGISTERS_reg[71][22]  ( .D(n7696), .CK(CLK), .QN(n15535) );
  DFF_X1 \REGISTERS_reg[71][21]  ( .D(n7695), .CK(CLK), .QN(n15536) );
  DFF_X1 \REGISTERS_reg[71][20]  ( .D(n7694), .CK(CLK), .QN(n15537) );
  DFF_X1 \REGISTERS_reg[71][19]  ( .D(n7693), .CK(CLK), .QN(n15538) );
  DFF_X1 \REGISTERS_reg[71][18]  ( .D(n7692), .CK(CLK), .QN(n15539) );
  DFF_X1 \REGISTERS_reg[71][17]  ( .D(n7691), .CK(CLK), .QN(n15540) );
  DFF_X1 \REGISTERS_reg[71][16]  ( .D(n7690), .CK(CLK), .QN(n15541) );
  DFF_X1 \REGISTERS_reg[71][15]  ( .D(n7689), .CK(CLK), .QN(n15542) );
  DFF_X1 \REGISTERS_reg[71][14]  ( .D(n7688), .CK(CLK), .QN(n15543) );
  DFF_X1 \REGISTERS_reg[71][13]  ( .D(n7687), .CK(CLK), .QN(n15544) );
  DFF_X1 \REGISTERS_reg[71][12]  ( .D(n7686), .CK(CLK), .QN(n15545) );
  DFF_X1 \REGISTERS_reg[71][11]  ( .D(n7685), .CK(CLK), .QN(n15546) );
  DFF_X1 \REGISTERS_reg[71][10]  ( .D(n7684), .CK(CLK), .QN(n15547) );
  DFF_X1 \REGISTERS_reg[71][9]  ( .D(n7683), .CK(CLK), .QN(n15548) );
  DFF_X1 \REGISTERS_reg[71][8]  ( .D(n7682), .CK(CLK), .QN(n15549) );
  DFF_X1 \REGISTERS_reg[71][7]  ( .D(n7681), .CK(CLK), .QN(n15550) );
  DFF_X1 \REGISTERS_reg[71][6]  ( .D(n7680), .CK(CLK), .QN(n15551) );
  DFF_X1 \REGISTERS_reg[71][5]  ( .D(n7679), .CK(CLK), .QN(n15552) );
  DFF_X1 \REGISTERS_reg[71][4]  ( .D(n7678), .CK(CLK), .QN(n15553) );
  DFF_X1 \REGISTERS_reg[71][3]  ( .D(n7677), .CK(CLK), .QN(n15554) );
  DFF_X1 \REGISTERS_reg[71][2]  ( .D(n7676), .CK(CLK), .QN(n15555) );
  DFF_X1 \REGISTERS_reg[71][1]  ( .D(n7675), .CK(CLK), .QN(n15556) );
  DFF_X1 \REGISTERS_reg[71][0]  ( .D(n7674), .CK(CLK), .QN(n15557) );
  DFF_X1 \OUT1_tri_enable_reg[31]  ( .D(n7672), .CK(CLK), .Q(n6659), .QN(n1513) );
  DFF_X1 \OUT1_tri_enable_reg[30]  ( .D(n7670), .CK(CLK), .Q(n6661), .QN(n1514) );
  DFF_X1 \OUT1_tri_enable_reg[29]  ( .D(n7668), .CK(CLK), .Q(n6663), .QN(n1515) );
  DFF_X1 \OUT1_tri_enable_reg[28]  ( .D(n7666), .CK(CLK), .Q(n6665), .QN(n1516) );
  DFF_X1 \OUT1_tri_enable_reg[27]  ( .D(n7664), .CK(CLK), .Q(n6667), .QN(n1517) );
  DFF_X1 \OUT1_tri_enable_reg[26]  ( .D(n7662), .CK(CLK), .Q(n6669), .QN(n1518) );
  DFF_X1 \OUT1_tri_enable_reg[25]  ( .D(n7660), .CK(CLK), .Q(n6671), .QN(n1519) );
  DFF_X1 \OUT1_tri_enable_reg[24]  ( .D(n7658), .CK(CLK), .Q(n6673), .QN(n1520) );
  DFF_X1 \OUT1_reg[23]  ( .D(n7657), .CK(CLK), .QN(n1457) );
  DFF_X1 \OUT1_tri_enable_reg[23]  ( .D(n7656), .CK(CLK), .Q(n6675), .QN(n1521) );
  DFF_X1 \OUT1_reg[22]  ( .D(n7655), .CK(CLK), .QN(n1458) );
  DFF_X1 \OUT1_tri_enable_reg[22]  ( .D(n7654), .CK(CLK), .Q(n6677), .QN(n1522) );
  DFF_X1 \OUT1_reg[21]  ( .D(n7653), .CK(CLK), .QN(n1459) );
  DFF_X1 \OUT1_tri_enable_reg[21]  ( .D(n7652), .CK(CLK), .Q(n6679), .QN(n1523) );
  DFF_X1 \OUT1_reg[20]  ( .D(n7651), .CK(CLK), .QN(n1460) );
  DFF_X1 \OUT1_tri_enable_reg[20]  ( .D(n7650), .CK(CLK), .Q(n6681), .QN(n1524) );
  DFF_X1 \OUT1_reg[19]  ( .D(n7649), .CK(CLK), .QN(n1461) );
  DFF_X1 \OUT1_tri_enable_reg[19]  ( .D(n7648), .CK(CLK), .Q(n6683), .QN(n1525) );
  DFF_X1 \OUT1_reg[18]  ( .D(n7647), .CK(CLK), .QN(n1462) );
  DFF_X1 \OUT1_tri_enable_reg[18]  ( .D(n7646), .CK(CLK), .Q(n6685), .QN(n1526) );
  DFF_X1 \OUT1_reg[17]  ( .D(n7645), .CK(CLK), .QN(n1463) );
  DFF_X1 \OUT1_tri_enable_reg[17]  ( .D(n7644), .CK(CLK), .Q(n6687), .QN(n1527) );
  DFF_X1 \OUT1_reg[16]  ( .D(n7643), .CK(CLK), .QN(n1464) );
  DFF_X1 \OUT1_tri_enable_reg[16]  ( .D(n7642), .CK(CLK), .Q(n6689), .QN(n1528) );
  DFF_X1 \OUT1_reg[15]  ( .D(n7641), .CK(CLK), .QN(n1465) );
  DFF_X1 \OUT1_tri_enable_reg[15]  ( .D(n7640), .CK(CLK), .Q(n6691), .QN(n1529) );
  DFF_X1 \OUT1_reg[14]  ( .D(n7639), .CK(CLK), .QN(n1466) );
  DFF_X1 \OUT1_tri_enable_reg[14]  ( .D(n7638), .CK(CLK), .Q(n6693), .QN(n1530) );
  DFF_X1 \OUT1_reg[13]  ( .D(n7637), .CK(CLK), .QN(n1467) );
  DFF_X1 \OUT1_tri_enable_reg[13]  ( .D(n7636), .CK(CLK), .Q(n6695), .QN(n1531) );
  DFF_X1 \OUT1_reg[12]  ( .D(n7635), .CK(CLK), .QN(n1468) );
  DFF_X1 \OUT1_tri_enable_reg[12]  ( .D(n7634), .CK(CLK), .Q(n6697), .QN(n1532) );
  DFF_X1 \OUT1_reg[11]  ( .D(n7633), .CK(CLK), .QN(n1469) );
  DFF_X1 \OUT1_tri_enable_reg[11]  ( .D(n7632), .CK(CLK), .Q(n6699), .QN(n1533) );
  DFF_X1 \OUT1_reg[10]  ( .D(n7631), .CK(CLK), .QN(n1470) );
  DFF_X1 \OUT1_tri_enable_reg[10]  ( .D(n7630), .CK(CLK), .Q(n6701), .QN(n1534) );
  DFF_X1 \OUT1_reg[9]  ( .D(n7629), .CK(CLK), .QN(n1471) );
  DFF_X1 \OUT1_tri_enable_reg[9]  ( .D(n7628), .CK(CLK), .Q(n6703), .QN(n1535)
         );
  DFF_X1 \OUT1_reg[8]  ( .D(n7627), .CK(CLK), .QN(n1472) );
  DFF_X1 \OUT1_tri_enable_reg[8]  ( .D(n7626), .CK(CLK), .Q(n6705), .QN(n1536)
         );
  DFF_X1 \OUT1_reg[7]  ( .D(n7625), .CK(CLK), .QN(n1473) );
  DFF_X1 \OUT1_tri_enable_reg[7]  ( .D(n7624), .CK(CLK), .Q(n6707), .QN(n1537)
         );
  DFF_X1 \OUT1_reg[6]  ( .D(n7623), .CK(CLK), .QN(n1474) );
  DFF_X1 \OUT1_tri_enable_reg[6]  ( .D(n7622), .CK(CLK), .Q(n6709), .QN(n1538)
         );
  DFF_X1 \OUT1_reg[5]  ( .D(n7621), .CK(CLK), .QN(n1475) );
  DFF_X1 \OUT1_tri_enable_reg[5]  ( .D(n7620), .CK(CLK), .Q(n6711), .QN(n1539)
         );
  DFF_X1 \OUT1_reg[4]  ( .D(n7619), .CK(CLK), .QN(n1476) );
  DFF_X1 \OUT1_tri_enable_reg[4]  ( .D(n7618), .CK(CLK), .Q(n6713), .QN(n1540)
         );
  DFF_X1 \OUT1_reg[3]  ( .D(n7617), .CK(CLK), .QN(n1477) );
  DFF_X1 \OUT1_tri_enable_reg[3]  ( .D(n7616), .CK(CLK), .Q(n6715), .QN(n1541)
         );
  DFF_X1 \OUT1_reg[2]  ( .D(n7615), .CK(CLK), .QN(n1478) );
  DFF_X1 \OUT1_tri_enable_reg[2]  ( .D(n7614), .CK(CLK), .Q(n6717), .QN(n1542)
         );
  DFF_X1 \OUT1_reg[1]  ( .D(n7613), .CK(CLK), .QN(n1479) );
  DFF_X1 \OUT1_tri_enable_reg[1]  ( .D(n7612), .CK(CLK), .Q(n6719), .QN(n1543)
         );
  DFF_X1 \OUT1_reg[0]  ( .D(n7611), .CK(CLK), .QN(n1480) );
  DFF_X1 \OUT1_tri_enable_reg[0]  ( .D(n7610), .CK(CLK), .Q(n6721), .QN(n1544)
         );
  DFF_X1 \OUT2_tri_enable_reg[31]  ( .D(n7608), .CK(CLK), .Q(n6723), .QN(n1545) );
  DFF_X1 \OUT2_tri_enable_reg[30]  ( .D(n7606), .CK(CLK), .Q(n6725), .QN(n1546) );
  DFF_X1 \OUT2_tri_enable_reg[29]  ( .D(n7604), .CK(CLK), .Q(n6727), .QN(n1547) );
  DFF_X1 \OUT2_tri_enable_reg[28]  ( .D(n7602), .CK(CLK), .Q(n6729), .QN(n1548) );
  DFF_X1 \OUT2_tri_enable_reg[27]  ( .D(n7600), .CK(CLK), .Q(n6731), .QN(n1549) );
  DFF_X1 \OUT2_tri_enable_reg[26]  ( .D(n7598), .CK(CLK), .Q(n6733), .QN(n1550) );
  DFF_X1 \OUT2_tri_enable_reg[25]  ( .D(n7596), .CK(CLK), .Q(n6735), .QN(n1551) );
  DFF_X1 \OUT2_tri_enable_reg[24]  ( .D(n7594), .CK(CLK), .Q(n6737), .QN(n1552) );
  DFF_X1 \OUT2_reg[23]  ( .D(n7593), .CK(CLK), .QN(n1489) );
  DFF_X1 \OUT2_tri_enable_reg[23]  ( .D(n7592), .CK(CLK), .Q(n6739), .QN(n1553) );
  DFF_X1 \OUT2_reg[22]  ( .D(n7591), .CK(CLK), .QN(n1490) );
  DFF_X1 \OUT2_tri_enable_reg[22]  ( .D(n7590), .CK(CLK), .Q(n6741), .QN(n1554) );
  DFF_X1 \OUT2_reg[21]  ( .D(n7589), .CK(CLK), .QN(n1491) );
  DFF_X1 \OUT2_tri_enable_reg[21]  ( .D(n7588), .CK(CLK), .Q(n6743), .QN(n1555) );
  DFF_X1 \OUT2_reg[20]  ( .D(n7587), .CK(CLK), .QN(n1492) );
  DFF_X1 \OUT2_tri_enable_reg[20]  ( .D(n7586), .CK(CLK), .Q(n6745), .QN(n1556) );
  DFF_X1 \OUT2_reg[19]  ( .D(n7585), .CK(CLK), .QN(n1493) );
  DFF_X1 \OUT2_tri_enable_reg[19]  ( .D(n7584), .CK(CLK), .Q(n6747), .QN(n1557) );
  DFF_X1 \OUT2_reg[18]  ( .D(n7583), .CK(CLK), .QN(n1494) );
  DFF_X1 \OUT2_tri_enable_reg[18]  ( .D(n7582), .CK(CLK), .Q(n6749), .QN(n1558) );
  DFF_X1 \OUT2_reg[17]  ( .D(n7581), .CK(CLK), .QN(n1495) );
  DFF_X1 \OUT2_tri_enable_reg[17]  ( .D(n7580), .CK(CLK), .Q(n6751), .QN(n1559) );
  DFF_X1 \OUT2_reg[16]  ( .D(n7579), .CK(CLK), .QN(n1496) );
  DFF_X1 \OUT2_tri_enable_reg[16]  ( .D(n7578), .CK(CLK), .Q(n6753), .QN(n1560) );
  DFF_X1 \OUT2_reg[15]  ( .D(n7577), .CK(CLK), .QN(n1497) );
  DFF_X1 \OUT2_tri_enable_reg[15]  ( .D(n7576), .CK(CLK), .Q(n6755), .QN(n1561) );
  DFF_X1 \OUT2_reg[14]  ( .D(n7575), .CK(CLK), .QN(n1498) );
  DFF_X1 \OUT2_tri_enable_reg[14]  ( .D(n7574), .CK(CLK), .Q(n6757), .QN(n1562) );
  DFF_X1 \OUT2_reg[13]  ( .D(n7573), .CK(CLK), .QN(n1499) );
  DFF_X1 \OUT2_tri_enable_reg[13]  ( .D(n7572), .CK(CLK), .Q(n6759), .QN(n1563) );
  DFF_X1 \OUT2_reg[12]  ( .D(n7571), .CK(CLK), .QN(n1500) );
  DFF_X1 \OUT2_tri_enable_reg[12]  ( .D(n7570), .CK(CLK), .Q(n6761), .QN(n1564) );
  DFF_X1 \OUT2_reg[11]  ( .D(n7569), .CK(CLK), .QN(n1501) );
  DFF_X1 \OUT2_tri_enable_reg[11]  ( .D(n7568), .CK(CLK), .Q(n6763), .QN(n1565) );
  DFF_X1 \OUT2_reg[10]  ( .D(n7567), .CK(CLK), .QN(n1502) );
  DFF_X1 \OUT2_tri_enable_reg[10]  ( .D(n7566), .CK(CLK), .Q(n6765), .QN(n1566) );
  DFF_X1 \OUT2_reg[9]  ( .D(n7565), .CK(CLK), .QN(n1503) );
  DFF_X1 \OUT2_tri_enable_reg[9]  ( .D(n7564), .CK(CLK), .Q(n6767), .QN(n1567)
         );
  DFF_X1 \OUT2_reg[8]  ( .D(n7563), .CK(CLK), .QN(n1504) );
  DFF_X1 \OUT2_tri_enable_reg[8]  ( .D(n7562), .CK(CLK), .Q(n6769), .QN(n1568)
         );
  DFF_X1 \OUT2_reg[7]  ( .D(n7561), .CK(CLK), .QN(n1505) );
  DFF_X1 \OUT2_tri_enable_reg[7]  ( .D(n7560), .CK(CLK), .Q(n6771), .QN(n1569)
         );
  DFF_X1 \OUT2_reg[6]  ( .D(n7559), .CK(CLK), .QN(n1506) );
  DFF_X1 \OUT2_tri_enable_reg[6]  ( .D(n7558), .CK(CLK), .Q(n6773), .QN(n1570)
         );
  DFF_X1 \OUT2_reg[5]  ( .D(n7557), .CK(CLK), .QN(n1507) );
  DFF_X1 \OUT2_tri_enable_reg[5]  ( .D(n7556), .CK(CLK), .Q(n6775), .QN(n1571)
         );
  DFF_X1 \OUT2_reg[4]  ( .D(n7555), .CK(CLK), .QN(n1508) );
  DFF_X1 \OUT2_tri_enable_reg[4]  ( .D(n7554), .CK(CLK), .Q(n6777), .QN(n1572)
         );
  DFF_X1 \OUT2_reg[3]  ( .D(n7553), .CK(CLK), .QN(n1509) );
  DFF_X1 \OUT2_tri_enable_reg[3]  ( .D(n7552), .CK(CLK), .Q(n6779), .QN(n1573)
         );
  DFF_X1 \OUT2_reg[2]  ( .D(n7551), .CK(CLK), .QN(n1510) );
  DFF_X1 \OUT2_tri_enable_reg[2]  ( .D(n7550), .CK(CLK), .Q(n6781), .QN(n1574)
         );
  DFF_X1 \OUT2_reg[1]  ( .D(n7549), .CK(CLK), .QN(n1511) );
  DFF_X1 \OUT2_tri_enable_reg[1]  ( .D(n7548), .CK(CLK), .Q(n6783), .QN(n1575)
         );
  DFF_X1 \OUT2_reg[0]  ( .D(n7547), .CK(CLK), .QN(n1512) );
  DFF_X1 \OUT2_tri_enable_reg[0]  ( .D(n7546), .CK(CLK), .Q(n6785), .QN(n1576)
         );
  DFF_X1 \REGISTERS_reg[48][31]  ( .D(n8441), .CK(CLK), .QN(n15923) );
  DFF_X1 \REGISTERS_reg[48][30]  ( .D(n8440), .CK(CLK), .QN(n15924) );
  DFF_X1 \REGISTERS_reg[48][29]  ( .D(n8439), .CK(CLK), .QN(n15925) );
  DFF_X1 \REGISTERS_reg[48][28]  ( .D(n8438), .CK(CLK), .QN(n15926) );
  DFF_X1 \REGISTERS_reg[48][27]  ( .D(n8437), .CK(CLK), .QN(n15927) );
  DFF_X1 \REGISTERS_reg[48][26]  ( .D(n8436), .CK(CLK), .QN(n15928) );
  DFF_X1 \REGISTERS_reg[48][25]  ( .D(n8435), .CK(CLK), .QN(n15929) );
  DFF_X1 \REGISTERS_reg[48][24]  ( .D(n8434), .CK(CLK), .QN(n15930) );
  DFF_X1 \REGISTERS_reg[48][23]  ( .D(n8433), .CK(CLK), .QN(n15947) );
  DFF_X1 \REGISTERS_reg[48][22]  ( .D(n8432), .CK(CLK), .QN(n15948) );
  DFF_X1 \REGISTERS_reg[48][21]  ( .D(n8431), .CK(CLK), .QN(n15949) );
  DFF_X1 \REGISTERS_reg[48][20]  ( .D(n8430), .CK(CLK), .QN(n15950) );
  DFF_X1 \REGISTERS_reg[48][19]  ( .D(n8429), .CK(CLK), .QN(n15951) );
  DFF_X1 \REGISTERS_reg[48][18]  ( .D(n8428), .CK(CLK), .QN(n15952) );
  DFF_X1 \REGISTERS_reg[48][17]  ( .D(n8427), .CK(CLK), .QN(n15953) );
  DFF_X1 \REGISTERS_reg[48][16]  ( .D(n8426), .CK(CLK), .QN(n15954) );
  DFF_X1 \REGISTERS_reg[48][15]  ( .D(n8425), .CK(CLK), .QN(n15955) );
  DFF_X1 \REGISTERS_reg[48][14]  ( .D(n8424), .CK(CLK), .QN(n15956) );
  DFF_X1 \REGISTERS_reg[48][13]  ( .D(n8423), .CK(CLK), .QN(n15957) );
  DFF_X1 \REGISTERS_reg[48][12]  ( .D(n8422), .CK(CLK), .QN(n15958) );
  DFF_X1 \REGISTERS_reg[48][11]  ( .D(n8421), .CK(CLK), .QN(n15959) );
  DFF_X1 \REGISTERS_reg[48][10]  ( .D(n8420), .CK(CLK), .QN(n15960) );
  DFF_X1 \REGISTERS_reg[48][9]  ( .D(n8419), .CK(CLK), .QN(n15961) );
  DFF_X1 \REGISTERS_reg[48][8]  ( .D(n8418), .CK(CLK), .QN(n15962) );
  DFF_X1 \REGISTERS_reg[48][7]  ( .D(n8417), .CK(CLK), .QN(n15963) );
  DFF_X1 \REGISTERS_reg[48][6]  ( .D(n8416), .CK(CLK), .QN(n15964) );
  DFF_X1 \REGISTERS_reg[48][5]  ( .D(n8415), .CK(CLK), .QN(n15965) );
  DFF_X1 \REGISTERS_reg[48][4]  ( .D(n8414), .CK(CLK), .QN(n15966) );
  DFF_X1 \REGISTERS_reg[48][3]  ( .D(n8413), .CK(CLK), .QN(n15967) );
  DFF_X1 \REGISTERS_reg[48][2]  ( .D(n8412), .CK(CLK), .QN(n15968) );
  DFF_X1 \REGISTERS_reg[48][1]  ( .D(n8411), .CK(CLK), .QN(n15969) );
  DFF_X1 \REGISTERS_reg[48][0]  ( .D(n8410), .CK(CLK), .QN(n15970) );
  TINV_X1 U5 ( .I(n1449), .EN(n6659), .ZN(OUT1[31]) );
  TINV_X1 U6 ( .I(n1450), .EN(n6661), .ZN(OUT1[30]) );
  TINV_X1 U7 ( .I(n1451), .EN(n6663), .ZN(OUT1[29]) );
  TINV_X1 U8 ( .I(n1452), .EN(n6665), .ZN(OUT1[28]) );
  TINV_X1 U9 ( .I(n1453), .EN(n6667), .ZN(OUT1[27]) );
  TINV_X1 U10 ( .I(n1454), .EN(n6669), .ZN(OUT1[26]) );
  TINV_X1 U11 ( .I(n1455), .EN(n6671), .ZN(OUT1[25]) );
  TINV_X1 U12 ( .I(n1456), .EN(n6673), .ZN(OUT1[24]) );
  TINV_X1 U13 ( .I(n1457), .EN(n6675), .ZN(OUT1[23]) );
  TINV_X1 U14 ( .I(n1458), .EN(n6677), .ZN(OUT1[22]) );
  TINV_X1 U15 ( .I(n1459), .EN(n6679), .ZN(OUT1[21]) );
  TINV_X1 U16 ( .I(n1460), .EN(n6681), .ZN(OUT1[20]) );
  TINV_X1 U17 ( .I(n1461), .EN(n6683), .ZN(OUT1[19]) );
  TINV_X1 U18 ( .I(n1462), .EN(n6685), .ZN(OUT1[18]) );
  TINV_X1 U19 ( .I(n1463), .EN(n6687), .ZN(OUT1[17]) );
  TINV_X1 U20 ( .I(n1464), .EN(n6689), .ZN(OUT1[16]) );
  TINV_X1 U21 ( .I(n1465), .EN(n6691), .ZN(OUT1[15]) );
  TINV_X1 U22 ( .I(n1466), .EN(n6693), .ZN(OUT1[14]) );
  TINV_X1 U23 ( .I(n1467), .EN(n6695), .ZN(OUT1[13]) );
  TINV_X1 U24 ( .I(n1468), .EN(n6697), .ZN(OUT1[12]) );
  TINV_X1 U25 ( .I(n1469), .EN(n6699), .ZN(OUT1[11]) );
  TINV_X1 U26 ( .I(n1470), .EN(n6701), .ZN(OUT1[10]) );
  TINV_X1 U27 ( .I(n1471), .EN(n6703), .ZN(OUT1[9]) );
  TINV_X1 U28 ( .I(n1472), .EN(n6705), .ZN(OUT1[8]) );
  TINV_X1 U29 ( .I(n1473), .EN(n6707), .ZN(OUT1[7]) );
  TINV_X1 U30 ( .I(n1474), .EN(n6709), .ZN(OUT1[6]) );
  TINV_X1 U31 ( .I(n1475), .EN(n6711), .ZN(OUT1[5]) );
  TINV_X1 U32 ( .I(n1476), .EN(n6713), .ZN(OUT1[4]) );
  TINV_X1 U33 ( .I(n1477), .EN(n6715), .ZN(OUT1[3]) );
  TINV_X1 U34 ( .I(n1478), .EN(n6717), .ZN(OUT1[2]) );
  TINV_X1 U35 ( .I(n1479), .EN(n6719), .ZN(OUT1[1]) );
  TINV_X1 U36 ( .I(n1480), .EN(n6721), .ZN(OUT1[0]) );
  TINV_X1 U37 ( .I(n1481), .EN(n6723), .ZN(OUT2[31]) );
  TINV_X1 U38 ( .I(n1482), .EN(n6725), .ZN(OUT2[30]) );
  TINV_X1 U39 ( .I(n1483), .EN(n6727), .ZN(OUT2[29]) );
  TINV_X1 U40 ( .I(n1484), .EN(n6729), .ZN(OUT2[28]) );
  TINV_X1 U41 ( .I(n1485), .EN(n6731), .ZN(OUT2[27]) );
  TINV_X1 U42 ( .I(n1486), .EN(n6733), .ZN(OUT2[26]) );
  TINV_X1 U43 ( .I(n1487), .EN(n6735), .ZN(OUT2[25]) );
  TINV_X1 U44 ( .I(n1488), .EN(n6737), .ZN(OUT2[24]) );
  TINV_X1 U45 ( .I(n1489), .EN(n6739), .ZN(OUT2[23]) );
  TINV_X1 U46 ( .I(n1490), .EN(n6741), .ZN(OUT2[22]) );
  TINV_X1 U47 ( .I(n1491), .EN(n6743), .ZN(OUT2[21]) );
  TINV_X1 U48 ( .I(n1492), .EN(n6745), .ZN(OUT2[20]) );
  TINV_X1 U49 ( .I(n1493), .EN(n6747), .ZN(OUT2[19]) );
  TINV_X1 U50 ( .I(n1494), .EN(n6749), .ZN(OUT2[18]) );
  TINV_X1 U51 ( .I(n1495), .EN(n6751), .ZN(OUT2[17]) );
  TINV_X1 U52 ( .I(n1496), .EN(n6753), .ZN(OUT2[16]) );
  TINV_X1 U53 ( .I(n1497), .EN(n6755), .ZN(OUT2[15]) );
  TINV_X1 U54 ( .I(n1498), .EN(n6757), .ZN(OUT2[14]) );
  TINV_X1 U55 ( .I(n1499), .EN(n6759), .ZN(OUT2[13]) );
  TINV_X1 U56 ( .I(n1500), .EN(n6761), .ZN(OUT2[12]) );
  TINV_X1 U57 ( .I(n1501), .EN(n6763), .ZN(OUT2[11]) );
  TINV_X1 U58 ( .I(n1502), .EN(n6765), .ZN(OUT2[10]) );
  TINV_X1 U59 ( .I(n1503), .EN(n6767), .ZN(OUT2[9]) );
  TINV_X1 U60 ( .I(n1504), .EN(n6769), .ZN(OUT2[8]) );
  TINV_X1 U61 ( .I(n1505), .EN(n6771), .ZN(OUT2[7]) );
  TINV_X1 U62 ( .I(n1506), .EN(n6773), .ZN(OUT2[6]) );
  TINV_X1 U63 ( .I(n1507), .EN(n6775), .ZN(OUT2[5]) );
  TINV_X1 U64 ( .I(n1508), .EN(n6777), .ZN(OUT2[4]) );
  TINV_X1 U65 ( .I(n1509), .EN(n6779), .ZN(OUT2[3]) );
  TINV_X1 U66 ( .I(n1510), .EN(n6781), .ZN(OUT2[2]) );
  TINV_X1 U67 ( .I(n1511), .EN(n6783), .ZN(OUT2[1]) );
  TINV_X1 U68 ( .I(n1512), .EN(n6785), .ZN(OUT2[0]) );
  NOR4_X2 U3817 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[5]), .A4(
        ADD_RD1[6]), .ZN(n4282) );
  NOR4_X2 U5158 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[5]), .A4(
        ADD_RD2[6]), .ZN(n5679) );
  NOR3_X2 U5252 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(ADD_RD2[0]), .ZN(n5660) );
  XOR2_X1 U7617 ( .A(ADD_WR[6]), .B(ADD_RD1[6]), .Z(n4320) );
  XOR2_X1 U7618 ( .A(ADD_WR[5]), .B(ADD_RD1[5]), .Z(n4319) );
  XOR2_X1 U7619 ( .A(ADD_WR[4]), .B(ADD_RD1[4]), .Z(n4318) );
  XOR2_X1 U7620 ( .A(ADD_WR[3]), .B(ADD_RD1[3]), .Z(n4317) );
  XOR2_X1 U7621 ( .A(ADD_WR[0]), .B(ADD_RD1[0]), .Z(n4321) );
  XOR2_X1 U7622 ( .A(n16071), .B(ADD_RD1[1]), .Z(n4314) );
  XOR2_X1 U7623 ( .A(n16072), .B(ADD_RD1[2]), .Z(n4313) );
  XOR2_X1 U7624 ( .A(ADD_WR[6]), .B(ADD_RD2[6]), .Z(n5752) );
  XOR2_X1 U7625 ( .A(ADD_WR[5]), .B(ADD_RD2[5]), .Z(n5750) );
  XOR2_X1 U7626 ( .A(ADD_WR[4]), .B(ADD_RD2[4]), .Z(n5748) );
  XOR2_X1 U7627 ( .A(ADD_WR[3]), .B(ADD_RD2[3]), .Z(n5746) );
  XOR2_X1 U7628 ( .A(ADD_WR[0]), .B(ADD_RD2[0]), .Z(n5754) );
  XOR2_X1 U7629 ( .A(n16071), .B(ADD_RD2[1]), .Z(n5740) );
  XOR2_X1 U7630 ( .A(n16072), .B(ADD_RD2[2]), .Z(n5738) );
  DFF_X1 \REGISTERS_reg[68][31]  ( .D(n7801), .CK(CLK), .Q(n15430), .QN(n6973)
         );
  DFF_X1 \REGISTERS_reg[68][30]  ( .D(n7800), .CK(CLK), .Q(n15431), .QN(n6972)
         );
  DFF_X1 \REGISTERS_reg[68][29]  ( .D(n7799), .CK(CLK), .Q(n15432), .QN(n6971)
         );
  DFF_X1 \REGISTERS_reg[68][28]  ( .D(n7798), .CK(CLK), .Q(n15433), .QN(n6970)
         );
  DFF_X1 \REGISTERS_reg[68][27]  ( .D(n7797), .CK(CLK), .Q(n15434), .QN(n6969)
         );
  DFF_X1 \REGISTERS_reg[68][26]  ( .D(n7796), .CK(CLK), .Q(n15435), .QN(n6968)
         );
  DFF_X1 \REGISTERS_reg[68][25]  ( .D(n7795), .CK(CLK), .Q(n15436), .QN(n6967)
         );
  DFF_X1 \REGISTERS_reg[68][24]  ( .D(n7794), .CK(CLK), .Q(n15437), .QN(n6966)
         );
  DFF_X1 \REGISTERS_reg[67][31]  ( .D(n7833), .CK(CLK), .Q(n15398), .QN(n7191)
         );
  DFF_X1 \REGISTERS_reg[67][30]  ( .D(n7832), .CK(CLK), .Q(n15399), .QN(n7190)
         );
  DFF_X1 \REGISTERS_reg[67][29]  ( .D(n7831), .CK(CLK), .Q(n15400), .QN(n7189)
         );
  DFF_X1 \REGISTERS_reg[67][28]  ( .D(n7830), .CK(CLK), .Q(n15401), .QN(n7188)
         );
  DFF_X1 \REGISTERS_reg[67][27]  ( .D(n7829), .CK(CLK), .Q(n15402), .QN(n7187)
         );
  DFF_X1 \REGISTERS_reg[67][26]  ( .D(n7828), .CK(CLK), .Q(n15403), .QN(n7186)
         );
  DFF_X1 \REGISTERS_reg[67][25]  ( .D(n7827), .CK(CLK), .Q(n15404), .QN(n7185)
         );
  DFF_X1 \REGISTERS_reg[67][24]  ( .D(n7826), .CK(CLK), .Q(n15405), .QN(n7184)
         );
  DFF_X1 \REGISTERS_reg[63][31]  ( .D(n7961), .CK(CLK), .Q(n15302), .QN(n7223)
         );
  DFF_X1 \REGISTERS_reg[63][30]  ( .D(n7960), .CK(CLK), .Q(n15303), .QN(n7222)
         );
  DFF_X1 \REGISTERS_reg[63][29]  ( .D(n7959), .CK(CLK), .Q(n15304), .QN(n7221)
         );
  DFF_X1 \REGISTERS_reg[63][28]  ( .D(n7958), .CK(CLK), .Q(n15305), .QN(n7220)
         );
  DFF_X1 \REGISTERS_reg[63][27]  ( .D(n7957), .CK(CLK), .Q(n15306), .QN(n7219)
         );
  DFF_X1 \REGISTERS_reg[63][26]  ( .D(n7956), .CK(CLK), .Q(n15307), .QN(n7218)
         );
  DFF_X1 \REGISTERS_reg[63][25]  ( .D(n7955), .CK(CLK), .Q(n15308), .QN(n7217)
         );
  DFF_X1 \REGISTERS_reg[63][24]  ( .D(n7954), .CK(CLK), .Q(n15309), .QN(n7216)
         );
  DFF_X1 \REGISTERS_reg[58][31]  ( .D(n8121), .CK(CLK), .Q(n15174), .QN(n7255)
         );
  DFF_X1 \REGISTERS_reg[58][30]  ( .D(n8120), .CK(CLK), .Q(n15175), .QN(n7254)
         );
  DFF_X1 \REGISTERS_reg[58][29]  ( .D(n8119), .CK(CLK), .Q(n15176), .QN(n7253)
         );
  DFF_X1 \REGISTERS_reg[58][28]  ( .D(n8118), .CK(CLK), .Q(n15177), .QN(n7252)
         );
  DFF_X1 \REGISTERS_reg[58][27]  ( .D(n8117), .CK(CLK), .Q(n15178), .QN(n7251)
         );
  DFF_X1 \REGISTERS_reg[58][26]  ( .D(n8116), .CK(CLK), .Q(n15179), .QN(n7250)
         );
  DFF_X1 \REGISTERS_reg[58][25]  ( .D(n8115), .CK(CLK), .Q(n15180), .QN(n7249)
         );
  DFF_X1 \REGISTERS_reg[58][24]  ( .D(n8114), .CK(CLK), .Q(n15181), .QN(n7248)
         );
  DFF_X1 \REGISTERS_reg[50][31]  ( .D(n8377), .CK(CLK), .Q(n14982), .QN(n6981)
         );
  DFF_X1 \REGISTERS_reg[50][30]  ( .D(n8376), .CK(CLK), .Q(n14983), .QN(n6980)
         );
  DFF_X1 \REGISTERS_reg[50][29]  ( .D(n8375), .CK(CLK), .Q(n14984), .QN(n6979)
         );
  DFF_X1 \REGISTERS_reg[50][28]  ( .D(n8374), .CK(CLK), .Q(n14985), .QN(n6978)
         );
  DFF_X1 \REGISTERS_reg[50][27]  ( .D(n8373), .CK(CLK), .Q(n14986), .QN(n6977)
         );
  DFF_X1 \REGISTERS_reg[50][26]  ( .D(n8372), .CK(CLK), .Q(n14987), .QN(n6976)
         );
  DFF_X1 \REGISTERS_reg[50][25]  ( .D(n8371), .CK(CLK), .Q(n14988), .QN(n6975)
         );
  DFF_X1 \REGISTERS_reg[50][24]  ( .D(n8370), .CK(CLK), .Q(n14989), .QN(n6974)
         );
  DFF_X1 \REGISTERS_reg[49][31]  ( .D(n8409), .CK(CLK), .Q(n15634), .QN(n969)
         );
  DFF_X1 \REGISTERS_reg[49][30]  ( .D(n8408), .CK(CLK), .Q(n15635), .QN(n970)
         );
  DFF_X1 \REGISTERS_reg[49][29]  ( .D(n8407), .CK(CLK), .Q(n15636), .QN(n971)
         );
  DFF_X1 \REGISTERS_reg[49][28]  ( .D(n8406), .CK(CLK), .Q(n15637), .QN(n972)
         );
  DFF_X1 \REGISTERS_reg[49][27]  ( .D(n8405), .CK(CLK), .Q(n15638), .QN(n973)
         );
  DFF_X1 \REGISTERS_reg[49][26]  ( .D(n8404), .CK(CLK), .Q(n15639), .QN(n974)
         );
  DFF_X1 \REGISTERS_reg[49][25]  ( .D(n8403), .CK(CLK), .Q(n15640), .QN(n975)
         );
  DFF_X1 \REGISTERS_reg[49][24]  ( .D(n8402), .CK(CLK), .Q(n15641), .QN(n976)
         );
  DFF_X1 \REGISTERS_reg[45][31]  ( .D(n8537), .CK(CLK), .Q(n14948), .QN(n7257)
         );
  DFF_X1 \REGISTERS_reg[45][30]  ( .D(n8536), .CK(CLK), .Q(n15613), .QN(n622)
         );
  DFF_X1 \REGISTERS_reg[45][29]  ( .D(n8535), .CK(CLK), .Q(n15614), .QN(n625)
         );
  DFF_X1 \REGISTERS_reg[45][28]  ( .D(n8534), .CK(CLK), .Q(n15615), .QN(n628)
         );
  DFF_X1 \REGISTERS_reg[45][27]  ( .D(n8533), .CK(CLK), .Q(n15616), .QN(n631)
         );
  DFF_X1 \REGISTERS_reg[45][26]  ( .D(n8532), .CK(CLK), .Q(n15617), .QN(n634)
         );
  DFF_X1 \REGISTERS_reg[45][25]  ( .D(n8531), .CK(CLK), .Q(n15618), .QN(n637)
         );
  DFF_X1 \REGISTERS_reg[45][24]  ( .D(n8530), .CK(CLK), .Q(n15619), .QN(n640)
         );
  DFF_X1 \REGISTERS_reg[40][31]  ( .D(n8697), .CK(CLK), .Q(n15558), .QN(n937)
         );
  DFF_X1 \REGISTERS_reg[40][30]  ( .D(n8696), .CK(CLK), .Q(n15559), .QN(n938)
         );
  DFF_X1 \REGISTERS_reg[40][29]  ( .D(n8695), .CK(CLK), .Q(n15560), .QN(n939)
         );
  DFF_X1 \REGISTERS_reg[40][28]  ( .D(n8694), .CK(CLK), .Q(n15561), .QN(n940)
         );
  DFF_X1 \REGISTERS_reg[40][27]  ( .D(n8693), .CK(CLK), .Q(n15562), .QN(n941)
         );
  DFF_X1 \REGISTERS_reg[40][26]  ( .D(n8692), .CK(CLK), .Q(n15563), .QN(n942)
         );
  DFF_X1 \REGISTERS_reg[40][25]  ( .D(n8691), .CK(CLK), .Q(n15564), .QN(n943)
         );
  DFF_X1 \REGISTERS_reg[40][24]  ( .D(n8690), .CK(CLK), .Q(n15565), .QN(n944)
         );
  DFF_X1 \REGISTERS_reg[32][31]  ( .D(n8953), .CK(CLK), .Q(n14660), .QN(n6989)
         );
  DFF_X1 \REGISTERS_reg[32][30]  ( .D(n8952), .CK(CLK), .Q(n14661), .QN(n6988)
         );
  DFF_X1 \REGISTERS_reg[32][29]  ( .D(n8951), .CK(CLK), .Q(n14662), .QN(n6987)
         );
  DFF_X1 \REGISTERS_reg[32][28]  ( .D(n8950), .CK(CLK), .Q(n14663), .QN(n6986)
         );
  DFF_X1 \REGISTERS_reg[32][27]  ( .D(n8949), .CK(CLK), .Q(n14664), .QN(n6985)
         );
  DFF_X1 \REGISTERS_reg[32][26]  ( .D(n8948), .CK(CLK), .Q(n14665), .QN(n6984)
         );
  DFF_X1 \REGISTERS_reg[32][25]  ( .D(n8947), .CK(CLK), .Q(n14666), .QN(n6983)
         );
  DFF_X1 \REGISTERS_reg[32][24]  ( .D(n8946), .CK(CLK), .Q(n14667), .QN(n6982)
         );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n8985), .CK(CLK), .Q(n15566), .QN(n905)
         );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n8984), .CK(CLK), .Q(n15567), .QN(n906)
         );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n8983), .CK(CLK), .Q(n15568), .QN(n907)
         );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n8982), .CK(CLK), .Q(n15569), .QN(n908)
         );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n8981), .CK(CLK), .Q(n15570), .QN(n909)
         );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n8980), .CK(CLK), .Q(n15571), .QN(n910)
         );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n8979), .CK(CLK), .Q(n15572), .QN(n911)
         );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n8978), .CK(CLK), .Q(n15573), .QN(n912)
         );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n9017), .CK(CLK), .Q(n15574), .QN(n5693)
         );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n9016), .CK(CLK), .Q(n15575), .QN(n5683)
         );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n9015), .CK(CLK), .Q(n15576), .QN(n5673)
         );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n9014), .CK(CLK), .Q(n15577), .QN(n5663)
         );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n9013), .CK(CLK), .Q(n15578), .QN(n5653)
         );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n9012), .CK(CLK), .Q(n15579), .QN(n5643)
         );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n9011), .CK(CLK), .Q(n15580), .QN(n5633)
         );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n9010), .CK(CLK), .Q(n15581), .QN(n5623)
         );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n9049), .CK(CLK), .Q(n15790), .QN(n5692)
         );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n9048), .CK(CLK), .Q(n15791), .QN(n5682)
         );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n9047), .CK(CLK), .Q(n15792), .QN(n5672)
         );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n9046), .CK(CLK), .Q(n15793), .QN(n5662)
         );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n9045), .CK(CLK), .Q(n15794), .QN(n5652)
         );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n9044), .CK(CLK), .Q(n15795), .QN(n5642)
         );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n9043), .CK(CLK), .Q(n15796), .QN(n5632)
         );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n9042), .CK(CLK), .Q(n15797), .QN(n5622)
         );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n9241), .CK(CLK), .Q(n14461), .QN(n6997)
         );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n9240), .CK(CLK), .Q(n14462), .QN(n6996)
         );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n9239), .CK(CLK), .Q(n14463), .QN(n6995)
         );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n9238), .CK(CLK), .Q(n14464), .QN(n6994)
         );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n9237), .CK(CLK), .Q(n14465), .QN(n6993)
         );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n9236), .CK(CLK), .Q(n14466), .QN(n6992)
         );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n9235), .CK(CLK), .Q(n14467), .QN(n6991)
         );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n9234), .CK(CLK), .Q(n14468), .QN(n6990)
         );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n9273), .CK(CLK), .Q(n15582), .QN(n873)
         );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n9272), .CK(CLK), .Q(n15583), .QN(n874)
         );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n9271), .CK(CLK), .Q(n15584), .QN(n875)
         );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n9270), .CK(CLK), .Q(n15585), .QN(n876)
         );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n9269), .CK(CLK), .Q(n15586), .QN(n877)
         );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n9268), .CK(CLK), .Q(n15587), .QN(n878)
         );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n9267), .CK(CLK), .Q(n15588), .QN(n879)
         );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n9266), .CK(CLK), .Q(n15589), .QN(n880)
         );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n9337), .CK(CLK), .Q(n15862), .QN(n5824)
         );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n9336), .CK(CLK), .Q(n15863), .QN(n5820)
         );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n9335), .CK(CLK), .Q(n15864), .QN(n5816)
         );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n9334), .CK(CLK), .Q(n15865), .QN(n5812)
         );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n9333), .CK(CLK), .Q(n15866), .QN(n5808)
         );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n9332), .CK(CLK), .Q(n15867), .QN(n5804)
         );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n9331), .CK(CLK), .Q(n15868), .QN(n5800)
         );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n9330), .CK(CLK), .Q(n15869), .QN(n5796)
         );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n9529), .CK(CLK), .Q(n14248), .QN(n7013)
         );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n9528), .CK(CLK), .Q(n14249), .QN(n7012)
         );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n9527), .CK(CLK), .Q(n14250), .QN(n7011)
         );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n9526), .CK(CLK), .Q(n14251), .QN(n7010)
         );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n9525), .CK(CLK), .Q(n14252), .QN(n7009)
         );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n9524), .CK(CLK), .Q(n14253), .QN(n7008)
         );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n9523), .CK(CLK), .Q(n14254), .QN(n7007)
         );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n9522), .CK(CLK), .Q(n14255), .QN(n7006)
         );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n9561), .CK(CLK), .Q(n15590), .QN(n841)
         );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n9560), .CK(CLK), .Q(n15591), .QN(n842)
         );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n9559), .CK(CLK), .Q(n15592), .QN(n843)
         );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n9558), .CK(CLK), .Q(n15593), .QN(n844)
         );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n9557), .CK(CLK), .Q(n15594), .QN(n845)
         );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n9556), .CK(CLK), .Q(n15595), .QN(n846)
         );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n9555), .CK(CLK), .Q(n15596), .QN(n847)
         );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n9554), .CK(CLK), .Q(n15597), .QN(n848)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n9817), .CK(CLK), .Q(n14076), .QN(n7021)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n9816), .CK(CLK), .Q(n14077), .QN(n7020)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n9815), .CK(CLK), .Q(n14078), .QN(n7019)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n9814), .CK(CLK), .Q(n14079), .QN(n7018)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n9813), .CK(CLK), .Q(n14080), .QN(n7017)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n9812), .CK(CLK), .Q(n14081), .QN(n7016)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n9811), .CK(CLK), .Q(n14082), .QN(n7015)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n9810), .CK(CLK), .Q(n14083), .QN(n7014)
         );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n9849), .CK(CLK), .Q(n15598), .QN(n809)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n9848), .CK(CLK), .Q(n15599), .QN(n810)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n9847), .CK(CLK), .Q(n15600), .QN(n811)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n9846), .CK(CLK), .Q(n15601), .QN(n812)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n9845), .CK(CLK), .Q(n15602), .QN(n813)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n9844), .CK(CLK), .Q(n15603), .QN(n814)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n9843), .CK(CLK), .Q(n15604), .QN(n815)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n9842), .CK(CLK), .Q(n15605), .QN(n816)
         );
  DFF_X1 \REGISTERS_reg[39][30]  ( .D(n8728), .CK(CLK), .Q(n15620), .QN(n5819)
         );
  DFF_X1 \REGISTERS_reg[39][29]  ( .D(n8727), .CK(CLK), .Q(n15621), .QN(n5815)
         );
  DFF_X1 \REGISTERS_reg[39][28]  ( .D(n8726), .CK(CLK), .Q(n15622), .QN(n5811)
         );
  DFF_X1 \REGISTERS_reg[39][27]  ( .D(n8725), .CK(CLK), .Q(n15623), .QN(n5807)
         );
  DFF_X1 \REGISTERS_reg[39][26]  ( .D(n8724), .CK(CLK), .Q(n15624), .QN(n5803)
         );
  DFF_X1 \REGISTERS_reg[39][25]  ( .D(n8723), .CK(CLK), .Q(n15625), .QN(n5799)
         );
  DFF_X1 \REGISTERS_reg[39][24]  ( .D(n8722), .CK(CLK), .Q(n15626), .QN(n5795)
         );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n9303), .CK(CLK), .Q(n15627), .QN(n5817)
         );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n9302), .CK(CLK), .Q(n15628), .QN(n5813)
         );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n9301), .CK(CLK), .Q(n15629), .QN(n5809)
         );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n9300), .CK(CLK), .Q(n15630), .QN(n5805)
         );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n9299), .CK(CLK), .Q(n15631), .QN(n5801)
         );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n9298), .CK(CLK), .Q(n15632), .QN(n5797)
         );
  DFF_X1 \REGISTERS_reg[68][23]  ( .D(n7793), .CK(CLK), .Q(n15438), .QN(n6965)
         );
  DFF_X1 \REGISTERS_reg[68][22]  ( .D(n7792), .CK(CLK), .Q(n15439), .QN(n6964)
         );
  DFF_X1 \REGISTERS_reg[68][21]  ( .D(n7791), .CK(CLK), .Q(n15440), .QN(n6963)
         );
  DFF_X1 \REGISTERS_reg[68][20]  ( .D(n7790), .CK(CLK), .Q(n15441), .QN(n6962)
         );
  DFF_X1 \REGISTERS_reg[68][19]  ( .D(n7789), .CK(CLK), .Q(n15442), .QN(n6961)
         );
  DFF_X1 \REGISTERS_reg[68][18]  ( .D(n7788), .CK(CLK), .Q(n15443), .QN(n6960)
         );
  DFF_X1 \REGISTERS_reg[68][17]  ( .D(n7787), .CK(CLK), .Q(n15444), .QN(n6959)
         );
  DFF_X1 \REGISTERS_reg[68][16]  ( .D(n7786), .CK(CLK), .Q(n15445), .QN(n6958)
         );
  DFF_X1 \REGISTERS_reg[68][15]  ( .D(n7785), .CK(CLK), .Q(n15446), .QN(n6957)
         );
  DFF_X1 \REGISTERS_reg[68][14]  ( .D(n7784), .CK(CLK), .Q(n15447), .QN(n6956)
         );
  DFF_X1 \REGISTERS_reg[68][13]  ( .D(n7783), .CK(CLK), .Q(n15448), .QN(n6955)
         );
  DFF_X1 \REGISTERS_reg[68][12]  ( .D(n7782), .CK(CLK), .Q(n15449), .QN(n6954)
         );
  DFF_X1 \REGISTERS_reg[68][11]  ( .D(n7781), .CK(CLK), .Q(n15450), .QN(n6953)
         );
  DFF_X1 \REGISTERS_reg[68][10]  ( .D(n7780), .CK(CLK), .Q(n15451), .QN(n6952)
         );
  DFF_X1 \REGISTERS_reg[68][9]  ( .D(n7779), .CK(CLK), .Q(n15452), .QN(n6951)
         );
  DFF_X1 \REGISTERS_reg[68][8]  ( .D(n7778), .CK(CLK), .Q(n15453), .QN(n6950)
         );
  DFF_X1 \REGISTERS_reg[68][7]  ( .D(n7777), .CK(CLK), .Q(n15454), .QN(n6949)
         );
  DFF_X1 \REGISTERS_reg[68][6]  ( .D(n7776), .CK(CLK), .Q(n15455), .QN(n6948)
         );
  DFF_X1 \REGISTERS_reg[68][5]  ( .D(n7775), .CK(CLK), .Q(n15456), .QN(n6947)
         );
  DFF_X1 \REGISTERS_reg[68][4]  ( .D(n7774), .CK(CLK), .Q(n15457), .QN(n6946)
         );
  DFF_X1 \REGISTERS_reg[68][3]  ( .D(n7773), .CK(CLK), .Q(n15458), .QN(n6945)
         );
  DFF_X1 \REGISTERS_reg[68][2]  ( .D(n7772), .CK(CLK), .Q(n15459), .QN(n6944)
         );
  DFF_X1 \REGISTERS_reg[68][1]  ( .D(n7771), .CK(CLK), .Q(n15460), .QN(n6943)
         );
  DFF_X1 \REGISTERS_reg[68][0]  ( .D(n7770), .CK(CLK), .Q(n15461), .QN(n6942)
         );
  DFF_X1 \REGISTERS_reg[67][23]  ( .D(n7825), .CK(CLK), .Q(n15406), .QN(n7183)
         );
  DFF_X1 \REGISTERS_reg[67][22]  ( .D(n7824), .CK(CLK), .Q(n15407), .QN(n7182)
         );
  DFF_X1 \REGISTERS_reg[67][21]  ( .D(n7823), .CK(CLK), .Q(n15408), .QN(n7181)
         );
  DFF_X1 \REGISTERS_reg[67][20]  ( .D(n7822), .CK(CLK), .Q(n15409), .QN(n7180)
         );
  DFF_X1 \REGISTERS_reg[67][19]  ( .D(n7821), .CK(CLK), .Q(n15410), .QN(n7179)
         );
  DFF_X1 \REGISTERS_reg[67][18]  ( .D(n7820), .CK(CLK), .Q(n15411), .QN(n7178)
         );
  DFF_X1 \REGISTERS_reg[67][17]  ( .D(n7819), .CK(CLK), .Q(n15412), .QN(n7177)
         );
  DFF_X1 \REGISTERS_reg[67][16]  ( .D(n7818), .CK(CLK), .Q(n15413), .QN(n7176)
         );
  DFF_X1 \REGISTERS_reg[67][15]  ( .D(n7817), .CK(CLK), .Q(n15414), .QN(n7175)
         );
  DFF_X1 \REGISTERS_reg[67][14]  ( .D(n7816), .CK(CLK), .Q(n15415), .QN(n7174)
         );
  DFF_X1 \REGISTERS_reg[67][13]  ( .D(n7815), .CK(CLK), .Q(n15416), .QN(n7173)
         );
  DFF_X1 \REGISTERS_reg[67][12]  ( .D(n7814), .CK(CLK), .Q(n15417), .QN(n7172)
         );
  DFF_X1 \REGISTERS_reg[67][11]  ( .D(n7813), .CK(CLK), .Q(n15418), .QN(n7171)
         );
  DFF_X1 \REGISTERS_reg[67][10]  ( .D(n7812), .CK(CLK), .Q(n15419), .QN(n7170)
         );
  DFF_X1 \REGISTERS_reg[67][9]  ( .D(n7811), .CK(CLK), .Q(n15420), .QN(n7169)
         );
  DFF_X1 \REGISTERS_reg[67][8]  ( .D(n7810), .CK(CLK), .Q(n15421), .QN(n7168)
         );
  DFF_X1 \REGISTERS_reg[67][7]  ( .D(n7809), .CK(CLK), .Q(n15422), .QN(n7167)
         );
  DFF_X1 \REGISTERS_reg[67][6]  ( .D(n7808), .CK(CLK), .Q(n15423), .QN(n7166)
         );
  DFF_X1 \REGISTERS_reg[67][5]  ( .D(n7807), .CK(CLK), .Q(n15424), .QN(n7165)
         );
  DFF_X1 \REGISTERS_reg[67][4]  ( .D(n7806), .CK(CLK), .Q(n15425), .QN(n7164)
         );
  DFF_X1 \REGISTERS_reg[67][3]  ( .D(n7805), .CK(CLK), .Q(n15426), .QN(n7163)
         );
  DFF_X1 \REGISTERS_reg[67][2]  ( .D(n7804), .CK(CLK), .Q(n15427), .QN(n7162)
         );
  DFF_X1 \REGISTERS_reg[67][1]  ( .D(n7803), .CK(CLK), .Q(n15428), .QN(n7161)
         );
  DFF_X1 \REGISTERS_reg[67][0]  ( .D(n7802), .CK(CLK), .Q(n15429), .QN(n7160)
         );
  DFF_X1 \REGISTERS_reg[63][23]  ( .D(n7953), .CK(CLK), .Q(n15310), .QN(n7215)
         );
  DFF_X1 \REGISTERS_reg[63][22]  ( .D(n7952), .CK(CLK), .Q(n15311), .QN(n7214)
         );
  DFF_X1 \REGISTERS_reg[63][21]  ( .D(n7951), .CK(CLK), .Q(n15312), .QN(n7213)
         );
  DFF_X1 \REGISTERS_reg[63][20]  ( .D(n7950), .CK(CLK), .Q(n15313), .QN(n7212)
         );
  DFF_X1 \REGISTERS_reg[63][19]  ( .D(n7949), .CK(CLK), .Q(n15314), .QN(n7211)
         );
  DFF_X1 \REGISTERS_reg[63][18]  ( .D(n7948), .CK(CLK), .Q(n15315), .QN(n7210)
         );
  DFF_X1 \REGISTERS_reg[63][17]  ( .D(n7947), .CK(CLK), .Q(n15316), .QN(n7209)
         );
  DFF_X1 \REGISTERS_reg[63][16]  ( .D(n7946), .CK(CLK), .Q(n15317), .QN(n7208)
         );
  DFF_X1 \REGISTERS_reg[63][15]  ( .D(n7945), .CK(CLK), .Q(n15318), .QN(n7207)
         );
  DFF_X1 \REGISTERS_reg[63][14]  ( .D(n7944), .CK(CLK), .Q(n15319), .QN(n7206)
         );
  DFF_X1 \REGISTERS_reg[63][13]  ( .D(n7943), .CK(CLK), .Q(n15320), .QN(n7205)
         );
  DFF_X1 \REGISTERS_reg[63][12]  ( .D(n7942), .CK(CLK), .Q(n15321), .QN(n7204)
         );
  DFF_X1 \REGISTERS_reg[63][11]  ( .D(n7941), .CK(CLK), .Q(n15322), .QN(n7203)
         );
  DFF_X1 \REGISTERS_reg[63][10]  ( .D(n7940), .CK(CLK), .Q(n15323), .QN(n7202)
         );
  DFF_X1 \REGISTERS_reg[63][9]  ( .D(n7939), .CK(CLK), .Q(n15324), .QN(n7201)
         );
  DFF_X1 \REGISTERS_reg[63][8]  ( .D(n7938), .CK(CLK), .Q(n15325), .QN(n7200)
         );
  DFF_X1 \REGISTERS_reg[63][7]  ( .D(n7937), .CK(CLK), .Q(n15326), .QN(n7199)
         );
  DFF_X1 \REGISTERS_reg[63][6]  ( .D(n7936), .CK(CLK), .Q(n15327), .QN(n7198)
         );
  DFF_X1 \REGISTERS_reg[63][5]  ( .D(n7935), .CK(CLK), .Q(n15328), .QN(n7197)
         );
  DFF_X1 \REGISTERS_reg[63][4]  ( .D(n7934), .CK(CLK), .Q(n15329), .QN(n7196)
         );
  DFF_X1 \REGISTERS_reg[63][3]  ( .D(n7933), .CK(CLK), .Q(n15330), .QN(n7195)
         );
  DFF_X1 \REGISTERS_reg[63][2]  ( .D(n7932), .CK(CLK), .Q(n15331), .QN(n7194)
         );
  DFF_X1 \REGISTERS_reg[63][1]  ( .D(n7931), .CK(CLK), .Q(n15332), .QN(n7193)
         );
  DFF_X1 \REGISTERS_reg[63][0]  ( .D(n7930), .CK(CLK), .Q(n15333), .QN(n7192)
         );
  DFF_X1 \REGISTERS_reg[58][23]  ( .D(n8113), .CK(CLK), .Q(n15182), .QN(n7247)
         );
  DFF_X1 \REGISTERS_reg[58][22]  ( .D(n8112), .CK(CLK), .Q(n15183), .QN(n7246)
         );
  DFF_X1 \REGISTERS_reg[58][21]  ( .D(n8111), .CK(CLK), .Q(n15184), .QN(n7245)
         );
  DFF_X1 \REGISTERS_reg[58][20]  ( .D(n8110), .CK(CLK), .Q(n15185), .QN(n7244)
         );
  DFF_X1 \REGISTERS_reg[58][19]  ( .D(n8109), .CK(CLK), .Q(n15186), .QN(n7243)
         );
  DFF_X1 \REGISTERS_reg[58][18]  ( .D(n8108), .CK(CLK), .Q(n15187), .QN(n7242)
         );
  DFF_X1 \REGISTERS_reg[58][17]  ( .D(n8107), .CK(CLK), .Q(n15188), .QN(n7241)
         );
  DFF_X1 \REGISTERS_reg[58][16]  ( .D(n8106), .CK(CLK), .Q(n15189), .QN(n7240)
         );
  DFF_X1 \REGISTERS_reg[58][15]  ( .D(n8105), .CK(CLK), .Q(n15190), .QN(n7239)
         );
  DFF_X1 \REGISTERS_reg[58][14]  ( .D(n8104), .CK(CLK), .Q(n15191), .QN(n7238)
         );
  DFF_X1 \REGISTERS_reg[58][13]  ( .D(n8103), .CK(CLK), .Q(n15192), .QN(n7237)
         );
  DFF_X1 \REGISTERS_reg[58][12]  ( .D(n8102), .CK(CLK), .Q(n15193), .QN(n7236)
         );
  DFF_X1 \REGISTERS_reg[58][11]  ( .D(n8101), .CK(CLK), .Q(n15194), .QN(n7235)
         );
  DFF_X1 \REGISTERS_reg[58][10]  ( .D(n8100), .CK(CLK), .Q(n15195), .QN(n7234)
         );
  DFF_X1 \REGISTERS_reg[58][9]  ( .D(n8099), .CK(CLK), .Q(n15196), .QN(n7233)
         );
  DFF_X1 \REGISTERS_reg[58][8]  ( .D(n8098), .CK(CLK), .Q(n15197), .QN(n7232)
         );
  DFF_X1 \REGISTERS_reg[58][7]  ( .D(n8097), .CK(CLK), .Q(n15198), .QN(n7231)
         );
  DFF_X1 \REGISTERS_reg[58][6]  ( .D(n8096), .CK(CLK), .Q(n15199), .QN(n7230)
         );
  DFF_X1 \REGISTERS_reg[58][5]  ( .D(n8095), .CK(CLK), .Q(n15200), .QN(n7229)
         );
  DFF_X1 \REGISTERS_reg[58][4]  ( .D(n8094), .CK(CLK), .Q(n15201), .QN(n7228)
         );
  DFF_X1 \REGISTERS_reg[58][3]  ( .D(n8093), .CK(CLK), .Q(n15202), .QN(n7227)
         );
  DFF_X1 \REGISTERS_reg[58][2]  ( .D(n8092), .CK(CLK), .Q(n15203), .QN(n7226)
         );
  DFF_X1 \REGISTERS_reg[58][1]  ( .D(n8091), .CK(CLK), .Q(n15204), .QN(n7225)
         );
  DFF_X1 \REGISTERS_reg[58][0]  ( .D(n8090), .CK(CLK), .Q(n15205), .QN(n7224)
         );
  DFF_X1 \REGISTERS_reg[50][23]  ( .D(n8369), .CK(CLK), .Q(n14990), .QN(n7045)
         );
  DFF_X1 \REGISTERS_reg[50][22]  ( .D(n8368), .CK(CLK), .Q(n14991), .QN(n7044)
         );
  DFF_X1 \REGISTERS_reg[50][21]  ( .D(n8367), .CK(CLK), .Q(n14992), .QN(n7043)
         );
  DFF_X1 \REGISTERS_reg[50][20]  ( .D(n8366), .CK(CLK), .Q(n14993), .QN(n7042)
         );
  DFF_X1 \REGISTERS_reg[50][19]  ( .D(n8365), .CK(CLK), .Q(n14994), .QN(n7041)
         );
  DFF_X1 \REGISTERS_reg[50][18]  ( .D(n8364), .CK(CLK), .Q(n14995), .QN(n7040)
         );
  DFF_X1 \REGISTERS_reg[50][17]  ( .D(n8363), .CK(CLK), .Q(n14996), .QN(n7039)
         );
  DFF_X1 \REGISTERS_reg[50][16]  ( .D(n8362), .CK(CLK), .Q(n14997), .QN(n7038)
         );
  DFF_X1 \REGISTERS_reg[50][15]  ( .D(n8361), .CK(CLK), .Q(n14998), .QN(n7037)
         );
  DFF_X1 \REGISTERS_reg[50][14]  ( .D(n8360), .CK(CLK), .Q(n14999), .QN(n7036)
         );
  DFF_X1 \REGISTERS_reg[50][13]  ( .D(n8359), .CK(CLK), .Q(n15000), .QN(n7035)
         );
  DFF_X1 \REGISTERS_reg[50][12]  ( .D(n8358), .CK(CLK), .Q(n15001), .QN(n7034)
         );
  DFF_X1 \REGISTERS_reg[50][11]  ( .D(n8357), .CK(CLK), .Q(n15002), .QN(n7033)
         );
  DFF_X1 \REGISTERS_reg[50][10]  ( .D(n8356), .CK(CLK), .Q(n15003), .QN(n7032)
         );
  DFF_X1 \REGISTERS_reg[50][9]  ( .D(n8355), .CK(CLK), .Q(n15004), .QN(n7031)
         );
  DFF_X1 \REGISTERS_reg[50][8]  ( .D(n8354), .CK(CLK), .Q(n15005), .QN(n7030)
         );
  DFF_X1 \REGISTERS_reg[50][7]  ( .D(n8353), .CK(CLK), .Q(n15006), .QN(n7029)
         );
  DFF_X1 \REGISTERS_reg[50][6]  ( .D(n8352), .CK(CLK), .Q(n15007), .QN(n7028)
         );
  DFF_X1 \REGISTERS_reg[50][5]  ( .D(n8351), .CK(CLK), .Q(n15008), .QN(n7027)
         );
  DFF_X1 \REGISTERS_reg[50][4]  ( .D(n8350), .CK(CLK), .Q(n15009), .QN(n7026)
         );
  DFF_X1 \REGISTERS_reg[50][3]  ( .D(n8349), .CK(CLK), .Q(n15010), .QN(n7025)
         );
  DFF_X1 \REGISTERS_reg[50][2]  ( .D(n8348), .CK(CLK), .Q(n15011), .QN(n7024)
         );
  DFF_X1 \REGISTERS_reg[50][1]  ( .D(n8347), .CK(CLK), .Q(n15012), .QN(n7023)
         );
  DFF_X1 \REGISTERS_reg[50][0]  ( .D(n8346), .CK(CLK), .Q(n15013), .QN(n7022)
         );
  DFF_X1 \REGISTERS_reg[49][23]  ( .D(n8401), .CK(CLK), .Q(n15642), .QN(n977)
         );
  DFF_X1 \REGISTERS_reg[49][22]  ( .D(n8400), .CK(CLK), .Q(n15643), .QN(n978)
         );
  DFF_X1 \REGISTERS_reg[49][21]  ( .D(n8399), .CK(CLK), .Q(n15644), .QN(n979)
         );
  DFF_X1 \REGISTERS_reg[49][20]  ( .D(n8398), .CK(CLK), .Q(n15645), .QN(n980)
         );
  DFF_X1 \REGISTERS_reg[49][19]  ( .D(n8397), .CK(CLK), .Q(n15646), .QN(n981)
         );
  DFF_X1 \REGISTERS_reg[49][18]  ( .D(n8396), .CK(CLK), .Q(n15647), .QN(n982)
         );
  DFF_X1 \REGISTERS_reg[49][17]  ( .D(n8395), .CK(CLK), .Q(n15648), .QN(n983)
         );
  DFF_X1 \REGISTERS_reg[49][16]  ( .D(n8394), .CK(CLK), .Q(n15649), .QN(n984)
         );
  DFF_X1 \REGISTERS_reg[49][15]  ( .D(n8393), .CK(CLK), .Q(n15650), .QN(n985)
         );
  DFF_X1 \REGISTERS_reg[49][14]  ( .D(n8392), .CK(CLK), .Q(n15651), .QN(n986)
         );
  DFF_X1 \REGISTERS_reg[49][13]  ( .D(n8391), .CK(CLK), .Q(n15652), .QN(n987)
         );
  DFF_X1 \REGISTERS_reg[49][12]  ( .D(n8390), .CK(CLK), .Q(n15653), .QN(n988)
         );
  DFF_X1 \REGISTERS_reg[49][11]  ( .D(n8389), .CK(CLK), .Q(n15654), .QN(n989)
         );
  DFF_X1 \REGISTERS_reg[49][10]  ( .D(n8388), .CK(CLK), .Q(n15655), .QN(n990)
         );
  DFF_X1 \REGISTERS_reg[49][9]  ( .D(n8387), .CK(CLK), .Q(n15656), .QN(n991)
         );
  DFF_X1 \REGISTERS_reg[49][8]  ( .D(n8386), .CK(CLK), .Q(n15657), .QN(n992)
         );
  DFF_X1 \REGISTERS_reg[49][7]  ( .D(n8385), .CK(CLK), .Q(n15606), .QN(n993)
         );
  DFF_X1 \REGISTERS_reg[49][6]  ( .D(n8384), .CK(CLK), .Q(n15607), .QN(n994)
         );
  DFF_X1 \REGISTERS_reg[49][5]  ( .D(n8383), .CK(CLK), .Q(n15608), .QN(n995)
         );
  DFF_X1 \REGISTERS_reg[49][4]  ( .D(n8382), .CK(CLK), .Q(n15609), .QN(n996)
         );
  DFF_X1 \REGISTERS_reg[49][3]  ( .D(n8381), .CK(CLK), .Q(n15610), .QN(n997)
         );
  DFF_X1 \REGISTERS_reg[49][2]  ( .D(n8380), .CK(CLK), .Q(n15611), .QN(n998)
         );
  DFF_X1 \REGISTERS_reg[49][1]  ( .D(n8379), .CK(CLK), .Q(n15612), .QN(n999)
         );
  DFF_X1 \REGISTERS_reg[49][0]  ( .D(n8378), .CK(CLK), .Q(n14981), .QN(n7256)
         );
  DFF_X1 \REGISTERS_reg[45][23]  ( .D(n8529), .CK(CLK), .Q(n15658), .QN(n643)
         );
  DFF_X1 \REGISTERS_reg[45][22]  ( .D(n8528), .CK(CLK), .Q(n15659), .QN(n646)
         );
  DFF_X1 \REGISTERS_reg[45][21]  ( .D(n8527), .CK(CLK), .Q(n15660), .QN(n649)
         );
  DFF_X1 \REGISTERS_reg[45][20]  ( .D(n8526), .CK(CLK), .Q(n15661), .QN(n652)
         );
  DFF_X1 \REGISTERS_reg[45][19]  ( .D(n8525), .CK(CLK), .Q(n15662), .QN(n655)
         );
  DFF_X1 \REGISTERS_reg[45][18]  ( .D(n8524), .CK(CLK), .Q(n15663), .QN(n658)
         );
  DFF_X1 \REGISTERS_reg[45][17]  ( .D(n8523), .CK(CLK), .Q(n15664), .QN(n661)
         );
  DFF_X1 \REGISTERS_reg[45][16]  ( .D(n8522), .CK(CLK), .Q(n15665), .QN(n664)
         );
  DFF_X1 \REGISTERS_reg[45][15]  ( .D(n8521), .CK(CLK), .Q(n15666), .QN(n667)
         );
  DFF_X1 \REGISTERS_reg[45][14]  ( .D(n8520), .CK(CLK), .Q(n15667), .QN(n670)
         );
  DFF_X1 \REGISTERS_reg[45][13]  ( .D(n8519), .CK(CLK), .Q(n15668), .QN(n673)
         );
  DFF_X1 \REGISTERS_reg[45][12]  ( .D(n8518), .CK(CLK), .Q(n15669), .QN(n676)
         );
  DFF_X1 \REGISTERS_reg[45][11]  ( .D(n8517), .CK(CLK), .Q(n15670), .QN(n679)
         );
  DFF_X1 \REGISTERS_reg[45][10]  ( .D(n8516), .CK(CLK), .Q(n15671), .QN(n682)
         );
  DFF_X1 \REGISTERS_reg[45][9]  ( .D(n8515), .CK(CLK), .Q(n15672), .QN(n685)
         );
  DFF_X1 \REGISTERS_reg[45][8]  ( .D(n8514), .CK(CLK), .Q(n15673), .QN(n688)
         );
  DFF_X1 \REGISTERS_reg[45][7]  ( .D(n8513), .CK(CLK), .Q(n15674), .QN(n691)
         );
  DFF_X1 \REGISTERS_reg[45][6]  ( .D(n8512), .CK(CLK), .Q(n15675), .QN(n694)
         );
  DFF_X1 \REGISTERS_reg[45][5]  ( .D(n8511), .CK(CLK), .Q(n15676), .QN(n697)
         );
  DFF_X1 \REGISTERS_reg[45][4]  ( .D(n8510), .CK(CLK), .Q(n15677), .QN(n700)
         );
  DFF_X1 \REGISTERS_reg[45][3]  ( .D(n8509), .CK(CLK), .Q(n15678), .QN(n703)
         );
  DFF_X1 \REGISTERS_reg[45][2]  ( .D(n8508), .CK(CLK), .Q(n15679), .QN(n706)
         );
  DFF_X1 \REGISTERS_reg[45][1]  ( .D(n8507), .CK(CLK), .Q(n15680), .QN(n709)
         );
  DFF_X1 \REGISTERS_reg[45][0]  ( .D(n8506), .CK(CLK), .Q(n15681), .QN(n712)
         );
  DFF_X1 \REGISTERS_reg[40][23]  ( .D(n8689), .CK(CLK), .Q(n15682), .QN(n945)
         );
  DFF_X1 \REGISTERS_reg[40][22]  ( .D(n8688), .CK(CLK), .Q(n15683), .QN(n946)
         );
  DFF_X1 \REGISTERS_reg[40][21]  ( .D(n8687), .CK(CLK), .Q(n15684), .QN(n947)
         );
  DFF_X1 \REGISTERS_reg[40][20]  ( .D(n8686), .CK(CLK), .Q(n15685), .QN(n948)
         );
  DFF_X1 \REGISTERS_reg[40][19]  ( .D(n8685), .CK(CLK), .Q(n15686), .QN(n949)
         );
  DFF_X1 \REGISTERS_reg[40][18]  ( .D(n8684), .CK(CLK), .Q(n15687), .QN(n950)
         );
  DFF_X1 \REGISTERS_reg[40][17]  ( .D(n8683), .CK(CLK), .Q(n15688), .QN(n951)
         );
  DFF_X1 \REGISTERS_reg[40][16]  ( .D(n8682), .CK(CLK), .Q(n15689), .QN(n952)
         );
  DFF_X1 \REGISTERS_reg[40][15]  ( .D(n8681), .CK(CLK), .Q(n15690), .QN(n953)
         );
  DFF_X1 \REGISTERS_reg[40][14]  ( .D(n8680), .CK(CLK), .Q(n15691), .QN(n954)
         );
  DFF_X1 \REGISTERS_reg[40][13]  ( .D(n8679), .CK(CLK), .Q(n15692), .QN(n955)
         );
  DFF_X1 \REGISTERS_reg[40][12]  ( .D(n8678), .CK(CLK), .Q(n15693), .QN(n956)
         );
  DFF_X1 \REGISTERS_reg[40][11]  ( .D(n8677), .CK(CLK), .Q(n15694), .QN(n957)
         );
  DFF_X1 \REGISTERS_reg[40][10]  ( .D(n8676), .CK(CLK), .Q(n15695), .QN(n958)
         );
  DFF_X1 \REGISTERS_reg[40][9]  ( .D(n8675), .CK(CLK), .Q(n15696), .QN(n959)
         );
  DFF_X1 \REGISTERS_reg[40][8]  ( .D(n8674), .CK(CLK), .Q(n15697), .QN(n960)
         );
  DFF_X1 \REGISTERS_reg[40][7]  ( .D(n8673), .CK(CLK), .Q(n15698), .QN(n961)
         );
  DFF_X1 \REGISTERS_reg[40][6]  ( .D(n8672), .CK(CLK), .Q(n15699), .QN(n962)
         );
  DFF_X1 \REGISTERS_reg[40][5]  ( .D(n8671), .CK(CLK), .Q(n15700), .QN(n963)
         );
  DFF_X1 \REGISTERS_reg[40][4]  ( .D(n8670), .CK(CLK), .Q(n15701), .QN(n964)
         );
  DFF_X1 \REGISTERS_reg[40][3]  ( .D(n8669), .CK(CLK), .Q(n15702), .QN(n965)
         );
  DFF_X1 \REGISTERS_reg[40][2]  ( .D(n8668), .CK(CLK), .Q(n15703), .QN(n966)
         );
  DFF_X1 \REGISTERS_reg[40][1]  ( .D(n8667), .CK(CLK), .Q(n15704), .QN(n967)
         );
  DFF_X1 \REGISTERS_reg[40][0]  ( .D(n8666), .CK(CLK), .Q(n15705), .QN(n968)
         );
  DFF_X1 \REGISTERS_reg[39][23]  ( .D(n8721), .CK(CLK), .Q(n15706), .QN(n5791)
         );
  DFF_X1 \REGISTERS_reg[39][22]  ( .D(n8720), .CK(CLK), .Q(n15707), .QN(n5787)
         );
  DFF_X1 \REGISTERS_reg[39][21]  ( .D(n8719), .CK(CLK), .Q(n15708), .QN(n5783)
         );
  DFF_X1 \REGISTERS_reg[39][20]  ( .D(n8718), .CK(CLK), .Q(n15709), .QN(n5779)
         );
  DFF_X1 \REGISTERS_reg[39][19]  ( .D(n8717), .CK(CLK), .Q(n15710), .QN(n5775)
         );
  DFF_X1 \REGISTERS_reg[39][18]  ( .D(n8716), .CK(CLK), .Q(n15711), .QN(n5771)
         );
  DFF_X1 \REGISTERS_reg[39][17]  ( .D(n8715), .CK(CLK), .Q(n15712), .QN(n5767)
         );
  DFF_X1 \REGISTERS_reg[39][16]  ( .D(n8714), .CK(CLK), .Q(n15713), .QN(n5763)
         );
  DFF_X1 \REGISTERS_reg[39][15]  ( .D(n8713), .CK(CLK), .Q(n15714), .QN(n5759)
         );
  DFF_X1 \REGISTERS_reg[39][14]  ( .D(n8712), .CK(CLK), .Q(n15715), .QN(n5755)
         );
  DFF_X1 \REGISTERS_reg[39][13]  ( .D(n8711), .CK(CLK), .Q(n15716), .QN(n5751)
         );
  DFF_X1 \REGISTERS_reg[39][12]  ( .D(n8710), .CK(CLK), .Q(n15717), .QN(n5747)
         );
  DFF_X1 \REGISTERS_reg[39][11]  ( .D(n8709), .CK(CLK), .Q(n15718), .QN(n5743)
         );
  DFF_X1 \REGISTERS_reg[39][10]  ( .D(n8708), .CK(CLK), .Q(n15719), .QN(n5739)
         );
  DFF_X1 \REGISTERS_reg[39][9]  ( .D(n8707), .CK(CLK), .Q(n15720), .QN(n5735)
         );
  DFF_X1 \REGISTERS_reg[39][8]  ( .D(n8706), .CK(CLK), .Q(n15721), .QN(n5731)
         );
  DFF_X1 \REGISTERS_reg[39][7]  ( .D(n8705), .CK(CLK), .Q(n15722), .QN(n5727)
         );
  DFF_X1 \REGISTERS_reg[39][6]  ( .D(n8704), .CK(CLK), .Q(n15723), .QN(n5723)
         );
  DFF_X1 \REGISTERS_reg[39][5]  ( .D(n8703), .CK(CLK), .Q(n15724), .QN(n5719)
         );
  DFF_X1 \REGISTERS_reg[39][4]  ( .D(n8702), .CK(CLK), .Q(n15725), .QN(n5715)
         );
  DFF_X1 \REGISTERS_reg[39][3]  ( .D(n8701), .CK(CLK), .Q(n15726), .QN(n5711)
         );
  DFF_X1 \REGISTERS_reg[39][2]  ( .D(n8700), .CK(CLK), .Q(n15727), .QN(n5707)
         );
  DFF_X1 \REGISTERS_reg[39][1]  ( .D(n8699), .CK(CLK), .Q(n15728), .QN(n5703)
         );
  DFF_X1 \REGISTERS_reg[39][0]  ( .D(n8698), .CK(CLK), .Q(n15729), .QN(n5699)
         );
  DFF_X1 \REGISTERS_reg[38][31]  ( .D(n8761), .CK(CLK), .Q(n15730), .QN(n5822)
         );
  DFF_X1 \REGISTERS_reg[38][30]  ( .D(n8760), .CK(CLK), .Q(n15731), .QN(n5818)
         );
  DFF_X1 \REGISTERS_reg[38][29]  ( .D(n8759), .CK(CLK), .Q(n15732), .QN(n5814)
         );
  DFF_X1 \REGISTERS_reg[38][28]  ( .D(n8758), .CK(CLK), .Q(n15733), .QN(n5810)
         );
  DFF_X1 \REGISTERS_reg[38][27]  ( .D(n8757), .CK(CLK), .Q(n15734), .QN(n5806)
         );
  DFF_X1 \REGISTERS_reg[38][26]  ( .D(n8756), .CK(CLK), .Q(n15735), .QN(n5802)
         );
  DFF_X1 \REGISTERS_reg[38][25]  ( .D(n8755), .CK(CLK), .Q(n15736), .QN(n5798)
         );
  DFF_X1 \REGISTERS_reg[38][24]  ( .D(n8754), .CK(CLK), .Q(n15737), .QN(n5794)
         );
  DFF_X1 \REGISTERS_reg[38][23]  ( .D(n8753), .CK(CLK), .Q(n15738), .QN(n5790)
         );
  DFF_X1 \REGISTERS_reg[38][22]  ( .D(n8752), .CK(CLK), .Q(n15739), .QN(n5786)
         );
  DFF_X1 \REGISTERS_reg[38][21]  ( .D(n8751), .CK(CLK), .Q(n15740), .QN(n5782)
         );
  DFF_X1 \REGISTERS_reg[38][20]  ( .D(n8750), .CK(CLK), .Q(n15741), .QN(n5778)
         );
  DFF_X1 \REGISTERS_reg[32][23]  ( .D(n8945), .CK(CLK), .Q(n14668), .QN(n7069)
         );
  DFF_X1 \REGISTERS_reg[32][22]  ( .D(n8944), .CK(CLK), .Q(n14669), .QN(n7068)
         );
  DFF_X1 \REGISTERS_reg[32][21]  ( .D(n8943), .CK(CLK), .Q(n14670), .QN(n7067)
         );
  DFF_X1 \REGISTERS_reg[32][20]  ( .D(n8942), .CK(CLK), .Q(n14671), .QN(n7066)
         );
  DFF_X1 \REGISTERS_reg[32][19]  ( .D(n8941), .CK(CLK), .Q(n14672), .QN(n7065)
         );
  DFF_X1 \REGISTERS_reg[32][18]  ( .D(n8940), .CK(CLK), .Q(n14673), .QN(n7064)
         );
  DFF_X1 \REGISTERS_reg[32][17]  ( .D(n8939), .CK(CLK), .Q(n14674), .QN(n7063)
         );
  DFF_X1 \REGISTERS_reg[32][16]  ( .D(n8938), .CK(CLK), .Q(n14675), .QN(n7062)
         );
  DFF_X1 \REGISTERS_reg[32][15]  ( .D(n8937), .CK(CLK), .Q(n14676), .QN(n7061)
         );
  DFF_X1 \REGISTERS_reg[32][14]  ( .D(n8936), .CK(CLK), .Q(n14677), .QN(n7060)
         );
  DFF_X1 \REGISTERS_reg[32][13]  ( .D(n8935), .CK(CLK), .Q(n14678), .QN(n7059)
         );
  DFF_X1 \REGISTERS_reg[32][12]  ( .D(n8934), .CK(CLK), .Q(n14679), .QN(n7058)
         );
  DFF_X1 \REGISTERS_reg[32][11]  ( .D(n8933), .CK(CLK), .Q(n14680), .QN(n7057)
         );
  DFF_X1 \REGISTERS_reg[32][10]  ( .D(n8932), .CK(CLK), .Q(n14681), .QN(n7056)
         );
  DFF_X1 \REGISTERS_reg[32][9]  ( .D(n8931), .CK(CLK), .Q(n14682), .QN(n7055)
         );
  DFF_X1 \REGISTERS_reg[32][8]  ( .D(n8930), .CK(CLK), .Q(n14683), .QN(n7054)
         );
  DFF_X1 \REGISTERS_reg[32][7]  ( .D(n8929), .CK(CLK), .Q(n14684), .QN(n7053)
         );
  DFF_X1 \REGISTERS_reg[32][6]  ( .D(n8928), .CK(CLK), .Q(n14685), .QN(n7052)
         );
  DFF_X1 \REGISTERS_reg[32][5]  ( .D(n8927), .CK(CLK), .Q(n14686), .QN(n7051)
         );
  DFF_X1 \REGISTERS_reg[32][4]  ( .D(n8926), .CK(CLK), .Q(n14687), .QN(n7050)
         );
  DFF_X1 \REGISTERS_reg[32][3]  ( .D(n8925), .CK(CLK), .Q(n14688), .QN(n7049)
         );
  DFF_X1 \REGISTERS_reg[32][2]  ( .D(n8924), .CK(CLK), .Q(n14689), .QN(n7048)
         );
  DFF_X1 \REGISTERS_reg[32][1]  ( .D(n8923), .CK(CLK), .Q(n14690), .QN(n7047)
         );
  DFF_X1 \REGISTERS_reg[32][0]  ( .D(n8922), .CK(CLK), .Q(n14691), .QN(n7046)
         );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n8977), .CK(CLK), .Q(n15742), .QN(n913)
         );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n8976), .CK(CLK), .Q(n15743), .QN(n914)
         );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n8975), .CK(CLK), .Q(n15744), .QN(n915)
         );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n8974), .CK(CLK), .Q(n15745), .QN(n916)
         );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n8973), .CK(CLK), .Q(n15746), .QN(n917)
         );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n8972), .CK(CLK), .Q(n15747), .QN(n918)
         );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n8971), .CK(CLK), .Q(n15748), .QN(n919)
         );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n8970), .CK(CLK), .Q(n15749), .QN(n920)
         );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n8969), .CK(CLK), .Q(n15750), .QN(n921)
         );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n8968), .CK(CLK), .Q(n15751), .QN(n922)
         );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n8967), .CK(CLK), .Q(n15752), .QN(n923)
         );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n8966), .CK(CLK), .Q(n15753), .QN(n924)
         );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n8965), .CK(CLK), .Q(n15754), .QN(n925)
         );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n8964), .CK(CLK), .Q(n15755), .QN(n926)
         );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n8963), .CK(CLK), .Q(n15756), .QN(n927)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n8962), .CK(CLK), .Q(n15757), .QN(n928)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n8961), .CK(CLK), .Q(n15758), .QN(n929)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n8960), .CK(CLK), .Q(n15759), .QN(n930)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n8959), .CK(CLK), .Q(n15760), .QN(n931)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n8958), .CK(CLK), .Q(n15761), .QN(n932)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n8957), .CK(CLK), .Q(n15762), .QN(n933)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n8956), .CK(CLK), .Q(n15763), .QN(n934)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n8955), .CK(CLK), .Q(n15764), .QN(n935)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n8954), .CK(CLK), .Q(n15765), .QN(n936)
         );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n9009), .CK(CLK), .Q(n15766), .QN(n5613)
         );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n9008), .CK(CLK), .Q(n15767), .QN(n5603)
         );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n9007), .CK(CLK), .Q(n15768), .QN(n5593)
         );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n9006), .CK(CLK), .Q(n15769), .QN(n5583)
         );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n9005), .CK(CLK), .Q(n15770), .QN(n5573)
         );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n9004), .CK(CLK), .Q(n15771), .QN(n5563)
         );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n9003), .CK(CLK), .Q(n15772), .QN(n5553)
         );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n9002), .CK(CLK), .Q(n15773), .QN(n5543)
         );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n9001), .CK(CLK), .Q(n15774), .QN(n5533)
         );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n9000), .CK(CLK), .Q(n15775), .QN(n5523)
         );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n8999), .CK(CLK), .Q(n15776), .QN(n5513)
         );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n8998), .CK(CLK), .Q(n15777), .QN(n5503)
         );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n8997), .CK(CLK), .Q(n15778), .QN(n5493)
         );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n8996), .CK(CLK), .Q(n15779), .QN(n5483)
         );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n8995), .CK(CLK), .Q(n15780), .QN(n5473)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n8994), .CK(CLK), .Q(n15781), .QN(n5463)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n8993), .CK(CLK), .Q(n15782), .QN(n5453)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n8992), .CK(CLK), .Q(n15783), .QN(n5443)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n8991), .CK(CLK), .Q(n15784), .QN(n5433)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n8990), .CK(CLK), .Q(n15785), .QN(n5423)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n8989), .CK(CLK), .Q(n15786), .QN(n5413)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n8988), .CK(CLK), .Q(n15787), .QN(n5403)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n8987), .CK(CLK), .Q(n15788), .QN(n5393)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n8986), .CK(CLK), .Q(n15789), .QN(n5383)
         );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n9041), .CK(CLK), .Q(n15798), .QN(n5612)
         );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n9040), .CK(CLK), .Q(n15799), .QN(n5602)
         );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n9039), .CK(CLK), .Q(n15800), .QN(n5592)
         );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n9038), .CK(CLK), .Q(n15801), .QN(n5582)
         );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n9037), .CK(CLK), .Q(n15802), .QN(n5572)
         );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n9036), .CK(CLK), .Q(n15803), .QN(n5562)
         );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n9035), .CK(CLK), .Q(n15804), .QN(n5552)
         );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n9034), .CK(CLK), .Q(n15805), .QN(n5542)
         );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n9033), .CK(CLK), .Q(n15806), .QN(n5532)
         );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n9032), .CK(CLK), .Q(n15807), .QN(n5522)
         );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n9031), .CK(CLK), .Q(n15808), .QN(n5512)
         );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n9030), .CK(CLK), .Q(n15809), .QN(n5502)
         );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n9029), .CK(CLK), .Q(n15810), .QN(n5492)
         );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n9028), .CK(CLK), .Q(n15811), .QN(n5482)
         );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n9027), .CK(CLK), .Q(n15812), .QN(n5472)
         );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n9026), .CK(CLK), .Q(n15813), .QN(n5462)
         );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n9025), .CK(CLK), .Q(n15633), .QN(n5452)
         );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n9024), .CK(CLK), .Q(n14653), .QN(n7159)
         );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n9023), .CK(CLK), .Q(n14654), .QN(n7158)
         );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n9022), .CK(CLK), .Q(n14655), .QN(n7157)
         );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n9021), .CK(CLK), .Q(n14656), .QN(n7156)
         );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n9020), .CK(CLK), .Q(n14657), .QN(n7155)
         );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n9019), .CK(CLK), .Q(n14658), .QN(n7154)
         );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n9018), .CK(CLK), .Q(n14659), .QN(n7153)
         );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n9233), .CK(CLK), .Q(n14469), .QN(n7093)
         );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n9232), .CK(CLK), .Q(n14470), .QN(n7092)
         );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n9231), .CK(CLK), .Q(n14471), .QN(n7091)
         );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n9230), .CK(CLK), .Q(n14472), .QN(n7090)
         );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n9229), .CK(CLK), .Q(n14473), .QN(n7089)
         );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n9228), .CK(CLK), .Q(n14474), .QN(n7088)
         );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n9227), .CK(CLK), .Q(n14475), .QN(n7087)
         );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n9226), .CK(CLK), .Q(n14476), .QN(n7086)
         );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n9225), .CK(CLK), .Q(n14477), .QN(n7085)
         );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n9224), .CK(CLK), .Q(n14478), .QN(n7084)
         );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n9223), .CK(CLK), .Q(n14479), .QN(n7083)
         );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n9222), .CK(CLK), .Q(n14480), .QN(n7082)
         );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n9221), .CK(CLK), .Q(n14481), .QN(n7081)
         );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n9220), .CK(CLK), .Q(n14482), .QN(n7080)
         );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n9219), .CK(CLK), .Q(n14483), .QN(n7079)
         );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n9218), .CK(CLK), .Q(n14484), .QN(n7078)
         );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n9217), .CK(CLK), .Q(n14485), .QN(n7077)
         );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n9216), .CK(CLK), .Q(n14486), .QN(n7076)
         );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n9215), .CK(CLK), .Q(n14487), .QN(n7075)
         );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n9214), .CK(CLK), .Q(n14488), .QN(n7074)
         );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n9213), .CK(CLK), .Q(n14489), .QN(n7073)
         );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n9212), .CK(CLK), .Q(n14490), .QN(n7072)
         );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n9211), .CK(CLK), .Q(n14491), .QN(n7071)
         );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n9210), .CK(CLK), .Q(n14492), .QN(n7070)
         );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n9265), .CK(CLK), .Q(n15814), .QN(n881)
         );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n9264), .CK(CLK), .Q(n15815), .QN(n882)
         );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n9263), .CK(CLK), .Q(n15816), .QN(n883)
         );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n9262), .CK(CLK), .Q(n15817), .QN(n884)
         );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n9261), .CK(CLK), .Q(n15818), .QN(n885)
         );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n9260), .CK(CLK), .Q(n15819), .QN(n886)
         );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n9259), .CK(CLK), .Q(n15820), .QN(n887)
         );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n9258), .CK(CLK), .Q(n15821), .QN(n888)
         );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n9257), .CK(CLK), .Q(n15822), .QN(n889)
         );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n9256), .CK(CLK), .Q(n15823), .QN(n890)
         );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n9255), .CK(CLK), .Q(n15824), .QN(n891)
         );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n9254), .CK(CLK), .Q(n15825), .QN(n892)
         );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n9253), .CK(CLK), .Q(n15826), .QN(n893)
         );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n9252), .CK(CLK), .Q(n15827), .QN(n894)
         );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n9251), .CK(CLK), .Q(n15828), .QN(n895)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n9250), .CK(CLK), .Q(n15829), .QN(n896)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n9249), .CK(CLK), .Q(n15830), .QN(n897)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n9248), .CK(CLK), .Q(n15831), .QN(n898)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n9247), .CK(CLK), .Q(n15832), .QN(n899)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n9246), .CK(CLK), .Q(n15833), .QN(n900)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n9245), .CK(CLK), .Q(n15834), .QN(n901)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n9244), .CK(CLK), .Q(n15835), .QN(n902)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n9243), .CK(CLK), .Q(n15836), .QN(n903)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n9242), .CK(CLK), .Q(n15837), .QN(n904)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n9297), .CK(CLK), .Q(n15838), .QN(n5793)
         );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n9296), .CK(CLK), .Q(n15839), .QN(n5789)
         );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n9295), .CK(CLK), .Q(n15840), .QN(n5785)
         );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n9294), .CK(CLK), .Q(n15841), .QN(n5781)
         );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n9293), .CK(CLK), .Q(n15842), .QN(n5777)
         );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n9292), .CK(CLK), .Q(n15843), .QN(n5773)
         );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n9291), .CK(CLK), .Q(n15844), .QN(n5769)
         );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n9290), .CK(CLK), .Q(n15845), .QN(n5765)
         );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n9289), .CK(CLK), .Q(n15846), .QN(n5761)
         );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n9288), .CK(CLK), .Q(n15847), .QN(n5757)
         );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n9287), .CK(CLK), .Q(n15848), .QN(n5753)
         );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n9286), .CK(CLK), .Q(n15849), .QN(n5749)
         );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n9285), .CK(CLK), .Q(n15850), .QN(n5745)
         );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n9284), .CK(CLK), .Q(n15851), .QN(n5741)
         );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n9283), .CK(CLK), .Q(n15852), .QN(n5737)
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n9282), .CK(CLK), .Q(n15853), .QN(n5733)
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n9281), .CK(CLK), .Q(n15854), .QN(n5729)
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n9280), .CK(CLK), .Q(n15855), .QN(n5725)
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n9279), .CK(CLK), .Q(n15856), .QN(n5721)
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n9278), .CK(CLK), .Q(n15857), .QN(n5717)
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n9277), .CK(CLK), .Q(n15858), .QN(n5713)
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n9276), .CK(CLK), .Q(n15859), .QN(n5709)
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n9275), .CK(CLK), .Q(n15860), .QN(n5705)
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n9274), .CK(CLK), .Q(n15861), .QN(n5701)
         );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n9329), .CK(CLK), .Q(n15870), .QN(n5792)
         );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n9328), .CK(CLK), .Q(n15871), .QN(n5788)
         );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n9327), .CK(CLK), .Q(n15872), .QN(n5784)
         );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n9326), .CK(CLK), .Q(n15873), .QN(n5780)
         );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n9325), .CK(CLK), .Q(n15922), .QN(n5776)
         );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n9324), .CK(CLK), .Q(n14440), .QN(n7104)
         );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n9323), .CK(CLK), .Q(n14441), .QN(n7103)
         );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n9322), .CK(CLK), .Q(n14442), .QN(n7102)
         );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n9321), .CK(CLK), .Q(n14443), .QN(n7101)
         );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n9320), .CK(CLK), .Q(n14444), .QN(n7100)
         );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n9319), .CK(CLK), .Q(n14445), .QN(n7099)
         );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n9318), .CK(CLK), .Q(n14446), .QN(n7098)
         );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n9317), .CK(CLK), .Q(n14447), .QN(n7097)
         );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n9316), .CK(CLK), .Q(n14448), .QN(n7096)
         );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n9315), .CK(CLK), .Q(n14449), .QN(n7095)
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n9314), .CK(CLK), .Q(n14450), .QN(n7094)
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n9313), .CK(CLK), .Q(n14451), .QN(n7005)
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n9312), .CK(CLK), .Q(n14452), .QN(n7004)
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n9311), .CK(CLK), .Q(n14453), .QN(n7003)
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n9310), .CK(CLK), .Q(n14454), .QN(n7002)
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n9309), .CK(CLK), .Q(n14455), .QN(n7001)
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n9308), .CK(CLK), .Q(n14456), .QN(n7000)
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n9307), .CK(CLK), .Q(n14457), .QN(n6999)
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n9306), .CK(CLK), .Q(n14458), .QN(n6998)
         );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n9521), .CK(CLK), .Q(n14256), .QN(n7128)
         );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n9520), .CK(CLK), .Q(n14257), .QN(n7127)
         );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n9519), .CK(CLK), .Q(n14258), .QN(n7126)
         );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n9518), .CK(CLK), .Q(n14259), .QN(n7125)
         );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n9517), .CK(CLK), .Q(n14260), .QN(n7124)
         );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n9516), .CK(CLK), .Q(n14261), .QN(n7123)
         );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n9515), .CK(CLK), .Q(n14262), .QN(n7122)
         );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n9514), .CK(CLK), .Q(n14263), .QN(n7121)
         );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n9513), .CK(CLK), .Q(n14264), .QN(n7120)
         );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n9512), .CK(CLK), .Q(n14265), .QN(n7119)
         );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n9511), .CK(CLK), .Q(n14266), .QN(n7118)
         );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n9510), .CK(CLK), .Q(n14267), .QN(n7117)
         );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n9509), .CK(CLK), .Q(n14268), .QN(n7116)
         );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n9508), .CK(CLK), .Q(n14269), .QN(n7115)
         );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n9507), .CK(CLK), .Q(n14270), .QN(n7114)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n9506), .CK(CLK), .Q(n14271), .QN(n7113)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n9505), .CK(CLK), .Q(n14272), .QN(n7112)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n9504), .CK(CLK), .Q(n14273), .QN(n7111)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n9503), .CK(CLK), .Q(n14274), .QN(n7110)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n9502), .CK(CLK), .Q(n14275), .QN(n7109)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n9501), .CK(CLK), .Q(n14276), .QN(n7108)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n9500), .CK(CLK), .Q(n14277), .QN(n7107)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n9499), .CK(CLK), .Q(n14278), .QN(n7106)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n9498), .CK(CLK), .Q(n14279), .QN(n7105)
         );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n9553), .CK(CLK), .Q(n15874), .QN(n849)
         );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n9552), .CK(CLK), .Q(n15875), .QN(n850)
         );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n9551), .CK(CLK), .Q(n15876), .QN(n851)
         );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n9550), .CK(CLK), .Q(n15877), .QN(n852)
         );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n9549), .CK(CLK), .Q(n15878), .QN(n853)
         );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n9548), .CK(CLK), .Q(n15879), .QN(n854)
         );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n9547), .CK(CLK), .Q(n15880), .QN(n855)
         );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n9546), .CK(CLK), .Q(n15881), .QN(n856)
         );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n9545), .CK(CLK), .Q(n15882), .QN(n857)
         );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n9544), .CK(CLK), .Q(n15883), .QN(n858)
         );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n9543), .CK(CLK), .Q(n15884), .QN(n859)
         );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n9542), .CK(CLK), .Q(n15885), .QN(n860)
         );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n9541), .CK(CLK), .Q(n15886), .QN(n861)
         );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n9540), .CK(CLK), .Q(n15887), .QN(n862)
         );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n9539), .CK(CLK), .Q(n15888), .QN(n863)
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n9538), .CK(CLK), .Q(n15889), .QN(n864)
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n9537), .CK(CLK), .Q(n15890), .QN(n865)
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n9536), .CK(CLK), .Q(n15891), .QN(n866)
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n9535), .CK(CLK), .Q(n15892), .QN(n867)
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n9534), .CK(CLK), .Q(n15893), .QN(n868)
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n9533), .CK(CLK), .Q(n15894), .QN(n869)
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n9532), .CK(CLK), .Q(n15895), .QN(n870)
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n9531), .CK(CLK), .Q(n15896), .QN(n871)
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n9530), .CK(CLK), .Q(n15897), .QN(n872)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n9809), .CK(CLK), .Q(n14084), .QN(n7152)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n9808), .CK(CLK), .Q(n14085), .QN(n7151)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n9807), .CK(CLK), .Q(n14086), .QN(n7150)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n9806), .CK(CLK), .Q(n14087), .QN(n7149)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n9805), .CK(CLK), .Q(n14088), .QN(n7148)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n9804), .CK(CLK), .Q(n14089), .QN(n7147)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n9803), .CK(CLK), .Q(n14090), .QN(n7146)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n9802), .CK(CLK), .Q(n14091), .QN(n7145)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n9801), .CK(CLK), .Q(n14092), .QN(n7144)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n9800), .CK(CLK), .Q(n14093), .QN(n7143)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n9799), .CK(CLK), .Q(n14094), .QN(n7142)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n9798), .CK(CLK), .Q(n14095), .QN(n7141)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n9797), .CK(CLK), .Q(n14096), .QN(n7140)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n9796), .CK(CLK), .Q(n14097), .QN(n7139)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n9795), .CK(CLK), .Q(n14098), .QN(n7138)
         );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n9794), .CK(CLK), .Q(n14099), .QN(n7137)
         );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n9793), .CK(CLK), .Q(n14100), .QN(n7136)
         );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n9792), .CK(CLK), .Q(n14101), .QN(n7135)
         );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n9791), .CK(CLK), .Q(n14102), .QN(n7134)
         );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n9790), .CK(CLK), .Q(n14103), .QN(n7133)
         );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n9789), .CK(CLK), .Q(n14104), .QN(n7132)
         );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n9788), .CK(CLK), .Q(n14105), .QN(n7131)
         );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n9787), .CK(CLK), .Q(n14106), .QN(n7130)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n9786), .CK(CLK), .Q(n14107), .QN(n7129)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n9841), .CK(CLK), .Q(n15898), .QN(n817)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n9840), .CK(CLK), .Q(n15899), .QN(n818)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n9839), .CK(CLK), .Q(n15900), .QN(n819)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n9838), .CK(CLK), .Q(n15901), .QN(n820)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n9837), .CK(CLK), .Q(n15902), .QN(n821)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n9836), .CK(CLK), .Q(n15903), .QN(n822)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n9835), .CK(CLK), .Q(n15904), .QN(n823)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n9834), .CK(CLK), .Q(n15905), .QN(n824)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n9833), .CK(CLK), .Q(n15906), .QN(n825)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n9832), .CK(CLK), .Q(n15907), .QN(n826)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n9831), .CK(CLK), .Q(n15908), .QN(n827)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n9830), .CK(CLK), .Q(n15909), .QN(n828)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n9829), .CK(CLK), .Q(n15910), .QN(n829)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n9828), .CK(CLK), .Q(n15911), .QN(n830)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n9827), .CK(CLK), .Q(n15912), .QN(n831) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n9826), .CK(CLK), .Q(n15913), .QN(n832) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n9825), .CK(CLK), .Q(n15914), .QN(n833) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n9824), .CK(CLK), .Q(n15915), .QN(n834) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n9823), .CK(CLK), .Q(n15916), .QN(n835) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n9822), .CK(CLK), .Q(n15917), .QN(n836) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n9821), .CK(CLK), .Q(n15918), .QN(n837) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n9820), .CK(CLK), .Q(n15919), .QN(n838) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n9819), .CK(CLK), .Q(n15920), .QN(n839) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n9818), .CK(CLK), .Q(n15921), .QN(n840) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n9593), .CK(CLK), .Q(n15931), .QN(n5695)
         );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n9592), .CK(CLK), .Q(n15932), .QN(n5685)
         );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n9591), .CK(CLK), .Q(n15933), .QN(n5675)
         );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n9590), .CK(CLK), .Q(n15934), .QN(n5665)
         );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n9589), .CK(CLK), .Q(n15935), .QN(n5655)
         );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n9588), .CK(CLK), .Q(n15936), .QN(n5645)
         );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n9587), .CK(CLK), .Q(n15937), .QN(n5635)
         );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n9586), .CK(CLK), .Q(n15938), .QN(n5625)
         );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n9689), .CK(CLK), .Q(n14204), .QN(n6921)
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n9688), .CK(CLK), .Q(n14205), .QN(n6920)
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n9687), .CK(CLK), .Q(n14206), .QN(n6919)
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n9686), .CK(CLK), .Q(n14207), .QN(n6918)
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n9685), .CK(CLK), .Q(n14208), .QN(n6917)
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n9684), .CK(CLK), .Q(n14209), .QN(n6916)
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n9683), .CK(CLK), .Q(n14210), .QN(n6915)
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n9682), .CK(CLK), .Q(n14211), .QN(n6914)
         );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n9881), .CK(CLK), .Q(n15939), .QN(n5697)
         );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n9880), .CK(CLK), .Q(n15940), .QN(n5687)
         );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n9879), .CK(CLK), .Q(n15941), .QN(n5677)
         );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n9878), .CK(CLK), .Q(n15942), .QN(n5667)
         );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n9877), .CK(CLK), .Q(n15943), .QN(n5657)
         );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n9876), .CK(CLK), .Q(n15944), .QN(n5647)
         );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n9875), .CK(CLK), .Q(n15945), .QN(n5637)
         );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n9874), .CK(CLK), .Q(n15946), .QN(n5627)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n9977), .CK(CLK), .Q(n14028), .QN(n6937)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n9976), .CK(CLK), .Q(n14029), .QN(n6936)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n9975), .CK(CLK), .Q(n14030), .QN(n6935)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n9974), .CK(CLK), .Q(n14031), .QN(n6934)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n9973), .CK(CLK), .Q(n14032), .QN(n6933)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n9972), .CK(CLK), .Q(n14033), .QN(n6932)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n9971), .CK(CLK), .Q(n14034), .QN(n6931)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n9970), .CK(CLK), .Q(n14035), .QN(n6930)
         );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n9657), .CK(CLK), .Q(n14216), .QN(n6793)
         );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n9656), .CK(CLK), .Q(n14217), .QN(n6792)
         );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n9655), .CK(CLK), .Q(n14218), .QN(n6791)
         );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n9654), .CK(CLK), .Q(n14219), .QN(n6790)
         );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n9653), .CK(CLK), .Q(n14220), .QN(n6789)
         );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n9652), .CK(CLK), .Q(n14221), .QN(n6788)
         );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n9651), .CK(CLK), .Q(n14222), .QN(n6787)
         );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n9650), .CK(CLK), .Q(n14223), .QN(n6786)
         );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n9945), .CK(CLK), .Q(n14044), .QN(n6809)
         );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n9944), .CK(CLK), .Q(n14045), .QN(n6808)
         );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n9943), .CK(CLK), .Q(n14046), .QN(n6807)
         );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n9942), .CK(CLK), .Q(n14047), .QN(n6806)
         );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n9941), .CK(CLK), .Q(n14048), .QN(n6805)
         );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n9940), .CK(CLK), .Q(n14049), .QN(n6804)
         );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n9939), .CK(CLK), .Q(n14050), .QN(n6803)
         );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n9938), .CK(CLK), .Q(n14051), .QN(n6802)
         );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n9585), .CK(CLK), .Q(n15971), .QN(n5615)
         );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n9584), .CK(CLK), .Q(n15972), .QN(n5605)
         );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n9583), .CK(CLK), .Q(n15973), .QN(n5595)
         );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n9582), .CK(CLK), .Q(n15974), .QN(n5585)
         );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n9581), .CK(CLK), .Q(n15975), .QN(n5575)
         );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n9580), .CK(CLK), .Q(n15976), .QN(n5565)
         );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n9579), .CK(CLK), .Q(n15977), .QN(n5555)
         );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n9578), .CK(CLK), .Q(n15978), .QN(n5545)
         );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n9577), .CK(CLK), .Q(n15979), .QN(n5535)
         );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n9576), .CK(CLK), .Q(n15980), .QN(n5525)
         );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n9575), .CK(CLK), .Q(n15981), .QN(n5515)
         );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n9574), .CK(CLK), .Q(n15982), .QN(n5505)
         );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n9573), .CK(CLK), .Q(n15983), .QN(n5495)
         );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n9572), .CK(CLK), .Q(n15984), .QN(n5485)
         );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n9571), .CK(CLK), .Q(n15985), .QN(n5475)
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n9570), .CK(CLK), .Q(n15986), .QN(n5465)
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n9569), .CK(CLK), .Q(n15987), .QN(n5455)
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n9568), .CK(CLK), .Q(n15988), .QN(n5445)
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n9567), .CK(CLK), .Q(n15989), .QN(n5435)
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n9566), .CK(CLK), .Q(n15990), .QN(n5425)
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n9565), .CK(CLK), .Q(n15991), .QN(n5415)
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n9564), .CK(CLK), .Q(n15992), .QN(n5405)
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n9563), .CK(CLK), .Q(n15993), .QN(n5395)
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n9562), .CK(CLK), .Q(n15994), .QN(n5385)
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n9681), .CK(CLK), .Q(n14212), .QN(n6941)
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n9680), .CK(CLK), .Q(n14213), .QN(n6940)
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n9679), .CK(CLK), .Q(n14214), .QN(n6939)
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n9678), .CK(CLK), .Q(n14215), .QN(n6938)
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n9677), .CK(CLK), .Q(n16043), .QN(n653)
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n9676), .CK(CLK), .Q(n16044), .QN(n656)
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n9675), .CK(CLK), .Q(n16045), .QN(n659)
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n9674), .CK(CLK), .Q(n16046), .QN(n662)
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n9673), .CK(CLK), .Q(n16047), .QN(n665)
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n9672), .CK(CLK), .Q(n16048), .QN(n668)
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n9671), .CK(CLK), .Q(n16049), .QN(n671)
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n9670), .CK(CLK), .Q(n16050), .QN(n674)
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n9669), .CK(CLK), .Q(n15995), .QN(n677)
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n9668), .CK(CLK), .Q(n15996), .QN(n680)
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n9667), .CK(CLK), .Q(n15997), .QN(n683) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n9666), .CK(CLK), .Q(n15998), .QN(n686) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n9665), .CK(CLK), .Q(n15999), .QN(n689) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n9664), .CK(CLK), .Q(n16000), .QN(n692) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n9663), .CK(CLK), .Q(n16001), .QN(n695) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n9662), .CK(CLK), .Q(n16002), .QN(n698) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n9661), .CK(CLK), .Q(n16003), .QN(n701) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n9660), .CK(CLK), .Q(n16004), .QN(n704) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n9659), .CK(CLK), .Q(n16005), .QN(n707) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n9658), .CK(CLK), .Q(n16006), .QN(n710) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n9873), .CK(CLK), .Q(n16007), .QN(n5617)
         );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n9872), .CK(CLK), .Q(n16008), .QN(n5607)
         );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n9871), .CK(CLK), .Q(n16009), .QN(n5597)
         );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n9870), .CK(CLK), .Q(n16010), .QN(n5587)
         );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n9869), .CK(CLK), .Q(n16011), .QN(n5577)
         );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n9868), .CK(CLK), .Q(n16012), .QN(n5567)
         );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n9867), .CK(CLK), .Q(n16013), .QN(n5557)
         );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n9866), .CK(CLK), .Q(n16014), .QN(n5547)
         );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n9865), .CK(CLK), .Q(n16015), .QN(n5537)
         );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n9864), .CK(CLK), .Q(n16016), .QN(n5527)
         );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n9863), .CK(CLK), .Q(n16017), .QN(n5517)
         );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n9862), .CK(CLK), .Q(n16018), .QN(n5507)
         );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n9861), .CK(CLK), .Q(n16019), .QN(n5497)
         );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n9860), .CK(CLK), .Q(n16020), .QN(n5487)
         );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n9859), .CK(CLK), .Q(n16021), .QN(n5477)
         );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n9858), .CK(CLK), .Q(n16022), .QN(n5467)
         );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n9857), .CK(CLK), .Q(n16023), .QN(n5457)
         );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n9856), .CK(CLK), .Q(n16024), .QN(n5447)
         );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n9855), .CK(CLK), .Q(n16025), .QN(n5437)
         );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n9854), .CK(CLK), .Q(n16026), .QN(n5427)
         );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n9853), .CK(CLK), .Q(n16027), .QN(n5417)
         );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n9852), .CK(CLK), .Q(n16028), .QN(n5407)
         );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n9851), .CK(CLK), .Q(n16029), .QN(n5397)
         );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n9850), .CK(CLK), .Q(n16030), .QN(n5387)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n9969), .CK(CLK), .Q(n14036), .QN(n6929)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n9968), .CK(CLK), .Q(n14037), .QN(n6928)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n9967), .CK(CLK), .Q(n14038), .QN(n6927)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n9966), .CK(CLK), .Q(n14039), .QN(n6926)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n9965), .CK(CLK), .Q(n14040), .QN(n6925)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n9964), .CK(CLK), .Q(n14041), .QN(n6924)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n9963), .CK(CLK), .Q(n14042), .QN(n6923)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n9962), .CK(CLK), .Q(n14043), .QN(n6922)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n9961), .CK(CLK), .Q(n16051), .QN(n666)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n9960), .CK(CLK), .Q(n16052), .QN(n669)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n9959), .CK(CLK), .Q(n16053), .QN(n672)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n9958), .CK(CLK), .Q(n16054), .QN(n675)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n9957), .CK(CLK), .Q(n16031), .QN(n678)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n9956), .CK(CLK), .Q(n16032), .QN(n681)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n9955), .CK(CLK), .Q(n16033), .QN(n684) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n9954), .CK(CLK), .Q(n16034), .QN(n687) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n9953), .CK(CLK), .Q(n16035), .QN(n690) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n9952), .CK(CLK), .Q(n16036), .QN(n693) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n9951), .CK(CLK), .Q(n16037), .QN(n696) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n9950), .CK(CLK), .Q(n16038), .QN(n699) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n9949), .CK(CLK), .Q(n16039), .QN(n702) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n9948), .CK(CLK), .Q(n16040), .QN(n705) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n9947), .CK(CLK), .Q(n16041), .QN(n708) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n9946), .CK(CLK), .Q(n16042), .QN(n711) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n9649), .CK(CLK), .Q(n14224), .QN(n6813)
         );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n9648), .CK(CLK), .Q(n14225), .QN(n6812)
         );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n9647), .CK(CLK), .Q(n14226), .QN(n6811)
         );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n9646), .CK(CLK), .Q(n14227), .QN(n6810)
         );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n9645), .CK(CLK), .Q(n14228), .QN(n6893)
         );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n9644), .CK(CLK), .Q(n14229), .QN(n6892)
         );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n9643), .CK(CLK), .Q(n14230), .QN(n6891)
         );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n9642), .CK(CLK), .Q(n14231), .QN(n6890)
         );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n9641), .CK(CLK), .Q(n14232), .QN(n6888)
         );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n9640), .CK(CLK), .Q(n14233), .QN(n6886)
         );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n9639), .CK(CLK), .Q(n14234), .QN(n6884)
         );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n9638), .CK(CLK), .Q(n14235), .QN(n6882)
         );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n9637), .CK(CLK), .Q(n14236), .QN(n6881)
         );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n9636), .CK(CLK), .Q(n14237), .QN(n6880)
         );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n9635), .CK(CLK), .Q(n14238), .QN(n6879)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n9634), .CK(CLK), .Q(n14239), .QN(n6878)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n9633), .CK(CLK), .Q(n14240), .QN(n6877)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n9632), .CK(CLK), .Q(n14241), .QN(n6876)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n9631), .CK(CLK), .Q(n14242), .QN(n6875)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n9630), .CK(CLK), .Q(n14243), .QN(n6874)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n9629), .CK(CLK), .Q(n14244), .QN(n6873)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n9628), .CK(CLK), .Q(n14245), .QN(n6872)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n9627), .CK(CLK), .Q(n14246), .QN(n6871)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n9626), .CK(CLK), .Q(n14247), .QN(n6870)
         );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n9937), .CK(CLK), .Q(n14052), .QN(n6801)
         );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n9936), .CK(CLK), .Q(n14053), .QN(n6800)
         );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n9935), .CK(CLK), .Q(n14054), .QN(n6799)
         );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n9934), .CK(CLK), .Q(n14055), .QN(n6798)
         );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n9933), .CK(CLK), .Q(n14056), .QN(n6797)
         );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n9932), .CK(CLK), .Q(n14057), .QN(n6796)
         );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n9931), .CK(CLK), .Q(n14058), .QN(n6795)
         );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n9930), .CK(CLK), .Q(n14059), .QN(n6794)
         );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n9929), .CK(CLK), .Q(n14060), .QN(n6889)
         );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n9928), .CK(CLK), .Q(n14061), .QN(n6887)
         );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n9927), .CK(CLK), .Q(n14062), .QN(n6885)
         );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n9926), .CK(CLK), .Q(n14063), .QN(n6883)
         );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n9925), .CK(CLK), .Q(n14064), .QN(n6841)
         );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n9924), .CK(CLK), .Q(n14065), .QN(n6840)
         );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n9923), .CK(CLK), .Q(n14066), .QN(n6839)
         );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n9922), .CK(CLK), .Q(n14067), .QN(n6838)
         );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n9921), .CK(CLK), .Q(n14068), .QN(n6837)
         );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n9920), .CK(CLK), .Q(n14069), .QN(n6836)
         );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n9919), .CK(CLK), .Q(n14070), .QN(n6835)
         );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n9918), .CK(CLK), .Q(n14071), .QN(n6834)
         );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n9917), .CK(CLK), .Q(n14072), .QN(n6833)
         );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n9916), .CK(CLK), .Q(n14073), .QN(n6832)
         );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n9915), .CK(CLK), .Q(n14074), .QN(n6831)
         );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n9914), .CK(CLK), .Q(n14075), .QN(n6830)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n7609), .CK(CLK), .QN(n1481) );
  DFF_X1 \OUT2_reg[30]  ( .D(n7607), .CK(CLK), .QN(n1482) );
  DFF_X1 \OUT2_reg[29]  ( .D(n7605), .CK(CLK), .QN(n1483) );
  DFF_X1 \OUT2_reg[28]  ( .D(n7603), .CK(CLK), .QN(n1484) );
  DFF_X1 \OUT2_reg[27]  ( .D(n7601), .CK(CLK), .QN(n1485) );
  DFF_X1 \OUT2_reg[26]  ( .D(n7599), .CK(CLK), .QN(n1486) );
  DFF_X1 \OUT2_reg[25]  ( .D(n7597), .CK(CLK), .QN(n1487) );
  DFF_X1 \OUT1_reg[31]  ( .D(n7673), .CK(CLK), .QN(n1449) );
  DFF_X1 \OUT1_reg[30]  ( .D(n7671), .CK(CLK), .QN(n1450) );
  DFF_X1 \OUT1_reg[29]  ( .D(n7669), .CK(CLK), .QN(n1451) );
  DFF_X1 \OUT1_reg[28]  ( .D(n7667), .CK(CLK), .QN(n1452) );
  DFF_X1 \OUT1_reg[27]  ( .D(n7665), .CK(CLK), .QN(n1453) );
  DFF_X1 \OUT1_reg[26]  ( .D(n7663), .CK(CLK), .QN(n1454) );
  DFF_X1 \OUT1_reg[25]  ( .D(n7661), .CK(CLK), .QN(n1455) );
  DFF_X1 \OUT2_reg[24]  ( .D(n7595), .CK(CLK), .QN(n1488) );
  DFF_X1 \OUT1_reg[24]  ( .D(n7659), .CK(CLK), .QN(n1456) );
  NOR3_X1 U3 ( .A1(n16058), .A2(ADD_RD2[3]), .A3(n16057), .ZN(n5710) );
  NOR3_X1 U4 ( .A1(n16068), .A2(ADD_RD2[0]), .A3(n16069), .ZN(n5669) );
  NOR3_X2 U69 ( .A1(n16064), .A2(ADD_RD1[2]), .A3(n16065), .ZN(n4279) );
  NOR3_X1 U70 ( .A1(n16056), .A2(ADD_RD1[3]), .A3(n16055), .ZN(n4299) );
  NOR3_X1 U71 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n16064), .ZN(n4274) );
  NOR3_X1 U72 ( .A1(n16065), .A2(ADD_RD1[0]), .A3(n16066), .ZN(n4276) );
  NOR3_X1 U73 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(ADD_RD1[0]), .ZN(n4271)
         );
  NOR3_X1 U74 ( .A1(n16067), .A2(ADD_RD2[1]), .A3(n16069), .ZN(n5668) );
  NOR3_X1 U75 ( .A1(n16064), .A2(ADD_RD1[1]), .A3(n16066), .ZN(n4275) );
  BUF_X1 U76 ( .A(n2875), .Z(n13797) );
  BUF_X1 U77 ( .A(n2902), .Z(n13743) );
  BUF_X1 U78 ( .A(n2878), .Z(n13791) );
  BUF_X1 U79 ( .A(n2905), .Z(n13737) );
  BUF_X1 U80 ( .A(n2911), .Z(n13725) );
  BUF_X1 U81 ( .A(n2908), .Z(n13731) );
  BUF_X1 U82 ( .A(n2899), .Z(n13749) );
  BUF_X1 U83 ( .A(n2896), .Z(n13755) );
  BUF_X1 U84 ( .A(n2893), .Z(n13761) );
  BUF_X1 U85 ( .A(n2890), .Z(n13767) );
  BUF_X1 U86 ( .A(n2887), .Z(n13773) );
  BUF_X1 U87 ( .A(n2884), .Z(n13779) );
  BUF_X1 U88 ( .A(n2881), .Z(n13785) );
  BUF_X1 U89 ( .A(n2872), .Z(n13803) );
  BUF_X1 U90 ( .A(n2869), .Z(n13809) );
  BUF_X1 U91 ( .A(n2980), .Z(n13527) );
  BUF_X1 U92 ( .A(n2927), .Z(n13683) );
  BUF_X1 U93 ( .A(n2943), .Z(n13635) );
  BUF_X1 U94 ( .A(n2945), .Z(n13629) );
  BUF_X1 U95 ( .A(n2964), .Z(n13575) );
  BUF_X1 U96 ( .A(n3017), .Z(n13437) );
  BUF_X1 U97 ( .A(n3015), .Z(n13443) );
  BUF_X1 U98 ( .A(n3013), .Z(n13449) );
  BUF_X1 U99 ( .A(n3010), .Z(n13455) );
  BUF_X1 U100 ( .A(n3007), .Z(n13461) );
  BUF_X1 U101 ( .A(n3004), .Z(n13467) );
  BUF_X1 U102 ( .A(n3001), .Z(n13473) );
  BUF_X1 U103 ( .A(n2997), .Z(n13479) );
  BUF_X1 U104 ( .A(n2995), .Z(n13485) );
  BUF_X1 U105 ( .A(n2993), .Z(n13491) );
  BUF_X1 U106 ( .A(n2991), .Z(n13497) );
  BUF_X1 U107 ( .A(n2989), .Z(n13503) );
  BUF_X1 U108 ( .A(n2987), .Z(n13509) );
  BUF_X1 U109 ( .A(n2985), .Z(n13515) );
  BUF_X1 U110 ( .A(n2983), .Z(n13521) );
  BUF_X1 U111 ( .A(n2978), .Z(n13533) );
  BUF_X1 U112 ( .A(n2976), .Z(n13539) );
  BUF_X1 U113 ( .A(n2974), .Z(n13545) );
  BUF_X1 U114 ( .A(n2972), .Z(n13551) );
  BUF_X1 U115 ( .A(n2970), .Z(n13557) );
  BUF_X1 U116 ( .A(n2968), .Z(n13563) );
  BUF_X1 U117 ( .A(n2966), .Z(n13569) );
  BUF_X1 U118 ( .A(n2962), .Z(n13581) );
  BUF_X1 U119 ( .A(n2960), .Z(n13587) );
  BUF_X1 U120 ( .A(n2958), .Z(n13593) );
  BUF_X1 U121 ( .A(n2956), .Z(n13599) );
  BUF_X1 U122 ( .A(n2954), .Z(n13605) );
  BUF_X1 U123 ( .A(n2952), .Z(n13611) );
  BUF_X1 U124 ( .A(n2950), .Z(n13617) );
  BUF_X1 U125 ( .A(n2947), .Z(n13623) );
  BUF_X1 U126 ( .A(n2941), .Z(n13641) );
  BUF_X1 U127 ( .A(n2939), .Z(n13647) );
  BUF_X1 U128 ( .A(n2937), .Z(n13653) );
  BUF_X1 U129 ( .A(n2935), .Z(n13659) );
  BUF_X1 U130 ( .A(n2933), .Z(n13665) );
  BUF_X1 U131 ( .A(n2931), .Z(n13671) );
  BUF_X1 U132 ( .A(n2929), .Z(n13677) );
  BUF_X1 U133 ( .A(n2925), .Z(n13689) );
  BUF_X1 U134 ( .A(n2923), .Z(n13695) );
  BUF_X1 U135 ( .A(n2921), .Z(n13701) );
  BUF_X1 U136 ( .A(n2919), .Z(n13707) );
  BUF_X1 U137 ( .A(n2917), .Z(n13713) );
  BUF_X1 U138 ( .A(n2914), .Z(n13719) );
  BUF_X1 U139 ( .A(n3034), .Z(n13395) );
  BUF_X1 U140 ( .A(n3032), .Z(n13401) );
  BUF_X1 U141 ( .A(n3029), .Z(n13407) );
  BUF_X1 U142 ( .A(n3027), .Z(n13413) );
  BUF_X1 U143 ( .A(n3025), .Z(n13419) );
  BUF_X1 U144 ( .A(n3023), .Z(n13425) );
  BUF_X1 U145 ( .A(n3019), .Z(n13431) );
  BUF_X1 U146 ( .A(n3037), .Z(n13386) );
  BUF_X1 U147 ( .A(n2875), .Z(n13796) );
  BUF_X1 U148 ( .A(n2893), .Z(n13760) );
  BUF_X1 U149 ( .A(n2902), .Z(n13742) );
  BUF_X1 U150 ( .A(n2875), .Z(n13795) );
  BUF_X1 U151 ( .A(n2902), .Z(n13741) );
  BUF_X1 U152 ( .A(n2878), .Z(n13790) );
  BUF_X1 U153 ( .A(n2905), .Z(n13736) );
  BUF_X1 U154 ( .A(n2878), .Z(n13789) );
  BUF_X1 U155 ( .A(n2905), .Z(n13735) );
  BUF_X1 U156 ( .A(n2911), .Z(n13724) );
  BUF_X1 U157 ( .A(n2911), .Z(n13723) );
  BUF_X1 U158 ( .A(n2908), .Z(n13730) );
  BUF_X1 U159 ( .A(n2908), .Z(n13729) );
  BUF_X1 U160 ( .A(n2899), .Z(n13748) );
  BUF_X1 U161 ( .A(n2899), .Z(n13747) );
  BUF_X1 U162 ( .A(n2896), .Z(n13754) );
  BUF_X1 U163 ( .A(n2896), .Z(n13753) );
  BUF_X1 U164 ( .A(n2893), .Z(n13759) );
  BUF_X1 U165 ( .A(n2890), .Z(n13766) );
  BUF_X1 U166 ( .A(n2890), .Z(n13765) );
  BUF_X1 U167 ( .A(n2887), .Z(n13772) );
  BUF_X1 U168 ( .A(n2887), .Z(n13771) );
  BUF_X1 U169 ( .A(n2884), .Z(n13778) );
  BUF_X1 U170 ( .A(n2884), .Z(n13777) );
  BUF_X1 U171 ( .A(n2881), .Z(n13784) );
  BUF_X1 U172 ( .A(n2881), .Z(n13783) );
  BUF_X1 U173 ( .A(n2872), .Z(n13802) );
  BUF_X1 U174 ( .A(n2872), .Z(n13801) );
  BUF_X1 U175 ( .A(n2869), .Z(n13808) );
  BUF_X1 U176 ( .A(n2869), .Z(n13807) );
  BUF_X1 U177 ( .A(n2980), .Z(n13526) );
  BUF_X1 U178 ( .A(n2980), .Z(n13525) );
  BUF_X1 U179 ( .A(n2923), .Z(n13693) );
  BUF_X1 U180 ( .A(n2925), .Z(n13688) );
  BUF_X1 U181 ( .A(n2927), .Z(n13682) );
  BUF_X1 U182 ( .A(n2941), .Z(n13640) );
  BUF_X1 U183 ( .A(n2941), .Z(n13639) );
  BUF_X1 U184 ( .A(n2943), .Z(n13634) );
  BUF_X1 U185 ( .A(n2945), .Z(n13628) );
  BUF_X1 U186 ( .A(n2960), .Z(n13585) );
  BUF_X1 U187 ( .A(n2962), .Z(n13580) );
  BUF_X1 U188 ( .A(n2964), .Z(n13574) );
  BUF_X1 U189 ( .A(n2974), .Z(n13544) );
  BUF_X1 U190 ( .A(n2983), .Z(n13520) );
  BUF_X1 U191 ( .A(n2983), .Z(n13519) );
  BUF_X1 U192 ( .A(n2927), .Z(n13681) );
  BUF_X1 U193 ( .A(n2943), .Z(n13633) );
  BUF_X1 U194 ( .A(n2945), .Z(n13627) );
  BUF_X1 U195 ( .A(n2964), .Z(n13573) );
  BUF_X1 U196 ( .A(n3017), .Z(n13436) );
  BUF_X1 U197 ( .A(n3017), .Z(n13435) );
  BUF_X1 U198 ( .A(n3015), .Z(n13442) );
  BUF_X1 U199 ( .A(n3015), .Z(n13441) );
  BUF_X1 U200 ( .A(n3013), .Z(n13448) );
  BUF_X1 U201 ( .A(n3013), .Z(n13447) );
  BUF_X1 U202 ( .A(n3010), .Z(n13454) );
  BUF_X1 U203 ( .A(n3010), .Z(n13453) );
  BUF_X1 U204 ( .A(n3007), .Z(n13460) );
  BUF_X1 U205 ( .A(n3007), .Z(n13459) );
  BUF_X1 U206 ( .A(n3004), .Z(n13466) );
  BUF_X1 U207 ( .A(n3004), .Z(n13465) );
  BUF_X1 U208 ( .A(n3001), .Z(n13472) );
  BUF_X1 U209 ( .A(n3001), .Z(n13471) );
  BUF_X1 U210 ( .A(n2997), .Z(n13478) );
  BUF_X1 U211 ( .A(n2997), .Z(n13477) );
  BUF_X1 U212 ( .A(n2995), .Z(n13484) );
  BUF_X1 U213 ( .A(n2995), .Z(n13483) );
  BUF_X1 U214 ( .A(n2993), .Z(n13490) );
  BUF_X1 U215 ( .A(n2993), .Z(n13489) );
  BUF_X1 U216 ( .A(n2991), .Z(n13496) );
  BUF_X1 U217 ( .A(n2991), .Z(n13495) );
  BUF_X1 U218 ( .A(n2989), .Z(n13502) );
  BUF_X1 U219 ( .A(n2989), .Z(n13501) );
  BUF_X1 U220 ( .A(n2987), .Z(n13508) );
  BUF_X1 U221 ( .A(n2987), .Z(n13507) );
  BUF_X1 U222 ( .A(n2985), .Z(n13514) );
  BUF_X1 U223 ( .A(n2985), .Z(n13513) );
  BUF_X1 U224 ( .A(n2978), .Z(n13532) );
  BUF_X1 U225 ( .A(n2978), .Z(n13531) );
  BUF_X1 U226 ( .A(n2976), .Z(n13538) );
  BUF_X1 U227 ( .A(n2976), .Z(n13537) );
  BUF_X1 U228 ( .A(n2974), .Z(n13543) );
  BUF_X1 U229 ( .A(n2972), .Z(n13550) );
  BUF_X1 U230 ( .A(n2972), .Z(n13549) );
  BUF_X1 U231 ( .A(n2970), .Z(n13556) );
  BUF_X1 U232 ( .A(n2970), .Z(n13555) );
  BUF_X1 U233 ( .A(n2968), .Z(n13562) );
  BUF_X1 U234 ( .A(n2968), .Z(n13561) );
  BUF_X1 U235 ( .A(n2966), .Z(n13568) );
  BUF_X1 U236 ( .A(n2966), .Z(n13567) );
  BUF_X1 U237 ( .A(n2962), .Z(n13579) );
  BUF_X1 U238 ( .A(n2960), .Z(n13586) );
  BUF_X1 U239 ( .A(n2958), .Z(n13592) );
  BUF_X1 U240 ( .A(n2958), .Z(n13591) );
  BUF_X1 U241 ( .A(n2956), .Z(n13598) );
  BUF_X1 U242 ( .A(n2956), .Z(n13597) );
  BUF_X1 U243 ( .A(n2954), .Z(n13604) );
  BUF_X1 U244 ( .A(n2954), .Z(n13603) );
  BUF_X1 U245 ( .A(n2952), .Z(n13610) );
  BUF_X1 U246 ( .A(n2952), .Z(n13609) );
  BUF_X1 U247 ( .A(n2950), .Z(n13616) );
  BUF_X1 U248 ( .A(n2950), .Z(n13615) );
  BUF_X1 U249 ( .A(n2947), .Z(n13622) );
  BUF_X1 U250 ( .A(n2947), .Z(n13621) );
  BUF_X1 U251 ( .A(n2939), .Z(n13646) );
  BUF_X1 U252 ( .A(n2939), .Z(n13645) );
  BUF_X1 U253 ( .A(n2937), .Z(n13652) );
  BUF_X1 U254 ( .A(n2937), .Z(n13651) );
  BUF_X1 U255 ( .A(n2935), .Z(n13658) );
  BUF_X1 U256 ( .A(n2935), .Z(n13657) );
  BUF_X1 U257 ( .A(n2933), .Z(n13664) );
  BUF_X1 U258 ( .A(n2933), .Z(n13663) );
  BUF_X1 U259 ( .A(n2931), .Z(n13670) );
  BUF_X1 U260 ( .A(n2931), .Z(n13669) );
  BUF_X1 U261 ( .A(n2929), .Z(n13676) );
  BUF_X1 U262 ( .A(n2929), .Z(n13675) );
  BUF_X1 U263 ( .A(n2925), .Z(n13687) );
  BUF_X1 U264 ( .A(n2923), .Z(n13694) );
  BUF_X1 U265 ( .A(n2921), .Z(n13700) );
  BUF_X1 U266 ( .A(n2921), .Z(n13699) );
  BUF_X1 U267 ( .A(n2919), .Z(n13706) );
  BUF_X1 U268 ( .A(n2919), .Z(n13705) );
  BUF_X1 U269 ( .A(n2917), .Z(n13712) );
  BUF_X1 U270 ( .A(n2917), .Z(n13711) );
  BUF_X1 U271 ( .A(n2914), .Z(n13718) );
  BUF_X1 U272 ( .A(n2914), .Z(n13717) );
  BUF_X1 U273 ( .A(n4395), .Z(n13012) );
  BUF_X1 U274 ( .A(n4432), .Z(n12931) );
  BUF_X1 U275 ( .A(n4395), .Z(n13013) );
  BUF_X1 U276 ( .A(n4432), .Z(n12932) );
  BUF_X1 U277 ( .A(n3111), .Z(n13240) );
  BUF_X1 U278 ( .A(n3111), .Z(n13241) );
  BUF_X1 U279 ( .A(n3034), .Z(n13394) );
  BUF_X1 U280 ( .A(n3034), .Z(n13393) );
  BUF_X1 U281 ( .A(n3032), .Z(n13400) );
  BUF_X1 U282 ( .A(n3032), .Z(n13399) );
  BUF_X1 U283 ( .A(n3029), .Z(n13406) );
  BUF_X1 U284 ( .A(n3029), .Z(n13405) );
  BUF_X1 U285 ( .A(n3027), .Z(n13412) );
  BUF_X1 U286 ( .A(n3027), .Z(n13411) );
  BUF_X1 U287 ( .A(n3025), .Z(n13418) );
  BUF_X1 U288 ( .A(n3025), .Z(n13417) );
  BUF_X1 U289 ( .A(n3023), .Z(n13424) );
  BUF_X1 U290 ( .A(n3023), .Z(n13423) );
  BUF_X1 U291 ( .A(n3019), .Z(n13430) );
  BUF_X1 U292 ( .A(n3019), .Z(n13429) );
  BUF_X1 U293 ( .A(n3037), .Z(n13384) );
  BUF_X1 U294 ( .A(n3149), .Z(n13156) );
  BUF_X1 U295 ( .A(n3149), .Z(n13157) );
  BUF_X1 U296 ( .A(n3037), .Z(n13385) );
  BUF_X1 U297 ( .A(n4371), .Z(n13060) );
  BUF_X1 U298 ( .A(n4371), .Z(n13061) );
  BUF_X1 U299 ( .A(n3087), .Z(n13288) );
  BUF_X1 U300 ( .A(n3087), .Z(n13289) );
  BUF_X1 U301 ( .A(n2832), .Z(n14021) );
  BUF_X1 U302 ( .A(n4361), .Z(n13084) );
  BUF_X1 U303 ( .A(n4404), .Z(n12988) );
  BUF_X1 U304 ( .A(n4419), .Z(n12961) );
  BUF_X1 U305 ( .A(n4361), .Z(n13085) );
  BUF_X1 U306 ( .A(n4404), .Z(n12989) );
  BUF_X1 U307 ( .A(n4419), .Z(n12962) );
  BUF_X1 U308 ( .A(n3077), .Z(n13312) );
  BUF_X1 U309 ( .A(n3120), .Z(n13216) );
  BUF_X1 U310 ( .A(n3135), .Z(n13189) );
  BUF_X1 U311 ( .A(n3077), .Z(n13313) );
  BUF_X1 U312 ( .A(n3120), .Z(n13217) );
  BUF_X1 U313 ( .A(n3135), .Z(n13190) );
  BUF_X1 U314 ( .A(n2832), .Z(n14020) );
  BUF_X1 U315 ( .A(n2832), .Z(n14019) );
  BUF_X1 U316 ( .A(n4350), .Z(n13102) );
  BUF_X1 U317 ( .A(n4350), .Z(n13103) );
  BUF_X1 U318 ( .A(n3066), .Z(n13330) );
  BUF_X1 U319 ( .A(n3066), .Z(n13331) );
  BUF_X1 U320 ( .A(n4395), .Z(n13014) );
  BUF_X1 U321 ( .A(n4432), .Z(n12933) );
  BUF_X1 U322 ( .A(n3111), .Z(n13242) );
  BUF_X1 U323 ( .A(n4324), .Z(n13150) );
  BUF_X1 U324 ( .A(n4324), .Z(n13151) );
  BUF_X1 U325 ( .A(n3040), .Z(n13378) );
  BUF_X1 U326 ( .A(n3040), .Z(n13379) );
  BUF_X1 U327 ( .A(n4338), .Z(n13132) );
  BUF_X1 U328 ( .A(n4338), .Z(n13133) );
  BUF_X1 U329 ( .A(n3054), .Z(n13360) );
  BUF_X1 U330 ( .A(n3054), .Z(n13361) );
  BUF_X1 U331 ( .A(n3149), .Z(n13158) );
  BUF_X1 U332 ( .A(n4371), .Z(n13062) );
  BUF_X1 U333 ( .A(n3087), .Z(n13290) );
  BUF_X1 U334 ( .A(n4361), .Z(n13086) );
  BUF_X1 U335 ( .A(n4404), .Z(n12990) );
  BUF_X1 U336 ( .A(n4419), .Z(n12963) );
  BUF_X1 U337 ( .A(n3077), .Z(n13314) );
  BUF_X1 U338 ( .A(n3120), .Z(n13218) );
  BUF_X1 U339 ( .A(n3135), .Z(n13191) );
  BUF_X1 U340 ( .A(n4350), .Z(n13104) );
  BUF_X1 U341 ( .A(n3066), .Z(n13332) );
  BUF_X1 U342 ( .A(n4324), .Z(n13152) );
  BUF_X1 U343 ( .A(n3040), .Z(n13380) );
  BUF_X1 U344 ( .A(n4338), .Z(n13134) );
  BUF_X1 U345 ( .A(n3054), .Z(n13362) );
  NOR3_X1 U346 ( .A1(n16058), .A2(n16062), .A3(n16057), .ZN(n5732) );
  NOR3_X1 U347 ( .A1(n16056), .A2(n16061), .A3(n16055), .ZN(n4310) );
  INV_X1 U348 ( .A(n13822), .ZN(n13813) );
  INV_X1 U349 ( .A(n13822), .ZN(n13812) );
  INV_X1 U350 ( .A(n13822), .ZN(n13811) );
  NAND2_X1 U351 ( .A1(n5679), .A2(n5664), .ZN(n4350) );
  NAND2_X1 U352 ( .A1(n4282), .A2(n4273), .ZN(n3066) );
  NAND2_X1 U353 ( .A1(n2982), .A2(n2867), .ZN(n2980) );
  NAND2_X1 U354 ( .A1(n2916), .A2(n2907), .ZN(n2941) );
  NAND2_X1 U355 ( .A1(n2982), .A2(n2871), .ZN(n2983) );
  NAND2_X1 U356 ( .A1(n2916), .A2(n2886), .ZN(n2927) );
  NAND2_X1 U357 ( .A1(n2916), .A2(n2910), .ZN(n2943) );
  NAND2_X1 U358 ( .A1(n2916), .A2(n2913), .ZN(n2945) );
  NAND2_X1 U359 ( .A1(n2949), .A2(n2892), .ZN(n2964) );
  NAND2_X1 U360 ( .A1(n2982), .A2(n2913), .ZN(n3017) );
  NAND2_X1 U361 ( .A1(n2982), .A2(n2910), .ZN(n3015) );
  NAND2_X1 U362 ( .A1(n2982), .A2(n2907), .ZN(n3013) );
  NAND2_X1 U363 ( .A1(n2982), .A2(n2904), .ZN(n3010) );
  NAND2_X1 U364 ( .A1(n2982), .A2(n2901), .ZN(n3007) );
  NAND2_X1 U365 ( .A1(n2982), .A2(n2898), .ZN(n3004) );
  NAND2_X1 U366 ( .A1(n2982), .A2(n2895), .ZN(n3001) );
  NAND2_X1 U367 ( .A1(n2982), .A2(n2892), .ZN(n2997) );
  NAND2_X1 U368 ( .A1(n2982), .A2(n2889), .ZN(n2995) );
  NAND2_X1 U369 ( .A1(n2982), .A2(n2886), .ZN(n2993) );
  NAND2_X1 U370 ( .A1(n2982), .A2(n2883), .ZN(n2991) );
  NAND2_X1 U371 ( .A1(n2982), .A2(n2880), .ZN(n2989) );
  NAND2_X1 U372 ( .A1(n2982), .A2(n2877), .ZN(n2987) );
  NAND2_X1 U373 ( .A1(n2982), .A2(n2874), .ZN(n2985) );
  NAND2_X1 U374 ( .A1(n2949), .A2(n2913), .ZN(n2978) );
  NAND2_X1 U375 ( .A1(n2949), .A2(n2910), .ZN(n2976) );
  NAND2_X1 U376 ( .A1(n2949), .A2(n2907), .ZN(n2974) );
  NAND2_X1 U377 ( .A1(n2949), .A2(n2904), .ZN(n2972) );
  NAND2_X1 U378 ( .A1(n2949), .A2(n2901), .ZN(n2970) );
  NAND2_X1 U379 ( .A1(n2949), .A2(n2898), .ZN(n2968) );
  NAND2_X1 U380 ( .A1(n2949), .A2(n2895), .ZN(n2966) );
  NAND2_X1 U381 ( .A1(n2949), .A2(n2889), .ZN(n2962) );
  NAND2_X1 U382 ( .A1(n2949), .A2(n2886), .ZN(n2960) );
  NAND2_X1 U383 ( .A1(n2949), .A2(n2883), .ZN(n2958) );
  NAND2_X1 U384 ( .A1(n2949), .A2(n2880), .ZN(n2956) );
  NAND2_X1 U385 ( .A1(n2949), .A2(n2877), .ZN(n2954) );
  NAND2_X1 U386 ( .A1(n2949), .A2(n2874), .ZN(n2952) );
  NAND2_X1 U387 ( .A1(n2949), .A2(n2871), .ZN(n2950) );
  NAND2_X1 U388 ( .A1(n2949), .A2(n2867), .ZN(n2947) );
  NAND2_X1 U389 ( .A1(n2916), .A2(n2904), .ZN(n2939) );
  NAND2_X1 U390 ( .A1(n2916), .A2(n2901), .ZN(n2937) );
  NAND2_X1 U391 ( .A1(n2916), .A2(n2898), .ZN(n2935) );
  NAND2_X1 U392 ( .A1(n2916), .A2(n2895), .ZN(n2933) );
  NAND2_X1 U393 ( .A1(n2916), .A2(n2892), .ZN(n2931) );
  NAND2_X1 U394 ( .A1(n2916), .A2(n2889), .ZN(n2929) );
  NAND2_X1 U395 ( .A1(n2916), .A2(n2883), .ZN(n2925) );
  NAND2_X1 U396 ( .A1(n2916), .A2(n2880), .ZN(n2923) );
  NAND2_X1 U397 ( .A1(n2916), .A2(n2877), .ZN(n2921) );
  NAND2_X1 U398 ( .A1(n2916), .A2(n2874), .ZN(n2919) );
  NAND2_X1 U399 ( .A1(n2916), .A2(n2871), .ZN(n2917) );
  NAND2_X1 U400 ( .A1(n2916), .A2(n2867), .ZN(n2914) );
  NAND2_X1 U401 ( .A1(n5710), .A2(n5664), .ZN(n4432) );
  NAND2_X1 U402 ( .A1(n4299), .A2(n4273), .ZN(n3149) );
  BUF_X1 U403 ( .A(n2961), .Z(n13583) );
  BUF_X1 U404 ( .A(n4354), .Z(n13093) );
  BUF_X1 U405 ( .A(n4354), .Z(n13094) );
  BUF_X1 U406 ( .A(n3070), .Z(n13321) );
  BUF_X1 U407 ( .A(n3070), .Z(n13322) );
  BUF_X1 U408 ( .A(n4343), .Z(n13120) );
  BUF_X1 U409 ( .A(n4369), .Z(n13066) );
  BUF_X1 U410 ( .A(n4380), .Z(n13039) );
  BUF_X1 U411 ( .A(n4406), .Z(n12985) );
  BUF_X1 U412 ( .A(n4421), .Z(n12958) );
  BUF_X1 U413 ( .A(n4343), .Z(n13121) );
  BUF_X1 U414 ( .A(n4369), .Z(n13067) );
  BUF_X1 U415 ( .A(n4380), .Z(n13040) );
  BUF_X1 U416 ( .A(n4406), .Z(n12986) );
  BUF_X1 U417 ( .A(n4421), .Z(n12959) );
  BUF_X1 U418 ( .A(n3059), .Z(n13348) );
  BUF_X1 U419 ( .A(n3085), .Z(n13294) );
  BUF_X1 U420 ( .A(n3096), .Z(n13267) );
  BUF_X1 U421 ( .A(n3122), .Z(n13213) );
  BUF_X1 U422 ( .A(n3137), .Z(n13186) );
  BUF_X1 U423 ( .A(n3148), .Z(n13159) );
  BUF_X1 U424 ( .A(n3059), .Z(n13349) );
  BUF_X1 U425 ( .A(n3085), .Z(n13295) );
  BUF_X1 U426 ( .A(n3096), .Z(n13268) );
  BUF_X1 U427 ( .A(n3122), .Z(n13214) );
  BUF_X1 U428 ( .A(n3137), .Z(n13187) );
  BUF_X1 U429 ( .A(n3148), .Z(n13160) );
  BUF_X1 U430 ( .A(n2834), .Z(n14010) );
  BUF_X1 U431 ( .A(n2876), .Z(n13792) );
  BUF_X1 U432 ( .A(n2876), .Z(n13793) );
  BUF_X1 U433 ( .A(n2894), .Z(n13756) );
  BUF_X1 U434 ( .A(n2903), .Z(n13738) );
  BUF_X1 U435 ( .A(n2903), .Z(n13739) );
  BUF_X1 U436 ( .A(n2879), .Z(n13786) );
  BUF_X1 U437 ( .A(n2879), .Z(n13787) );
  BUF_X1 U438 ( .A(n2834), .Z(n14011) );
  BUF_X1 U439 ( .A(n2906), .Z(n13732) );
  BUF_X1 U440 ( .A(n2906), .Z(n13733) );
  BUF_X1 U441 ( .A(n2926), .Z(n13684) );
  BUF_X1 U442 ( .A(n2926), .Z(n13685) );
  BUF_X1 U443 ( .A(n2928), .Z(n13678) );
  BUF_X1 U444 ( .A(n2928), .Z(n13679) );
  BUF_X1 U445 ( .A(n2942), .Z(n13637) );
  BUF_X1 U446 ( .A(n2944), .Z(n13630) );
  BUF_X1 U447 ( .A(n2944), .Z(n13631) );
  BUF_X1 U448 ( .A(n2946), .Z(n13624) );
  BUF_X1 U449 ( .A(n2946), .Z(n13625) );
  BUF_X1 U450 ( .A(n2961), .Z(n13582) );
  BUF_X1 U451 ( .A(n2963), .Z(n13576) );
  BUF_X1 U452 ( .A(n2963), .Z(n13577) );
  BUF_X1 U453 ( .A(n2965), .Z(n13570) );
  BUF_X1 U454 ( .A(n2965), .Z(n13571) );
  BUF_X1 U455 ( .A(n2975), .Z(n13540) );
  BUF_X1 U456 ( .A(n2975), .Z(n13541) );
  BUF_X1 U457 ( .A(n2984), .Z(n13517) );
  BUF_X1 U458 ( .A(n3030), .Z(n13402) );
  BUF_X1 U459 ( .A(n3030), .Z(n13403) );
  BUF_X1 U460 ( .A(n3028), .Z(n13408) );
  BUF_X1 U461 ( .A(n3028), .Z(n13409) );
  BUF_X1 U462 ( .A(n3018), .Z(n13432) );
  BUF_X1 U463 ( .A(n3018), .Z(n13433) );
  BUF_X1 U464 ( .A(n3005), .Z(n13462) );
  BUF_X1 U465 ( .A(n3005), .Z(n13463) );
  BUF_X1 U466 ( .A(n2986), .Z(n13510) );
  BUF_X1 U467 ( .A(n2986), .Z(n13511) );
  BUF_X1 U468 ( .A(n2984), .Z(n13516) );
  BUF_X1 U469 ( .A(n2948), .Z(n13618) );
  BUF_X1 U470 ( .A(n2948), .Z(n13619) );
  BUF_X1 U471 ( .A(n2942), .Z(n13636) );
  BUF_X1 U472 ( .A(n2930), .Z(n13672) );
  BUF_X1 U473 ( .A(n2930), .Z(n13673) );
  BUF_X1 U474 ( .A(n2924), .Z(n13690) );
  BUF_X1 U475 ( .A(n2924), .Z(n13691) );
  BUF_X1 U476 ( .A(n2909), .Z(n13726) );
  BUF_X1 U477 ( .A(n2909), .Z(n13727) );
  BUF_X1 U478 ( .A(n2897), .Z(n13750) );
  BUF_X1 U479 ( .A(n2897), .Z(n13751) );
  BUF_X1 U480 ( .A(n2894), .Z(n13757) );
  BUF_X1 U481 ( .A(n2882), .Z(n13780) );
  BUF_X1 U482 ( .A(n2882), .Z(n13781) );
  BUF_X1 U483 ( .A(n2870), .Z(n13804) );
  BUF_X1 U484 ( .A(n2870), .Z(n13805) );
  BUF_X1 U485 ( .A(n4355), .Z(n13090) );
  BUF_X1 U486 ( .A(n4355), .Z(n13091) );
  BUF_X1 U487 ( .A(n3071), .Z(n13318) );
  BUF_X1 U488 ( .A(n3071), .Z(n13319) );
  BUF_X1 U489 ( .A(n4396), .Z(n13009) );
  BUF_X1 U490 ( .A(n4396), .Z(n13010) );
  BUF_X1 U491 ( .A(n4344), .Z(n13117) );
  BUF_X1 U492 ( .A(n4370), .Z(n13063) );
  BUF_X1 U493 ( .A(n4381), .Z(n13036) );
  BUF_X1 U494 ( .A(n4407), .Z(n12982) );
  BUF_X1 U495 ( .A(n4422), .Z(n12955) );
  BUF_X1 U496 ( .A(n4433), .Z(n12928) );
  BUF_X1 U497 ( .A(n4344), .Z(n13118) );
  BUF_X1 U498 ( .A(n4370), .Z(n13064) );
  BUF_X1 U499 ( .A(n4381), .Z(n13037) );
  BUF_X1 U500 ( .A(n4407), .Z(n12983) );
  BUF_X1 U501 ( .A(n4422), .Z(n12956) );
  BUF_X1 U502 ( .A(n4433), .Z(n12929) );
  BUF_X1 U503 ( .A(n3060), .Z(n13345) );
  BUF_X1 U504 ( .A(n3086), .Z(n13291) );
  BUF_X1 U505 ( .A(n3097), .Z(n13264) );
  BUF_X1 U506 ( .A(n3112), .Z(n13237) );
  BUF_X1 U507 ( .A(n3123), .Z(n13210) );
  BUF_X1 U508 ( .A(n3138), .Z(n13183) );
  BUF_X1 U509 ( .A(n3060), .Z(n13346) );
  BUF_X1 U510 ( .A(n3086), .Z(n13292) );
  BUF_X1 U511 ( .A(n3097), .Z(n13265) );
  BUF_X1 U512 ( .A(n3112), .Z(n13238) );
  BUF_X1 U513 ( .A(n3123), .Z(n13211) );
  BUF_X1 U514 ( .A(n3138), .Z(n13184) );
  NAND2_X1 U515 ( .A1(n5661), .A2(n5664), .ZN(n4338) );
  NAND2_X1 U516 ( .A1(n5714), .A2(n5664), .ZN(n4395) );
  NAND2_X1 U517 ( .A1(n4272), .A2(n4273), .ZN(n3054) );
  NAND2_X1 U518 ( .A1(n4301), .A2(n4273), .ZN(n3111) );
  BUF_X1 U519 ( .A(n4345), .Z(n13114) );
  BUF_X1 U520 ( .A(n4351), .Z(n13099) );
  BUF_X1 U521 ( .A(n4345), .Z(n13115) );
  BUF_X1 U522 ( .A(n4351), .Z(n13100) );
  BUF_X1 U523 ( .A(n3061), .Z(n13342) );
  BUF_X1 U524 ( .A(n3067), .Z(n13327) );
  BUF_X1 U525 ( .A(n3061), .Z(n13343) );
  BUF_X1 U526 ( .A(n3067), .Z(n13328) );
  BUF_X1 U527 ( .A(n4334), .Z(n13141) );
  BUF_X1 U528 ( .A(n4340), .Z(n13126) );
  BUF_X1 U529 ( .A(n4360), .Z(n13087) );
  BUF_X1 U530 ( .A(n4366), .Z(n13072) );
  BUF_X1 U531 ( .A(n4377), .Z(n13045) );
  BUF_X1 U532 ( .A(n4386), .Z(n13033) );
  BUF_X1 U533 ( .A(n4397), .Z(n13006) );
  BUF_X1 U534 ( .A(n4392), .Z(n13018) );
  BUF_X1 U535 ( .A(n4403), .Z(n12991) );
  BUF_X1 U536 ( .A(n4412), .Z(n12979) );
  BUF_X1 U537 ( .A(n4423), .Z(n12952) );
  BUF_X1 U538 ( .A(n4418), .Z(n12964) );
  BUF_X1 U539 ( .A(n4429), .Z(n12937) );
  BUF_X1 U540 ( .A(n4334), .Z(n13142) );
  BUF_X1 U541 ( .A(n4340), .Z(n13127) );
  BUF_X1 U542 ( .A(n4360), .Z(n13088) );
  BUF_X1 U543 ( .A(n4366), .Z(n13073) );
  BUF_X1 U544 ( .A(n4377), .Z(n13046) );
  BUF_X1 U545 ( .A(n4386), .Z(n13034) );
  BUF_X1 U546 ( .A(n4397), .Z(n13007) );
  BUF_X1 U547 ( .A(n4392), .Z(n13019) );
  BUF_X1 U548 ( .A(n4403), .Z(n12992) );
  BUF_X1 U549 ( .A(n4412), .Z(n12980) );
  BUF_X1 U550 ( .A(n4423), .Z(n12953) );
  BUF_X1 U551 ( .A(n4418), .Z(n12965) );
  BUF_X1 U552 ( .A(n4429), .Z(n12938) );
  BUF_X1 U553 ( .A(n3050), .Z(n13369) );
  BUF_X1 U554 ( .A(n3056), .Z(n13354) );
  BUF_X1 U555 ( .A(n3076), .Z(n13315) );
  BUF_X1 U556 ( .A(n3082), .Z(n13300) );
  BUF_X1 U557 ( .A(n3093), .Z(n13273) );
  BUF_X1 U558 ( .A(n3102), .Z(n13261) );
  BUF_X1 U559 ( .A(n3113), .Z(n13234) );
  BUF_X1 U560 ( .A(n3108), .Z(n13246) );
  BUF_X1 U561 ( .A(n3119), .Z(n13219) );
  BUF_X1 U562 ( .A(n3128), .Z(n13207) );
  BUF_X1 U563 ( .A(n3139), .Z(n13180) );
  BUF_X1 U564 ( .A(n3134), .Z(n13192) );
  BUF_X1 U565 ( .A(n3145), .Z(n13165) );
  BUF_X1 U566 ( .A(n3050), .Z(n13370) );
  BUF_X1 U567 ( .A(n3056), .Z(n13355) );
  BUF_X1 U568 ( .A(n3076), .Z(n13316) );
  BUF_X1 U569 ( .A(n3082), .Z(n13301) );
  BUF_X1 U570 ( .A(n3093), .Z(n13274) );
  BUF_X1 U571 ( .A(n3102), .Z(n13262) );
  BUF_X1 U572 ( .A(n3113), .Z(n13235) );
  BUF_X1 U573 ( .A(n3108), .Z(n13247) );
  BUF_X1 U574 ( .A(n3119), .Z(n13220) );
  BUF_X1 U575 ( .A(n3128), .Z(n13208) );
  BUF_X1 U576 ( .A(n3139), .Z(n13181) );
  BUF_X1 U577 ( .A(n3134), .Z(n13193) );
  BUF_X1 U578 ( .A(n3145), .Z(n13166) );
  BUF_X1 U579 ( .A(n2981), .Z(n13522) );
  BUF_X1 U580 ( .A(n2981), .Z(n13523) );
  BUF_X1 U581 ( .A(n3035), .Z(n13390) );
  BUF_X1 U582 ( .A(n3035), .Z(n13391) );
  BUF_X1 U583 ( .A(n3033), .Z(n13396) );
  BUF_X1 U584 ( .A(n3033), .Z(n13397) );
  BUF_X1 U585 ( .A(n3026), .Z(n13414) );
  BUF_X1 U586 ( .A(n3026), .Z(n13415) );
  BUF_X1 U587 ( .A(n3024), .Z(n13420) );
  BUF_X1 U588 ( .A(n3024), .Z(n13421) );
  BUF_X1 U589 ( .A(n3020), .Z(n13426) );
  BUF_X1 U590 ( .A(n3020), .Z(n13427) );
  BUF_X1 U591 ( .A(n3016), .Z(n13438) );
  BUF_X1 U592 ( .A(n3016), .Z(n13439) );
  BUF_X1 U593 ( .A(n3014), .Z(n13444) );
  BUF_X1 U594 ( .A(n3014), .Z(n13445) );
  BUF_X1 U595 ( .A(n3011), .Z(n13450) );
  BUF_X1 U596 ( .A(n3011), .Z(n13451) );
  BUF_X1 U597 ( .A(n3008), .Z(n13456) );
  BUF_X1 U598 ( .A(n3008), .Z(n13457) );
  BUF_X1 U599 ( .A(n3002), .Z(n13468) );
  BUF_X1 U600 ( .A(n3002), .Z(n13469) );
  BUF_X1 U601 ( .A(n2998), .Z(n13474) );
  BUF_X1 U602 ( .A(n2998), .Z(n13475) );
  BUF_X1 U603 ( .A(n2996), .Z(n13480) );
  BUF_X1 U604 ( .A(n2996), .Z(n13481) );
  BUF_X1 U605 ( .A(n2994), .Z(n13486) );
  BUF_X1 U606 ( .A(n2994), .Z(n13487) );
  BUF_X1 U607 ( .A(n2992), .Z(n13492) );
  BUF_X1 U608 ( .A(n2992), .Z(n13493) );
  BUF_X1 U609 ( .A(n2990), .Z(n13498) );
  BUF_X1 U610 ( .A(n2990), .Z(n13499) );
  BUF_X1 U611 ( .A(n2988), .Z(n13504) );
  BUF_X1 U612 ( .A(n2988), .Z(n13505) );
  BUF_X1 U613 ( .A(n2979), .Z(n13528) );
  BUF_X1 U614 ( .A(n2979), .Z(n13529) );
  BUF_X1 U615 ( .A(n2977), .Z(n13534) );
  BUF_X1 U616 ( .A(n2977), .Z(n13535) );
  BUF_X1 U617 ( .A(n2973), .Z(n13546) );
  BUF_X1 U618 ( .A(n2973), .Z(n13547) );
  BUF_X1 U619 ( .A(n2971), .Z(n13552) );
  BUF_X1 U620 ( .A(n2971), .Z(n13553) );
  BUF_X1 U621 ( .A(n2969), .Z(n13558) );
  BUF_X1 U622 ( .A(n2969), .Z(n13559) );
  BUF_X1 U623 ( .A(n2967), .Z(n13564) );
  BUF_X1 U624 ( .A(n2967), .Z(n13565) );
  BUF_X1 U625 ( .A(n2959), .Z(n13588) );
  BUF_X1 U626 ( .A(n2959), .Z(n13589) );
  BUF_X1 U627 ( .A(n2957), .Z(n13594) );
  BUF_X1 U628 ( .A(n2957), .Z(n13595) );
  BUF_X1 U629 ( .A(n2955), .Z(n13600) );
  BUF_X1 U630 ( .A(n2955), .Z(n13601) );
  BUF_X1 U631 ( .A(n2953), .Z(n13606) );
  BUF_X1 U632 ( .A(n2953), .Z(n13607) );
  BUF_X1 U633 ( .A(n2951), .Z(n13612) );
  BUF_X1 U634 ( .A(n2951), .Z(n13613) );
  BUF_X1 U635 ( .A(n2940), .Z(n13642) );
  BUF_X1 U636 ( .A(n2940), .Z(n13643) );
  BUF_X1 U637 ( .A(n2938), .Z(n13648) );
  BUF_X1 U638 ( .A(n2938), .Z(n13649) );
  BUF_X1 U639 ( .A(n2936), .Z(n13654) );
  BUF_X1 U640 ( .A(n2936), .Z(n13655) );
  BUF_X1 U641 ( .A(n2934), .Z(n13660) );
  BUF_X1 U642 ( .A(n2934), .Z(n13661) );
  BUF_X1 U643 ( .A(n2932), .Z(n13666) );
  BUF_X1 U644 ( .A(n2932), .Z(n13667) );
  BUF_X1 U645 ( .A(n2922), .Z(n13696) );
  BUF_X1 U646 ( .A(n2922), .Z(n13697) );
  BUF_X1 U647 ( .A(n2920), .Z(n13702) );
  BUF_X1 U648 ( .A(n2920), .Z(n13703) );
  BUF_X1 U649 ( .A(n2918), .Z(n13708) );
  BUF_X1 U650 ( .A(n2918), .Z(n13709) );
  BUF_X1 U651 ( .A(n2915), .Z(n13714) );
  BUF_X1 U652 ( .A(n2915), .Z(n13715) );
  BUF_X1 U653 ( .A(n2912), .Z(n13720) );
  BUF_X1 U654 ( .A(n2912), .Z(n13721) );
  BUF_X1 U655 ( .A(n2900), .Z(n13744) );
  BUF_X1 U656 ( .A(n2900), .Z(n13745) );
  BUF_X1 U657 ( .A(n2891), .Z(n13762) );
  BUF_X1 U658 ( .A(n2891), .Z(n13763) );
  BUF_X1 U659 ( .A(n2888), .Z(n13768) );
  BUF_X1 U660 ( .A(n2888), .Z(n13769) );
  BUF_X1 U661 ( .A(n2885), .Z(n13774) );
  BUF_X1 U662 ( .A(n2885), .Z(n13775) );
  BUF_X1 U663 ( .A(n2873), .Z(n13798) );
  BUF_X1 U664 ( .A(n2873), .Z(n13799) );
  BUF_X1 U665 ( .A(n3036), .Z(n13387) );
  BUF_X1 U666 ( .A(n4346), .Z(n13111) );
  BUF_X1 U667 ( .A(n4352), .Z(n13096) );
  BUF_X1 U668 ( .A(n4346), .Z(n13112) );
  BUF_X1 U669 ( .A(n4352), .Z(n13097) );
  BUF_X1 U670 ( .A(n3062), .Z(n13339) );
  BUF_X1 U671 ( .A(n3068), .Z(n13324) );
  BUF_X1 U672 ( .A(n3062), .Z(n13340) );
  BUF_X1 U673 ( .A(n3068), .Z(n13325) );
  BUF_X1 U674 ( .A(n3036), .Z(n13388) );
  BUF_X1 U675 ( .A(n4335), .Z(n13138) );
  BUF_X1 U676 ( .A(n4341), .Z(n13123) );
  BUF_X1 U677 ( .A(n4372), .Z(n13057) );
  BUF_X1 U678 ( .A(n4367), .Z(n13069) );
  BUF_X1 U679 ( .A(n4378), .Z(n13042) );
  BUF_X1 U680 ( .A(n4387), .Z(n13030) );
  BUF_X1 U681 ( .A(n4398), .Z(n13003) );
  BUF_X1 U682 ( .A(n4393), .Z(n13015) );
  BUF_X1 U683 ( .A(n4413), .Z(n12976) );
  BUF_X1 U684 ( .A(n4424), .Z(n12949) );
  BUF_X1 U685 ( .A(n4430), .Z(n12934) );
  BUF_X1 U686 ( .A(n4335), .Z(n13139) );
  BUF_X1 U687 ( .A(n4341), .Z(n13124) );
  BUF_X1 U688 ( .A(n4372), .Z(n13058) );
  BUF_X1 U689 ( .A(n4367), .Z(n13070) );
  BUF_X1 U690 ( .A(n4378), .Z(n13043) );
  BUF_X1 U691 ( .A(n4387), .Z(n13031) );
  BUF_X1 U692 ( .A(n4398), .Z(n13004) );
  BUF_X1 U693 ( .A(n4393), .Z(n13016) );
  BUF_X1 U694 ( .A(n4413), .Z(n12977) );
  BUF_X1 U695 ( .A(n4424), .Z(n12950) );
  BUF_X1 U696 ( .A(n4430), .Z(n12935) );
  BUF_X1 U697 ( .A(n3051), .Z(n13366) );
  BUF_X1 U698 ( .A(n3057), .Z(n13351) );
  BUF_X1 U699 ( .A(n3088), .Z(n13285) );
  BUF_X1 U700 ( .A(n3083), .Z(n13297) );
  BUF_X1 U701 ( .A(n3094), .Z(n13270) );
  BUF_X1 U702 ( .A(n3103), .Z(n13258) );
  BUF_X1 U703 ( .A(n3114), .Z(n13231) );
  BUF_X1 U704 ( .A(n3109), .Z(n13243) );
  BUF_X1 U705 ( .A(n3129), .Z(n13204) );
  BUF_X1 U706 ( .A(n3140), .Z(n13177) );
  BUF_X1 U707 ( .A(n3146), .Z(n13162) );
  BUF_X1 U708 ( .A(n3051), .Z(n13367) );
  BUF_X1 U709 ( .A(n3057), .Z(n13352) );
  BUF_X1 U710 ( .A(n3088), .Z(n13286) );
  BUF_X1 U711 ( .A(n3083), .Z(n13298) );
  BUF_X1 U712 ( .A(n3094), .Z(n13271) );
  BUF_X1 U713 ( .A(n3103), .Z(n13259) );
  BUF_X1 U714 ( .A(n3114), .Z(n13232) );
  BUF_X1 U715 ( .A(n3109), .Z(n13244) );
  BUF_X1 U716 ( .A(n3129), .Z(n13205) );
  BUF_X1 U717 ( .A(n3140), .Z(n13178) );
  BUF_X1 U718 ( .A(n3146), .Z(n13163) );
  BUF_X1 U719 ( .A(n4339), .Z(n13129) );
  BUF_X1 U720 ( .A(n4339), .Z(n13130) );
  BUF_X1 U721 ( .A(n4365), .Z(n13075) );
  BUF_X1 U722 ( .A(n4376), .Z(n13048) );
  BUF_X1 U723 ( .A(n4391), .Z(n13021) );
  BUF_X1 U724 ( .A(n4402), .Z(n12994) );
  BUF_X1 U725 ( .A(n4417), .Z(n12967) );
  BUF_X1 U726 ( .A(n4428), .Z(n12940) );
  BUF_X1 U727 ( .A(n4365), .Z(n13076) );
  BUF_X1 U728 ( .A(n4376), .Z(n13049) );
  BUF_X1 U729 ( .A(n4391), .Z(n13022) );
  BUF_X1 U730 ( .A(n4402), .Z(n12995) );
  BUF_X1 U731 ( .A(n4417), .Z(n12968) );
  BUF_X1 U732 ( .A(n4428), .Z(n12941) );
  BUF_X1 U733 ( .A(n3055), .Z(n13357) );
  BUF_X1 U734 ( .A(n3081), .Z(n13303) );
  BUF_X1 U735 ( .A(n3092), .Z(n13276) );
  BUF_X1 U736 ( .A(n3107), .Z(n13249) );
  BUF_X1 U737 ( .A(n3118), .Z(n13222) );
  BUF_X1 U738 ( .A(n3133), .Z(n13195) );
  BUF_X1 U739 ( .A(n3144), .Z(n13168) );
  BUF_X1 U740 ( .A(n3055), .Z(n13358) );
  BUF_X1 U741 ( .A(n3081), .Z(n13304) );
  BUF_X1 U742 ( .A(n3092), .Z(n13277) );
  BUF_X1 U743 ( .A(n3107), .Z(n13250) );
  BUF_X1 U744 ( .A(n3118), .Z(n13223) );
  BUF_X1 U745 ( .A(n3133), .Z(n13196) );
  BUF_X1 U746 ( .A(n3144), .Z(n13169) );
  BUF_X1 U747 ( .A(n4354), .Z(n13095) );
  BUF_X1 U748 ( .A(n3070), .Z(n13323) );
  BUF_X1 U749 ( .A(n4343), .Z(n13122) );
  BUF_X1 U750 ( .A(n4369), .Z(n13068) );
  BUF_X1 U751 ( .A(n4380), .Z(n13041) );
  BUF_X1 U752 ( .A(n4406), .Z(n12987) );
  BUF_X1 U753 ( .A(n4421), .Z(n12960) );
  BUF_X1 U754 ( .A(n3059), .Z(n13350) );
  BUF_X1 U755 ( .A(n3085), .Z(n13296) );
  BUF_X1 U756 ( .A(n3096), .Z(n13269) );
  BUF_X1 U757 ( .A(n3137), .Z(n13188) );
  BUF_X1 U758 ( .A(n3148), .Z(n13161) );
  BUF_X1 U759 ( .A(n3122), .Z(n13215) );
  NAND2_X1 U760 ( .A1(n2877), .A2(n2868), .ZN(n2875) );
  NAND2_X1 U761 ( .A1(n2904), .A2(n2868), .ZN(n2902) );
  NAND2_X1 U762 ( .A1(n2880), .A2(n2868), .ZN(n2878) );
  NAND2_X1 U763 ( .A1(n2907), .A2(n2868), .ZN(n2905) );
  NAND2_X1 U764 ( .A1(n2913), .A2(n2868), .ZN(n2911) );
  NAND2_X1 U765 ( .A1(n2910), .A2(n2868), .ZN(n2908) );
  NAND2_X1 U766 ( .A1(n2901), .A2(n2868), .ZN(n2899) );
  NAND2_X1 U767 ( .A1(n2898), .A2(n2868), .ZN(n2896) );
  NAND2_X1 U768 ( .A1(n2895), .A2(n2868), .ZN(n2893) );
  NAND2_X1 U769 ( .A1(n2892), .A2(n2868), .ZN(n2890) );
  NAND2_X1 U770 ( .A1(n2889), .A2(n2868), .ZN(n2887) );
  NAND2_X1 U771 ( .A1(n2886), .A2(n2868), .ZN(n2884) );
  NAND2_X1 U772 ( .A1(n2883), .A2(n2868), .ZN(n2881) );
  NAND2_X1 U773 ( .A1(n2874), .A2(n2868), .ZN(n2872) );
  NAND2_X1 U774 ( .A1(n2871), .A2(n2868), .ZN(n2869) );
  NAND2_X1 U775 ( .A1(n2867), .A2(n2868), .ZN(n2832) );
  BUF_X1 U776 ( .A(n3030), .Z(n13404) );
  BUF_X1 U777 ( .A(n3028), .Z(n13410) );
  BUF_X1 U778 ( .A(n2834), .Z(n14012) );
  BUF_X1 U779 ( .A(n2876), .Z(n13794) );
  BUF_X1 U780 ( .A(n2903), .Z(n13740) );
  BUF_X1 U781 ( .A(n2924), .Z(n13692) );
  BUF_X1 U782 ( .A(n2942), .Z(n13638) );
  BUF_X1 U783 ( .A(n2984), .Z(n13518) );
  BUF_X1 U784 ( .A(n2879), .Z(n13788) );
  BUF_X1 U785 ( .A(n2906), .Z(n13734) );
  BUF_X1 U786 ( .A(n2928), .Z(n13680) );
  BUF_X1 U787 ( .A(n2944), .Z(n13632) );
  BUF_X1 U788 ( .A(n2946), .Z(n13626) );
  BUF_X1 U789 ( .A(n2965), .Z(n13572) );
  BUF_X1 U790 ( .A(n3018), .Z(n13434) );
  BUF_X1 U791 ( .A(n3005), .Z(n13464) );
  BUF_X1 U792 ( .A(n2986), .Z(n13512) );
  BUF_X1 U793 ( .A(n2975), .Z(n13542) );
  BUF_X1 U794 ( .A(n2948), .Z(n13620) );
  BUF_X1 U795 ( .A(n2930), .Z(n13674) );
  BUF_X1 U796 ( .A(n2909), .Z(n13728) );
  BUF_X1 U797 ( .A(n2897), .Z(n13752) );
  BUF_X1 U798 ( .A(n2894), .Z(n13758) );
  BUF_X1 U799 ( .A(n2882), .Z(n13782) );
  BUF_X1 U800 ( .A(n2870), .Z(n13806) );
  BUF_X1 U801 ( .A(n4348), .Z(n13108) );
  BUF_X1 U802 ( .A(n4348), .Z(n13109) );
  BUF_X1 U803 ( .A(n4337), .Z(n13135) );
  BUF_X1 U804 ( .A(n4363), .Z(n13081) );
  BUF_X1 U805 ( .A(n4374), .Z(n13054) );
  BUF_X1 U806 ( .A(n4389), .Z(n13027) );
  BUF_X1 U807 ( .A(n4400), .Z(n13000) );
  BUF_X1 U808 ( .A(n4415), .Z(n12973) );
  BUF_X1 U809 ( .A(n4426), .Z(n12946) );
  BUF_X1 U810 ( .A(n4337), .Z(n13136) );
  BUF_X1 U811 ( .A(n4363), .Z(n13082) );
  BUF_X1 U812 ( .A(n4374), .Z(n13055) );
  BUF_X1 U813 ( .A(n4389), .Z(n13028) );
  BUF_X1 U814 ( .A(n4400), .Z(n13001) );
  BUF_X1 U815 ( .A(n4415), .Z(n12974) );
  BUF_X1 U816 ( .A(n4426), .Z(n12947) );
  BUF_X1 U817 ( .A(n3053), .Z(n13363) );
  BUF_X1 U818 ( .A(n3064), .Z(n13336) );
  BUF_X1 U819 ( .A(n3079), .Z(n13309) );
  BUF_X1 U820 ( .A(n3090), .Z(n13282) );
  BUF_X1 U821 ( .A(n3105), .Z(n13255) );
  BUF_X1 U822 ( .A(n3116), .Z(n13228) );
  BUF_X1 U823 ( .A(n3131), .Z(n13201) );
  BUF_X1 U824 ( .A(n3142), .Z(n13174) );
  BUF_X1 U825 ( .A(n3053), .Z(n13364) );
  BUF_X1 U826 ( .A(n3064), .Z(n13337) );
  BUF_X1 U827 ( .A(n3079), .Z(n13310) );
  BUF_X1 U828 ( .A(n3090), .Z(n13283) );
  BUF_X1 U829 ( .A(n3105), .Z(n13256) );
  BUF_X1 U830 ( .A(n3116), .Z(n13229) );
  BUF_X1 U831 ( .A(n3131), .Z(n13202) );
  BUF_X1 U832 ( .A(n3142), .Z(n13175) );
  BUF_X1 U833 ( .A(n4349), .Z(n13105) );
  BUF_X1 U834 ( .A(n4349), .Z(n13106) );
  BUF_X1 U835 ( .A(n3065), .Z(n13333) );
  BUF_X1 U836 ( .A(n3065), .Z(n13334) );
  BUF_X1 U837 ( .A(n4375), .Z(n13051) );
  BUF_X1 U838 ( .A(n4375), .Z(n13052) );
  BUF_X1 U839 ( .A(n4364), .Z(n13078) );
  BUF_X1 U840 ( .A(n4390), .Z(n13024) );
  BUF_X1 U841 ( .A(n4401), .Z(n12997) );
  BUF_X1 U842 ( .A(n4416), .Z(n12970) );
  BUF_X1 U843 ( .A(n4427), .Z(n12943) );
  BUF_X1 U844 ( .A(n4364), .Z(n13079) );
  BUF_X1 U845 ( .A(n4390), .Z(n13025) );
  BUF_X1 U846 ( .A(n4401), .Z(n12998) );
  BUF_X1 U847 ( .A(n4416), .Z(n12971) );
  BUF_X1 U848 ( .A(n4427), .Z(n12944) );
  BUF_X1 U849 ( .A(n3080), .Z(n13306) );
  BUF_X1 U850 ( .A(n3091), .Z(n13279) );
  BUF_X1 U851 ( .A(n3106), .Z(n13252) );
  BUF_X1 U852 ( .A(n3117), .Z(n13225) );
  BUF_X1 U853 ( .A(n3132), .Z(n13198) );
  BUF_X1 U854 ( .A(n3143), .Z(n13171) );
  BUF_X1 U855 ( .A(n3080), .Z(n13307) );
  BUF_X1 U856 ( .A(n3091), .Z(n13280) );
  BUF_X1 U857 ( .A(n3106), .Z(n13253) );
  BUF_X1 U858 ( .A(n3117), .Z(n13226) );
  BUF_X1 U859 ( .A(n3132), .Z(n13199) );
  BUF_X1 U860 ( .A(n3143), .Z(n13172) );
  BUF_X1 U861 ( .A(n4355), .Z(n13092) );
  BUF_X1 U862 ( .A(n3071), .Z(n13320) );
  BUF_X1 U863 ( .A(n2963), .Z(n13578) );
  BUF_X1 U864 ( .A(n4396), .Z(n13011) );
  BUF_X1 U865 ( .A(n4344), .Z(n13119) );
  BUF_X1 U866 ( .A(n4370), .Z(n13065) );
  BUF_X1 U867 ( .A(n4381), .Z(n13038) );
  BUF_X1 U868 ( .A(n4407), .Z(n12984) );
  BUF_X1 U869 ( .A(n4422), .Z(n12957) );
  BUF_X1 U870 ( .A(n4433), .Z(n12930) );
  BUF_X1 U871 ( .A(n3060), .Z(n13347) );
  BUF_X1 U872 ( .A(n3086), .Z(n13293) );
  BUF_X1 U873 ( .A(n3097), .Z(n13266) );
  BUF_X1 U874 ( .A(n3138), .Z(n13185) );
  BUF_X1 U875 ( .A(n3112), .Z(n13239) );
  BUF_X1 U876 ( .A(n3123), .Z(n13212) );
  BUF_X1 U877 ( .A(n2926), .Z(n13686) );
  BUF_X1 U878 ( .A(n4345), .Z(n13116) );
  BUF_X1 U879 ( .A(n4351), .Z(n13101) );
  BUF_X1 U880 ( .A(n3061), .Z(n13344) );
  BUF_X1 U881 ( .A(n3067), .Z(n13329) );
  BUF_X1 U882 ( .A(n4418), .Z(n12966) );
  BUF_X1 U883 ( .A(n4334), .Z(n13143) );
  BUF_X1 U884 ( .A(n4340), .Z(n13128) );
  BUF_X1 U885 ( .A(n4360), .Z(n13089) );
  BUF_X1 U886 ( .A(n4366), .Z(n13074) );
  BUF_X1 U887 ( .A(n4377), .Z(n13047) );
  BUF_X1 U888 ( .A(n4386), .Z(n13035) );
  BUF_X1 U889 ( .A(n4397), .Z(n13008) );
  BUF_X1 U890 ( .A(n4392), .Z(n13020) );
  BUF_X1 U891 ( .A(n4403), .Z(n12993) );
  BUF_X1 U892 ( .A(n4423), .Z(n12954) );
  BUF_X1 U893 ( .A(n4429), .Z(n12939) );
  BUF_X1 U894 ( .A(n3050), .Z(n13371) );
  BUF_X1 U895 ( .A(n3056), .Z(n13356) );
  BUF_X1 U896 ( .A(n3076), .Z(n13317) );
  BUF_X1 U897 ( .A(n3082), .Z(n13302) );
  BUF_X1 U898 ( .A(n3093), .Z(n13275) );
  BUF_X1 U899 ( .A(n3102), .Z(n13263) );
  BUF_X1 U900 ( .A(n3113), .Z(n13236) );
  BUF_X1 U901 ( .A(n3108), .Z(n13248) );
  BUF_X1 U902 ( .A(n3119), .Z(n13221) );
  BUF_X1 U903 ( .A(n4412), .Z(n12981) );
  BUF_X1 U904 ( .A(n3128), .Z(n13209) );
  BUF_X1 U905 ( .A(n3139), .Z(n13182) );
  BUF_X1 U906 ( .A(n3134), .Z(n13194) );
  BUF_X1 U907 ( .A(n3145), .Z(n13167) );
  BUF_X1 U908 ( .A(n3035), .Z(n13392) );
  BUF_X1 U909 ( .A(n3033), .Z(n13398) );
  BUF_X1 U910 ( .A(n3026), .Z(n13416) );
  BUF_X1 U911 ( .A(n3024), .Z(n13422) );
  BUF_X1 U912 ( .A(n2981), .Z(n13524) );
  BUF_X1 U913 ( .A(n3020), .Z(n13428) );
  BUF_X1 U914 ( .A(n3016), .Z(n13440) );
  BUF_X1 U915 ( .A(n3014), .Z(n13446) );
  BUF_X1 U916 ( .A(n3011), .Z(n13452) );
  BUF_X1 U917 ( .A(n3008), .Z(n13458) );
  BUF_X1 U918 ( .A(n3002), .Z(n13470) );
  BUF_X1 U919 ( .A(n2998), .Z(n13476) );
  BUF_X1 U920 ( .A(n2996), .Z(n13482) );
  BUF_X1 U921 ( .A(n2994), .Z(n13488) );
  BUF_X1 U922 ( .A(n2992), .Z(n13494) );
  BUF_X1 U923 ( .A(n2990), .Z(n13500) );
  BUF_X1 U924 ( .A(n2988), .Z(n13506) );
  BUF_X1 U925 ( .A(n2979), .Z(n13530) );
  BUF_X1 U926 ( .A(n2977), .Z(n13536) );
  BUF_X1 U927 ( .A(n2973), .Z(n13548) );
  BUF_X1 U928 ( .A(n2971), .Z(n13554) );
  BUF_X1 U929 ( .A(n2969), .Z(n13560) );
  BUF_X1 U930 ( .A(n2967), .Z(n13566) );
  BUF_X1 U931 ( .A(n2959), .Z(n13590) );
  BUF_X1 U932 ( .A(n2957), .Z(n13596) );
  BUF_X1 U933 ( .A(n2955), .Z(n13602) );
  BUF_X1 U934 ( .A(n2953), .Z(n13608) );
  BUF_X1 U935 ( .A(n2951), .Z(n13614) );
  BUF_X1 U936 ( .A(n2940), .Z(n13644) );
  BUF_X1 U937 ( .A(n2938), .Z(n13650) );
  BUF_X1 U938 ( .A(n2936), .Z(n13656) );
  BUF_X1 U939 ( .A(n2934), .Z(n13662) );
  BUF_X1 U940 ( .A(n2932), .Z(n13668) );
  BUF_X1 U941 ( .A(n2922), .Z(n13698) );
  BUF_X1 U942 ( .A(n2920), .Z(n13704) );
  BUF_X1 U943 ( .A(n2918), .Z(n13710) );
  BUF_X1 U944 ( .A(n2915), .Z(n13716) );
  BUF_X1 U945 ( .A(n2912), .Z(n13722) );
  BUF_X1 U946 ( .A(n2900), .Z(n13746) );
  BUF_X1 U947 ( .A(n2891), .Z(n13764) );
  BUF_X1 U948 ( .A(n2888), .Z(n13770) );
  BUF_X1 U949 ( .A(n2885), .Z(n13776) );
  BUF_X1 U950 ( .A(n2873), .Z(n13800) );
  BUF_X1 U951 ( .A(n3036), .Z(n13389) );
  BUF_X1 U952 ( .A(n4346), .Z(n13113) );
  BUF_X1 U953 ( .A(n4352), .Z(n13098) );
  BUF_X1 U954 ( .A(n3062), .Z(n13341) );
  BUF_X1 U955 ( .A(n3068), .Z(n13326) );
  BUF_X1 U956 ( .A(n4335), .Z(n13140) );
  BUF_X1 U957 ( .A(n4341), .Z(n13125) );
  BUF_X1 U958 ( .A(n4372), .Z(n13059) );
  BUF_X1 U959 ( .A(n4367), .Z(n13071) );
  BUF_X1 U960 ( .A(n4378), .Z(n13044) );
  BUF_X1 U961 ( .A(n4387), .Z(n13032) );
  BUF_X1 U962 ( .A(n4398), .Z(n13005) );
  BUF_X1 U963 ( .A(n4393), .Z(n13017) );
  BUF_X1 U964 ( .A(n4424), .Z(n12951) );
  BUF_X1 U965 ( .A(n4430), .Z(n12936) );
  BUF_X1 U966 ( .A(n3051), .Z(n13368) );
  BUF_X1 U967 ( .A(n3057), .Z(n13353) );
  BUF_X1 U968 ( .A(n3088), .Z(n13287) );
  BUF_X1 U969 ( .A(n3083), .Z(n13299) );
  BUF_X1 U970 ( .A(n3094), .Z(n13272) );
  BUF_X1 U971 ( .A(n3103), .Z(n13260) );
  BUF_X1 U972 ( .A(n3114), .Z(n13233) );
  BUF_X1 U973 ( .A(n3109), .Z(n13245) );
  BUF_X1 U974 ( .A(n4413), .Z(n12978) );
  BUF_X1 U975 ( .A(n3129), .Z(n13206) );
  BUF_X1 U976 ( .A(n3140), .Z(n13179) );
  BUF_X1 U977 ( .A(n3146), .Z(n13164) );
  AND2_X1 U978 ( .A1(n3031), .A2(n3009), .ZN(n2889) );
  BUF_X1 U979 ( .A(n4339), .Z(n13131) );
  BUF_X1 U980 ( .A(n4376), .Z(n13050) );
  BUF_X1 U981 ( .A(n3133), .Z(n13197) );
  BUF_X1 U982 ( .A(n4365), .Z(n13077) );
  BUF_X1 U983 ( .A(n4391), .Z(n13023) );
  BUF_X1 U984 ( .A(n4402), .Z(n12996) );
  BUF_X1 U985 ( .A(n4417), .Z(n12969) );
  BUF_X1 U986 ( .A(n4428), .Z(n12942) );
  BUF_X1 U987 ( .A(n3055), .Z(n13359) );
  BUF_X1 U988 ( .A(n3092), .Z(n13278) );
  BUF_X1 U989 ( .A(n3081), .Z(n13305) );
  BUF_X1 U990 ( .A(n3107), .Z(n13251) );
  BUF_X1 U991 ( .A(n3118), .Z(n13224) );
  BUF_X1 U992 ( .A(n3144), .Z(n13170) );
  BUF_X1 U993 ( .A(n4349), .Z(n13107) );
  BUF_X1 U994 ( .A(n3065), .Z(n13335) );
  BUF_X1 U995 ( .A(n4348), .Z(n13110) );
  BUF_X1 U996 ( .A(n4337), .Z(n13137) );
  BUF_X1 U997 ( .A(n4374), .Z(n13056) );
  BUF_X1 U998 ( .A(n4415), .Z(n12975) );
  BUF_X1 U999 ( .A(n4426), .Z(n12948) );
  BUF_X1 U1000 ( .A(n3053), .Z(n13365) );
  BUF_X1 U1001 ( .A(n3090), .Z(n13284) );
  BUF_X1 U1002 ( .A(n3131), .Z(n13203) );
  BUF_X1 U1003 ( .A(n3142), .Z(n13176) );
  BUF_X1 U1004 ( .A(n4363), .Z(n13083) );
  BUF_X1 U1005 ( .A(n4389), .Z(n13029) );
  BUF_X1 U1006 ( .A(n4400), .Z(n13002) );
  BUF_X1 U1007 ( .A(n3064), .Z(n13338) );
  BUF_X1 U1008 ( .A(n3079), .Z(n13311) );
  BUF_X1 U1009 ( .A(n3105), .Z(n13257) );
  BUF_X1 U1010 ( .A(n3116), .Z(n13230) );
  BUF_X1 U1011 ( .A(n4375), .Z(n13053) );
  BUF_X1 U1012 ( .A(n4416), .Z(n12972) );
  BUF_X1 U1013 ( .A(n3080), .Z(n13308) );
  BUF_X1 U1014 ( .A(n3091), .Z(n13281) );
  BUF_X1 U1015 ( .A(n3132), .Z(n13200) );
  BUF_X1 U1016 ( .A(n4364), .Z(n13080) );
  BUF_X1 U1017 ( .A(n4390), .Z(n13026) );
  BUF_X1 U1018 ( .A(n4401), .Z(n12999) );
  BUF_X1 U1019 ( .A(n4427), .Z(n12945) );
  BUF_X1 U1020 ( .A(n3106), .Z(n13254) );
  BUF_X1 U1021 ( .A(n3117), .Z(n13227) );
  BUF_X1 U1022 ( .A(n3143), .Z(n13173) );
  BUF_X1 U1023 ( .A(n2961), .Z(n13584) );
  AND2_X1 U1024 ( .A1(n2999), .A2(n3009), .ZN(n2901) );
  NAND2_X1 U1025 ( .A1(n13149), .A2(n13153), .ZN(n4324) );
  NAND2_X1 U1026 ( .A1(n13377), .A2(n13381), .ZN(n3040) );
  NAND2_X1 U1027 ( .A1(n3021), .A2(n2889), .ZN(n3037) );
  NAND2_X1 U1028 ( .A1(n3021), .A2(n2886), .ZN(n3034) );
  NAND2_X1 U1029 ( .A1(n3021), .A2(n2883), .ZN(n3032) );
  NAND2_X1 U1030 ( .A1(n3021), .A2(n2880), .ZN(n3029) );
  NAND2_X1 U1031 ( .A1(n3021), .A2(n2877), .ZN(n3027) );
  NAND2_X1 U1032 ( .A1(n3021), .A2(n2874), .ZN(n3025) );
  NAND2_X1 U1033 ( .A1(n3021), .A2(n2871), .ZN(n3023) );
  NAND2_X1 U1034 ( .A1(n3021), .A2(n2867), .ZN(n3019) );
  AND2_X1 U1035 ( .A1(n5691), .A2(n5664), .ZN(n4361) );
  AND2_X1 U1036 ( .A1(n5690), .A2(n5664), .ZN(n4404) );
  AND2_X1 U1037 ( .A1(n4290), .A2(n4273), .ZN(n3077) );
  AND2_X1 U1038 ( .A1(n4289), .A2(n4273), .ZN(n3120) );
  AND2_X1 U1039 ( .A1(n5659), .A2(n5664), .ZN(n4371) );
  AND2_X1 U1040 ( .A1(n4270), .A2(n4273), .ZN(n3087) );
  AND2_X1 U1041 ( .A1(n5732), .A2(n5664), .ZN(n4419) );
  AND2_X1 U1042 ( .A1(n4310), .A2(n4273), .ZN(n3135) );
  NOR3_X1 U1043 ( .A1(n16062), .A2(ADD_RD2[5]), .A3(n16058), .ZN(n5691) );
  NOR3_X1 U1044 ( .A1(n16061), .A2(ADD_RD1[5]), .A3(n16056), .ZN(n4290) );
  NOR3_X1 U1045 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n16057), .ZN(n5690) );
  NOR3_X1 U1046 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n16055), .ZN(n4289) );
  NOR3_X1 U1047 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[5]), .A3(n16062), .ZN(n5661) );
  NOR3_X1 U1048 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[5]), .A3(n16061), .ZN(n4272) );
  NOR3_X1 U1049 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[5]), .A3(n16058), .ZN(n5659) );
  NOR3_X1 U1050 ( .A1(n16062), .A2(ADD_RD2[4]), .A3(n16057), .ZN(n5714) );
  NOR3_X1 U1051 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[5]), .A3(n16056), .ZN(n4270) );
  NOR3_X1 U1052 ( .A1(n16061), .A2(ADD_RD1[4]), .A3(n16055), .ZN(n4301) );
  NOR3_X2 U1053 ( .A1(n16068), .A2(n16067), .A3(n16069), .ZN(n5664) );
  NOR3_X2 U1054 ( .A1(n16065), .A2(n16064), .A3(n16066), .ZN(n4273) );
  NOR4_X1 U1055 ( .A1(n5746), .A2(n5748), .A3(n5750), .A4(n5752), .ZN(n5744)
         );
  NOR4_X1 U1056 ( .A1(n4317), .A2(n4318), .A3(n4319), .A4(n4320), .ZN(n4316)
         );
  AND3_X1 U1057 ( .A1(n16060), .A2(n16059), .A3(ADD_WR[6]), .ZN(n3021) );
  NAND2_X1 U1058 ( .A1(n5679), .A2(n5669), .ZN(n4349) );
  NAND2_X1 U1059 ( .A1(n5679), .A2(n5666), .ZN(n4354) );
  NAND2_X1 U1060 ( .A1(n5679), .A2(n5660), .ZN(n4355) );
  NAND2_X1 U1061 ( .A1(n4282), .A2(n4276), .ZN(n3065) );
  NAND2_X1 U1062 ( .A1(n4282), .A2(n4280), .ZN(n3070) );
  NAND2_X1 U1063 ( .A1(n4282), .A2(n4279), .ZN(n3071) );
  OAI21_X1 U1064 ( .B1(n14021), .B2(n13810), .A(n12927), .ZN(n2834) );
  OAI21_X1 U1065 ( .B1(n2866), .B2(n13386), .A(n12922), .ZN(n3036) );
  OAI21_X1 U1066 ( .B1(n13810), .B2(n13395), .A(n12922), .ZN(n3035) );
  OAI21_X1 U1067 ( .B1(n2866), .B2(n13401), .A(n12922), .ZN(n3033) );
  OAI21_X1 U1068 ( .B1(n13810), .B2(n13407), .A(n12922), .ZN(n3030) );
  OAI21_X1 U1069 ( .B1(n2866), .B2(n13413), .A(n12922), .ZN(n3028) );
  OAI21_X1 U1070 ( .B1(n13810), .B2(n13419), .A(n12922), .ZN(n3026) );
  OAI21_X1 U1071 ( .B1(n2866), .B2(n13425), .A(n12922), .ZN(n3024) );
  OAI21_X1 U1072 ( .B1(n13810), .B2(n13797), .A(n12927), .ZN(n2876) );
  OAI21_X1 U1073 ( .B1(n2866), .B2(n13743), .A(n12926), .ZN(n2903) );
  OAI21_X1 U1074 ( .B1(n13810), .B2(n13791), .A(n12927), .ZN(n2879) );
  OAI21_X1 U1075 ( .B1(n2866), .B2(n13749), .A(n12927), .ZN(n2900) );
  OAI21_X1 U1076 ( .B1(n13810), .B2(n13755), .A(n12927), .ZN(n2897) );
  OAI21_X1 U1077 ( .B1(n2866), .B2(n13761), .A(n12927), .ZN(n2894) );
  OAI21_X1 U1078 ( .B1(n13810), .B2(n13767), .A(n12927), .ZN(n2891) );
  OAI21_X1 U1079 ( .B1(n2866), .B2(n13773), .A(n12927), .ZN(n2888) );
  OAI21_X1 U1080 ( .B1(n13810), .B2(n13779), .A(n12927), .ZN(n2885) );
  OAI21_X1 U1081 ( .B1(n2866), .B2(n13785), .A(n12927), .ZN(n2882) );
  OAI21_X1 U1082 ( .B1(n13810), .B2(n13803), .A(n12927), .ZN(n2873) );
  OAI21_X1 U1083 ( .B1(n2866), .B2(n13809), .A(n12927), .ZN(n2870) );
  OAI21_X1 U1084 ( .B1(n13812), .B2(n13527), .A(n12923), .ZN(n2981) );
  OAI21_X1 U1085 ( .B1(n2866), .B2(n13737), .A(n12926), .ZN(n2906) );
  OAI21_X1 U1086 ( .B1(n13810), .B2(n13683), .A(n12926), .ZN(n2928) );
  OAI21_X1 U1087 ( .B1(n13811), .B2(n13635), .A(n12925), .ZN(n2944) );
  OAI21_X1 U1088 ( .B1(n13811), .B2(n13629), .A(n12925), .ZN(n2946) );
  OAI21_X1 U1089 ( .B1(n13812), .B2(n13575), .A(n12924), .ZN(n2965) );
  OAI21_X1 U1090 ( .B1(n13813), .B2(n13431), .A(n12922), .ZN(n3020) );
  OAI21_X1 U1091 ( .B1(n13813), .B2(n13437), .A(n12922), .ZN(n3018) );
  OAI21_X1 U1092 ( .B1(n13813), .B2(n13443), .A(n12922), .ZN(n3016) );
  OAI21_X1 U1093 ( .B1(n13813), .B2(n13449), .A(n12922), .ZN(n3014) );
  OAI21_X1 U1094 ( .B1(n13813), .B2(n13455), .A(n12922), .ZN(n3011) );
  OAI21_X1 U1095 ( .B1(n13813), .B2(n13461), .A(n12923), .ZN(n3008) );
  OAI21_X1 U1096 ( .B1(n13813), .B2(n13467), .A(n12923), .ZN(n3005) );
  OAI21_X1 U1097 ( .B1(n13813), .B2(n13473), .A(n12923), .ZN(n3002) );
  OAI21_X1 U1098 ( .B1(n13813), .B2(n13479), .A(n12923), .ZN(n2998) );
  OAI21_X1 U1099 ( .B1(n13813), .B2(n13485), .A(n12923), .ZN(n2996) );
  OAI21_X1 U1100 ( .B1(n13813), .B2(n13491), .A(n12923), .ZN(n2994) );
  OAI21_X1 U1101 ( .B1(n13813), .B2(n13497), .A(n12923), .ZN(n2992) );
  OAI21_X1 U1102 ( .B1(n13813), .B2(n13503), .A(n12923), .ZN(n2990) );
  OAI21_X1 U1103 ( .B1(n13812), .B2(n13509), .A(n12923), .ZN(n2988) );
  OAI21_X1 U1104 ( .B1(n13812), .B2(n13515), .A(n12923), .ZN(n2986) );
  OAI21_X1 U1105 ( .B1(n13812), .B2(n13521), .A(n12923), .ZN(n2984) );
  OAI21_X1 U1106 ( .B1(n13812), .B2(n13533), .A(n12924), .ZN(n2979) );
  OAI21_X1 U1107 ( .B1(n13812), .B2(n13539), .A(n12924), .ZN(n2977) );
  OAI21_X1 U1108 ( .B1(n13812), .B2(n13545), .A(n12924), .ZN(n2975) );
  OAI21_X1 U1109 ( .B1(n13812), .B2(n13551), .A(n12924), .ZN(n2973) );
  OAI21_X1 U1110 ( .B1(n13812), .B2(n13557), .A(n12924), .ZN(n2971) );
  OAI21_X1 U1111 ( .B1(n13812), .B2(n13563), .A(n12924), .ZN(n2969) );
  OAI21_X1 U1112 ( .B1(n13812), .B2(n13569), .A(n12924), .ZN(n2967) );
  OAI21_X1 U1113 ( .B1(n13812), .B2(n13581), .A(n12924), .ZN(n2963) );
  OAI21_X1 U1114 ( .B1(n13811), .B2(n13587), .A(n12924), .ZN(n2961) );
  OAI21_X1 U1115 ( .B1(n13811), .B2(n13593), .A(n12924), .ZN(n2959) );
  OAI21_X1 U1116 ( .B1(n13811), .B2(n13599), .A(n12924), .ZN(n2957) );
  OAI21_X1 U1117 ( .B1(n13811), .B2(n13605), .A(n12925), .ZN(n2955) );
  OAI21_X1 U1118 ( .B1(n13811), .B2(n13611), .A(n12925), .ZN(n2953) );
  OAI21_X1 U1119 ( .B1(n13811), .B2(n13617), .A(n12925), .ZN(n2951) );
  OAI21_X1 U1120 ( .B1(n13811), .B2(n13623), .A(n12925), .ZN(n2948) );
  OAI21_X1 U1121 ( .B1(n13811), .B2(n13641), .A(n12925), .ZN(n2942) );
  OAI21_X1 U1122 ( .B1(n13811), .B2(n13647), .A(n12925), .ZN(n2940) );
  OAI21_X1 U1123 ( .B1(n13811), .B2(n13653), .A(n12925), .ZN(n2938) );
  OAI21_X1 U1124 ( .B1(n13811), .B2(n13659), .A(n12925), .ZN(n2936) );
  OAI21_X1 U1125 ( .B1(n2866), .B2(n13665), .A(n12925), .ZN(n2934) );
  OAI21_X1 U1126 ( .B1(n13810), .B2(n13671), .A(n12925), .ZN(n2932) );
  OAI21_X1 U1127 ( .B1(n2866), .B2(n13677), .A(n12926), .ZN(n2930) );
  OAI21_X1 U1128 ( .B1(n13810), .B2(n13689), .A(n12926), .ZN(n2926) );
  OAI21_X1 U1129 ( .B1(n13813), .B2(n13695), .A(n12926), .ZN(n2924) );
  OAI21_X1 U1130 ( .B1(n13812), .B2(n13701), .A(n12926), .ZN(n2922) );
  OAI21_X1 U1131 ( .B1(n13811), .B2(n13707), .A(n12926), .ZN(n2920) );
  OAI21_X1 U1132 ( .B1(n2866), .B2(n13713), .A(n12926), .ZN(n2918) );
  OAI21_X1 U1133 ( .B1(n13810), .B2(n13719), .A(n12926), .ZN(n2915) );
  OAI21_X1 U1134 ( .B1(n13813), .B2(n13725), .A(n12926), .ZN(n2912) );
  OAI21_X1 U1135 ( .B1(n13812), .B2(n13731), .A(n12926), .ZN(n2909) );
  NAND2_X1 U1136 ( .A1(n5669), .A2(ADD_RD2[6]), .ZN(n4417) );
  NAND2_X1 U1137 ( .A1(n4276), .A2(ADD_RD1[6]), .ZN(n3133) );
  NAND2_X1 U1138 ( .A1(n4274), .A2(ADD_RD1[6]), .ZN(n3137) );
  NAND2_X1 U1139 ( .A1(n5710), .A2(n5674), .ZN(n4391) );
  NAND2_X1 U1140 ( .A1(n5710), .A2(n5668), .ZN(n4389) );
  NAND2_X1 U1141 ( .A1(n5710), .A2(n5676), .ZN(n4390) );
  NAND2_X1 U1142 ( .A1(n5710), .A2(n5660), .ZN(n4396) );
  NAND2_X1 U1143 ( .A1(n5710), .A2(n5669), .ZN(n4433) );
  NAND2_X1 U1144 ( .A1(n4299), .A2(n4278), .ZN(n3107) );
  NAND2_X1 U1145 ( .A1(n4299), .A2(n4275), .ZN(n3105) );
  NAND2_X1 U1146 ( .A1(n4299), .A2(n4279), .ZN(n3106) );
  NAND2_X1 U1147 ( .A1(n4299), .A2(n4271), .ZN(n3112) );
  NAND2_X1 U1148 ( .A1(n4299), .A2(n4276), .ZN(n3148) );
  BUF_X1 U1149 ( .A(n4325), .Z(n13147) );
  BUF_X1 U1150 ( .A(n4325), .Z(n13148) );
  BUF_X1 U1151 ( .A(n3041), .Z(n13375) );
  BUF_X1 U1152 ( .A(n3041), .Z(n13376) );
  NAND2_X1 U1153 ( .A1(n5690), .A2(n5671), .ZN(n4365) );
  NAND2_X1 U1154 ( .A1(n5690), .A2(n5676), .ZN(n4363) );
  NAND2_X1 U1155 ( .A1(n5690), .A2(n5666), .ZN(n4364) );
  NAND2_X1 U1156 ( .A1(n5691), .A2(n5666), .ZN(n4376) );
  NAND2_X1 U1157 ( .A1(n5691), .A2(n5671), .ZN(n4374) );
  NAND2_X1 U1158 ( .A1(n5691), .A2(n5660), .ZN(n4375) );
  NAND2_X1 U1159 ( .A1(n5691), .A2(n5674), .ZN(n4369) );
  NAND2_X1 U1160 ( .A1(n5691), .A2(n5676), .ZN(n4370) );
  NAND2_X1 U1161 ( .A1(n5690), .A2(n5668), .ZN(n4406) );
  NAND2_X1 U1162 ( .A1(n5690), .A2(n5674), .ZN(n4407) );
  NAND2_X1 U1163 ( .A1(n4289), .A2(n4280), .ZN(n3081) );
  NAND2_X1 U1164 ( .A1(n4289), .A2(n4279), .ZN(n3079) );
  NAND2_X1 U1165 ( .A1(n4289), .A2(n4274), .ZN(n3080) );
  NAND2_X1 U1166 ( .A1(n4290), .A2(n4274), .ZN(n3092) );
  NAND2_X1 U1167 ( .A1(n4290), .A2(n4280), .ZN(n3090) );
  NAND2_X1 U1168 ( .A1(n4290), .A2(n4271), .ZN(n3091) );
  NAND2_X1 U1169 ( .A1(n4290), .A2(n4279), .ZN(n3085) );
  NAND2_X1 U1170 ( .A1(n4290), .A2(n4278), .ZN(n3086) );
  NAND2_X1 U1171 ( .A1(n4289), .A2(n4275), .ZN(n3122) );
  NAND2_X1 U1172 ( .A1(n4289), .A2(n4278), .ZN(n3123) );
  BUF_X1 U1173 ( .A(n4325), .Z(n13145) );
  BUF_X1 U1174 ( .A(n4325), .Z(n13144) );
  BUF_X1 U1175 ( .A(n3041), .Z(n13373) );
  BUF_X1 U1176 ( .A(n3041), .Z(n13372) );
  BUF_X1 U1177 ( .A(n4322), .Z(n13153) );
  BUF_X1 U1178 ( .A(n3038), .Z(n13381) );
  BUF_X1 U1179 ( .A(n4322), .Z(n13154) );
  BUF_X1 U1180 ( .A(n3038), .Z(n13382) );
  NAND2_X1 U1181 ( .A1(n5659), .A2(n5660), .ZN(n4339) );
  NAND2_X1 U1182 ( .A1(n5659), .A2(n5666), .ZN(n4337) );
  NAND2_X1 U1183 ( .A1(n5661), .A2(n5660), .ZN(n4348) );
  NAND2_X1 U1184 ( .A1(n5661), .A2(n5671), .ZN(n4343) );
  NAND2_X1 U1185 ( .A1(n5661), .A2(n5666), .ZN(n4344) );
  NAND2_X1 U1186 ( .A1(n5659), .A2(n5676), .ZN(n4380) );
  NAND2_X1 U1187 ( .A1(n5659), .A2(n5671), .ZN(n4381) );
  NAND2_X1 U1188 ( .A1(n5714), .A2(n5676), .ZN(n4402) );
  NAND2_X1 U1189 ( .A1(n5714), .A2(n5674), .ZN(n4400) );
  NAND2_X1 U1190 ( .A1(n5714), .A2(n5671), .ZN(n4401) );
  NAND2_X1 U1191 ( .A1(n4270), .A2(n4271), .ZN(n3055) );
  NAND2_X1 U1192 ( .A1(n4270), .A2(n4274), .ZN(n3053) );
  NAND2_X1 U1193 ( .A1(n4272), .A2(n4271), .ZN(n3064) );
  NAND2_X1 U1194 ( .A1(n4272), .A2(n4279), .ZN(n3059) );
  NAND2_X1 U1195 ( .A1(n4272), .A2(n4278), .ZN(n3060) );
  NAND2_X1 U1196 ( .A1(n4270), .A2(n4279), .ZN(n3096) );
  NAND2_X1 U1197 ( .A1(n4270), .A2(n4280), .ZN(n3097) );
  NAND2_X1 U1198 ( .A1(n4301), .A2(n4279), .ZN(n3118) );
  NAND2_X1 U1199 ( .A1(n4301), .A2(n4278), .ZN(n3116) );
  NAND2_X1 U1200 ( .A1(n4301), .A2(n4280), .ZN(n3117) );
  BUF_X1 U1201 ( .A(n4325), .Z(n13146) );
  BUF_X1 U1202 ( .A(n3041), .Z(n13374) );
  NAND2_X1 U1203 ( .A1(n5732), .A2(n5668), .ZN(n4428) );
  NAND2_X1 U1204 ( .A1(n5732), .A2(n5669), .ZN(n4426) );
  NAND2_X1 U1205 ( .A1(n5732), .A2(n5674), .ZN(n4427) );
  NAND2_X1 U1206 ( .A1(n4310), .A2(n4275), .ZN(n3144) );
  NAND2_X1 U1207 ( .A1(n4310), .A2(n4276), .ZN(n3142) );
  NAND2_X1 U1208 ( .A1(n4310), .A2(n4278), .ZN(n3143) );
  NOR2_X1 U1209 ( .A1(n16071), .A2(n16070), .ZN(n3009) );
  NOR2_X1 U1210 ( .A1(n16072), .A2(ADD_WR[3]), .ZN(n3031) );
  AND2_X1 U1211 ( .A1(n3009), .A2(n3022), .ZN(n2877) );
  AND2_X1 U1212 ( .A1(n3006), .A2(n3022), .ZN(n2874) );
  AND2_X1 U1213 ( .A1(n3003), .A2(n3022), .ZN(n2871) );
  AND2_X1 U1214 ( .A1(n3022), .A2(n3000), .ZN(n2867) );
  AND2_X1 U1215 ( .A1(n3031), .A2(n3000), .ZN(n2880) );
  AND2_X1 U1216 ( .A1(n3031), .A2(n3006), .ZN(n2886) );
  AND2_X1 U1217 ( .A1(n3031), .A2(n3003), .ZN(n2883) );
  NAND2_X1 U1218 ( .A1(n5666), .A2(ADD_RD2[6]), .ZN(n4421) );
  NAND2_X1 U1219 ( .A1(n5671), .A2(ADD_RD2[6]), .ZN(n4422) );
  NAND2_X1 U1220 ( .A1(n4280), .A2(ADD_RD1[6]), .ZN(n3138) );
  NAND2_X1 U1221 ( .A1(n5664), .A2(ADD_RD2[6]), .ZN(n4415) );
  NAND2_X1 U1222 ( .A1(n4273), .A2(ADD_RD1[6]), .ZN(n3131) );
  NAND2_X1 U1223 ( .A1(n5668), .A2(ADD_RD2[6]), .ZN(n4416) );
  NAND2_X1 U1224 ( .A1(n4275), .A2(ADD_RD1[6]), .ZN(n3132) );
  BUF_X1 U1225 ( .A(n4322), .Z(n13155) );
  BUF_X1 U1226 ( .A(n3038), .Z(n13383) );
  AND2_X1 U1227 ( .A1(n3012), .A2(n3000), .ZN(n2904) );
  AND2_X1 U1228 ( .A1(n2999), .A2(n3000), .ZN(n2892) );
  AND2_X1 U1229 ( .A1(n3012), .A2(n3003), .ZN(n2907) );
  AND2_X1 U1230 ( .A1(n3012), .A2(n3009), .ZN(n2913) );
  AND2_X1 U1231 ( .A1(n3012), .A2(n3006), .ZN(n2910) );
  AND2_X1 U1232 ( .A1(n2999), .A2(n3006), .ZN(n2898) );
  AND2_X1 U1233 ( .A1(n2999), .A2(n3003), .ZN(n2895) );
  INV_X1 U1234 ( .A(ADD_WR[5]), .ZN(n16059) );
  INV_X1 U1235 ( .A(ADD_RD2[5]), .ZN(n16057) );
  INV_X1 U1236 ( .A(ADD_RD1[5]), .ZN(n16055) );
  INV_X1 U1237 ( .A(ADD_WR[4]), .ZN(n16060) );
  INV_X1 U1238 ( .A(ADD_RD2[4]), .ZN(n16058) );
  INV_X1 U1239 ( .A(ADD_RD1[4]), .ZN(n16056) );
  INV_X1 U1240 ( .A(ADD_RD2[3]), .ZN(n16062) );
  INV_X1 U1241 ( .A(ADD_RD1[3]), .ZN(n16061) );
  BUF_X1 U1242 ( .A(n13823), .Z(n13822) );
  AND2_X1 U1243 ( .A1(n5679), .A2(n5668), .ZN(n4345) );
  AND2_X1 U1244 ( .A1(n5679), .A2(n5674), .ZN(n4346) );
  AND2_X1 U1245 ( .A1(n5679), .A2(n5671), .ZN(n4351) );
  AND2_X1 U1246 ( .A1(n5679), .A2(n5676), .ZN(n4352) );
  AND2_X1 U1247 ( .A1(n4282), .A2(n4275), .ZN(n3061) );
  AND2_X1 U1248 ( .A1(n4282), .A2(n4278), .ZN(n3062) );
  AND2_X1 U1249 ( .A1(n4282), .A2(n4274), .ZN(n3067) );
  AND2_X1 U1250 ( .A1(n4282), .A2(n4271), .ZN(n3068) );
  AND2_X1 U1251 ( .A1(n5660), .A2(ADD_RD2[6]), .ZN(n4418) );
  AND2_X1 U1252 ( .A1(n5710), .A2(n5671), .ZN(n4386) );
  AND2_X1 U1253 ( .A1(n5710), .A2(n5666), .ZN(n4387) );
  AND2_X1 U1254 ( .A1(n4299), .A2(n4280), .ZN(n3102) );
  AND2_X1 U1255 ( .A1(n4299), .A2(n4274), .ZN(n3103) );
  AND2_X1 U1256 ( .A1(n5690), .A2(n5660), .ZN(n4360) );
  AND2_X1 U1257 ( .A1(n5691), .A2(n5668), .ZN(n4366) );
  AND2_X1 U1258 ( .A1(n5691), .A2(n5669), .ZN(n4367) );
  AND2_X1 U1259 ( .A1(n5690), .A2(n5669), .ZN(n4403) );
  AND2_X1 U1260 ( .A1(n4289), .A2(n4271), .ZN(n3076) );
  AND2_X1 U1261 ( .A1(n4290), .A2(n4276), .ZN(n3082) );
  AND2_X1 U1262 ( .A1(n4290), .A2(n4275), .ZN(n3083) );
  AND2_X1 U1263 ( .A1(n4289), .A2(n4276), .ZN(n3119) );
  AND2_X1 U1264 ( .A1(n5661), .A2(n5669), .ZN(n4334) );
  AND2_X1 U1265 ( .A1(n5661), .A2(n5668), .ZN(n4335) );
  AND2_X1 U1266 ( .A1(n5661), .A2(n5676), .ZN(n4340) );
  AND2_X1 U1267 ( .A1(n5661), .A2(n5674), .ZN(n4341) );
  AND2_X1 U1268 ( .A1(n5659), .A2(n5669), .ZN(n4372) );
  AND2_X1 U1269 ( .A1(n5659), .A2(n5674), .ZN(n4377) );
  AND2_X1 U1270 ( .A1(n5659), .A2(n5668), .ZN(n4378) );
  AND2_X1 U1271 ( .A1(n5714), .A2(n5666), .ZN(n4397) );
  AND2_X1 U1272 ( .A1(n5714), .A2(n5660), .ZN(n4398) );
  AND2_X1 U1273 ( .A1(n5714), .A2(n5669), .ZN(n4392) );
  AND2_X1 U1274 ( .A1(n5714), .A2(n5668), .ZN(n4393) );
  AND2_X1 U1275 ( .A1(n4272), .A2(n4276), .ZN(n3050) );
  AND2_X1 U1276 ( .A1(n4272), .A2(n4275), .ZN(n3051) );
  AND2_X1 U1277 ( .A1(n4272), .A2(n4280), .ZN(n3056) );
  AND2_X1 U1278 ( .A1(n4272), .A2(n4274), .ZN(n3057) );
  AND2_X1 U1279 ( .A1(n4270), .A2(n4276), .ZN(n3088) );
  AND2_X1 U1280 ( .A1(n4270), .A2(n4278), .ZN(n3093) );
  AND2_X1 U1281 ( .A1(n4270), .A2(n4275), .ZN(n3094) );
  AND2_X1 U1282 ( .A1(n4301), .A2(n4274), .ZN(n3113) );
  AND2_X1 U1283 ( .A1(n4301), .A2(n4271), .ZN(n3114) );
  AND2_X1 U1284 ( .A1(n4301), .A2(n4276), .ZN(n3108) );
  AND2_X1 U1285 ( .A1(n4301), .A2(n4275), .ZN(n3109) );
  AND2_X1 U1286 ( .A1(n5732), .A2(n5660), .ZN(n4429) );
  AND2_X1 U1287 ( .A1(n5732), .A2(n5676), .ZN(n4423) );
  AND2_X1 U1288 ( .A1(n5732), .A2(n5671), .ZN(n4424) );
  AND2_X1 U1289 ( .A1(n5732), .A2(n5666), .ZN(n4430) );
  AND2_X1 U1290 ( .A1(n4310), .A2(n4279), .ZN(n3139) );
  AND2_X1 U1291 ( .A1(n4310), .A2(n4280), .ZN(n3140) );
  AND2_X1 U1292 ( .A1(n4310), .A2(n4274), .ZN(n3145) );
  AND2_X1 U1293 ( .A1(n4310), .A2(n4271), .ZN(n3146) );
  AND2_X1 U1294 ( .A1(n4279), .A2(ADD_RD1[6]), .ZN(n3129) );
  AND2_X1 U1295 ( .A1(n4278), .A2(ADD_RD1[6]), .ZN(n3128) );
  AND2_X1 U1296 ( .A1(n5674), .A2(ADD_RD2[6]), .ZN(n4412) );
  AND2_X1 U1297 ( .A1(n5676), .A2(ADD_RD2[6]), .ZN(n4413) );
  AND2_X1 U1298 ( .A1(n4271), .A2(ADD_RD1[6]), .ZN(n3134) );
  BUF_X1 U1299 ( .A(n13823), .Z(n13821) );
  BUF_X1 U1300 ( .A(n13823), .Z(n13820) );
  BUF_X1 U1301 ( .A(n13816), .Z(n13819) );
  BUF_X1 U1302 ( .A(n13814), .Z(n13818) );
  BUF_X1 U1303 ( .A(n13821), .Z(n13817) );
  BUF_X1 U1304 ( .A(n13823), .Z(n13816) );
  BUF_X1 U1305 ( .A(n13823), .Z(n13815) );
  BUF_X1 U1306 ( .A(n13823), .Z(n13814) );
  AND2_X1 U1307 ( .A1(ADD_WR[3]), .A2(n16072), .ZN(n2999) );
  OAI222_X1 U1308 ( .A1(n14175), .A2(n13338), .B1(n14111), .B2(n13335), .C1(
        n14143), .C2(n13332), .ZN(n3235) );
  OAI222_X1 U1309 ( .A1(n14560), .A2(n13284), .B1(n14496), .B2(n13281), .C1(
        n14528), .C2(n13278), .ZN(n3243) );
  OAI222_X1 U1310 ( .A1(n14174), .A2(n13338), .B1(n14110), .B2(n13335), .C1(
        n14142), .C2(n13332), .ZN(n3198) );
  OAI222_X1 U1311 ( .A1(n14559), .A2(n13284), .B1(n14495), .B2(n13281), .C1(
        n14527), .C2(n13278), .ZN(n3206) );
  OAI222_X1 U1312 ( .A1(n14173), .A2(n13338), .B1(n14109), .B2(n13335), .C1(
        n14141), .C2(n13332), .ZN(n3161) );
  OAI222_X1 U1313 ( .A1(n14558), .A2(n13284), .B1(n14494), .B2(n13281), .C1(
        n14526), .C2(n13278), .ZN(n3169) );
  OAI222_X1 U1314 ( .A1(n14172), .A2(n13338), .B1(n14108), .B2(n13335), .C1(
        n14140), .C2(n13332), .ZN(n3063) );
  OAI222_X1 U1315 ( .A1(n14557), .A2(n13284), .B1(n14493), .B2(n13281), .C1(
        n14525), .C2(n13278), .ZN(n3089) );
  OAI222_X1 U1316 ( .A1(n14178), .A2(n13110), .B1(n14114), .B2(n13107), .C1(
        n14146), .C2(n13104), .ZN(n4630) );
  OAI222_X1 U1317 ( .A1(n14563), .A2(n13056), .B1(n14499), .B2(n13053), .C1(
        n14531), .C2(n13050), .ZN(n4638) );
  OAI222_X1 U1318 ( .A1(n14177), .A2(n13110), .B1(n14113), .B2(n13107), .C1(
        n14145), .C2(n13104), .ZN(n4593) );
  OAI222_X1 U1319 ( .A1(n14562), .A2(n13056), .B1(n14498), .B2(n13053), .C1(
        n14530), .C2(n13050), .ZN(n4601) );
  OAI222_X1 U1320 ( .A1(n14176), .A2(n13110), .B1(n14112), .B2(n13107), .C1(
        n14144), .C2(n13104), .ZN(n4556) );
  OAI222_X1 U1321 ( .A1(n14561), .A2(n13056), .B1(n14497), .B2(n13053), .C1(
        n14529), .C2(n13050), .ZN(n4564) );
  OAI222_X1 U1322 ( .A1(n14175), .A2(n13110), .B1(n14111), .B2(n13107), .C1(
        n14143), .C2(n13104), .ZN(n4519) );
  OAI222_X1 U1323 ( .A1(n14560), .A2(n13056), .B1(n14496), .B2(n13053), .C1(
        n14528), .C2(n13050), .ZN(n4527) );
  OAI222_X1 U1324 ( .A1(n14174), .A2(n13110), .B1(n14110), .B2(n13107), .C1(
        n14142), .C2(n13104), .ZN(n4482) );
  OAI222_X1 U1325 ( .A1(n14559), .A2(n13056), .B1(n14495), .B2(n13053), .C1(
        n14527), .C2(n13050), .ZN(n4490) );
  OAI222_X1 U1326 ( .A1(n14173), .A2(n13110), .B1(n14109), .B2(n13107), .C1(
        n14141), .C2(n13104), .ZN(n4445) );
  OAI222_X1 U1327 ( .A1(n14558), .A2(n13056), .B1(n14494), .B2(n13053), .C1(
        n14526), .C2(n13050), .ZN(n4453) );
  OAI222_X1 U1328 ( .A1(n14172), .A2(n13110), .B1(n14108), .B2(n13107), .C1(
        n14140), .C2(n13104), .ZN(n4347) );
  OAI222_X1 U1329 ( .A1(n14557), .A2(n13056), .B1(n14493), .B2(n13053), .C1(
        n14525), .C2(n13050), .ZN(n4373) );
  OAI222_X1 U1330 ( .A1(n14179), .A2(n13110), .B1(n14115), .B2(n13107), .C1(
        n14147), .C2(n13104), .ZN(n4667) );
  OAI222_X1 U1331 ( .A1(n14564), .A2(n13056), .B1(n14500), .B2(n13053), .C1(
        n14532), .C2(n13050), .ZN(n4675) );
  OAI222_X1 U1332 ( .A1(n14179), .A2(n13338), .B1(n14115), .B2(n13335), .C1(
        n14147), .C2(n13332), .ZN(n3383) );
  OAI222_X1 U1333 ( .A1(n14564), .A2(n13284), .B1(n14500), .B2(n13281), .C1(
        n14532), .C2(n13278), .ZN(n3391) );
  OAI222_X1 U1334 ( .A1(n14178), .A2(n13338), .B1(n14114), .B2(n13335), .C1(
        n14146), .C2(n13332), .ZN(n3346) );
  OAI222_X1 U1335 ( .A1(n14563), .A2(n13284), .B1(n14499), .B2(n13281), .C1(
        n14531), .C2(n13278), .ZN(n3354) );
  OAI222_X1 U1336 ( .A1(n14177), .A2(n13338), .B1(n14113), .B2(n13335), .C1(
        n14145), .C2(n13332), .ZN(n3309) );
  OAI222_X1 U1337 ( .A1(n14562), .A2(n13284), .B1(n14498), .B2(n13281), .C1(
        n14530), .C2(n13278), .ZN(n3317) );
  OAI222_X1 U1338 ( .A1(n14176), .A2(n13338), .B1(n14112), .B2(n13335), .C1(
        n14144), .C2(n13332), .ZN(n3272) );
  OAI222_X1 U1339 ( .A1(n14561), .A2(n13284), .B1(n14497), .B2(n13281), .C1(
        n14529), .C2(n13278), .ZN(n3280) );
  OAI222_X1 U1340 ( .A1(n14203), .A2(n13108), .B1(n14139), .B2(n13105), .C1(
        n14171), .C2(n13102), .ZN(n5678) );
  OAI222_X1 U1341 ( .A1(n14588), .A2(n13054), .B1(n14524), .B2(n13051), .C1(
        n14556), .C2(n13048), .ZN(n5696) );
  OAI222_X1 U1342 ( .A1(n14202), .A2(n13108), .B1(n14138), .B2(n13105), .C1(
        n14170), .C2(n13102), .ZN(n5599) );
  OAI222_X1 U1343 ( .A1(n14587), .A2(n13054), .B1(n14523), .B2(n13051), .C1(
        n14555), .C2(n13048), .ZN(n5611) );
  OAI222_X1 U1344 ( .A1(n14201), .A2(n13108), .B1(n14137), .B2(n13105), .C1(
        n14169), .C2(n13102), .ZN(n5538) );
  OAI222_X1 U1345 ( .A1(n14586), .A2(n13054), .B1(n14522), .B2(n13051), .C1(
        n14554), .C2(n13048), .ZN(n5550) );
  OAI222_X1 U1346 ( .A1(n14200), .A2(n13108), .B1(n14136), .B2(n13105), .C1(
        n14168), .C2(n13102), .ZN(n5476) );
  OAI222_X1 U1347 ( .A1(n14585), .A2(n13054), .B1(n14521), .B2(n13051), .C1(
        n14553), .C2(n13048), .ZN(n5489) );
  OAI222_X1 U1348 ( .A1(n14199), .A2(n13108), .B1(n14135), .B2(n13105), .C1(
        n14167), .C2(n13102), .ZN(n5419) );
  OAI222_X1 U1349 ( .A1(n14584), .A2(n13054), .B1(n14520), .B2(n13051), .C1(
        n14552), .C2(n13048), .ZN(n5430) );
  OAI222_X1 U1350 ( .A1(n14198), .A2(n13108), .B1(n14134), .B2(n13105), .C1(
        n14166), .C2(n13102), .ZN(n5370) );
  OAI222_X1 U1351 ( .A1(n14583), .A2(n13054), .B1(n14519), .B2(n13051), .C1(
        n14551), .C2(n13048), .ZN(n5378) );
  OAI222_X1 U1352 ( .A1(n14197), .A2(n13108), .B1(n14133), .B2(n13105), .C1(
        n14165), .C2(n13102), .ZN(n5333) );
  OAI222_X1 U1353 ( .A1(n14582), .A2(n13054), .B1(n14518), .B2(n13051), .C1(
        n14550), .C2(n13048), .ZN(n5341) );
  OAI222_X1 U1354 ( .A1(n14196), .A2(n13108), .B1(n14132), .B2(n13105), .C1(
        n14164), .C2(n13102), .ZN(n5296) );
  OAI222_X1 U1355 ( .A1(n14581), .A2(n13054), .B1(n14517), .B2(n13051), .C1(
        n14549), .C2(n13048), .ZN(n5304) );
  OAI222_X1 U1356 ( .A1(n14195), .A2(n13108), .B1(n14131), .B2(n13105), .C1(
        n14163), .C2(n13102), .ZN(n5259) );
  OAI222_X1 U1357 ( .A1(n14580), .A2(n13054), .B1(n14516), .B2(n13051), .C1(
        n14548), .C2(n13048), .ZN(n5267) );
  OAI222_X1 U1358 ( .A1(n14194), .A2(n13108), .B1(n14130), .B2(n13105), .C1(
        n14162), .C2(n13102), .ZN(n5222) );
  OAI222_X1 U1359 ( .A1(n14579), .A2(n13054), .B1(n14515), .B2(n13051), .C1(
        n14547), .C2(n13048), .ZN(n5230) );
  OAI222_X1 U1360 ( .A1(n14193), .A2(n13108), .B1(n14129), .B2(n13105), .C1(
        n14161), .C2(n13102), .ZN(n5185) );
  OAI222_X1 U1361 ( .A1(n14578), .A2(n13054), .B1(n14514), .B2(n13051), .C1(
        n14546), .C2(n13048), .ZN(n5193) );
  OAI222_X1 U1362 ( .A1(n14192), .A2(n13108), .B1(n14128), .B2(n13105), .C1(
        n14160), .C2(n13102), .ZN(n5148) );
  OAI222_X1 U1363 ( .A1(n14577), .A2(n13054), .B1(n14513), .B2(n13051), .C1(
        n14545), .C2(n13048), .ZN(n5156) );
  OAI222_X1 U1364 ( .A1(n14191), .A2(n13109), .B1(n14127), .B2(n13106), .C1(
        n14159), .C2(n13103), .ZN(n5111) );
  OAI222_X1 U1365 ( .A1(n14576), .A2(n13055), .B1(n14512), .B2(n13052), .C1(
        n14544), .C2(n13049), .ZN(n5119) );
  OAI222_X1 U1366 ( .A1(n14190), .A2(n13109), .B1(n14126), .B2(n13106), .C1(
        n14158), .C2(n13103), .ZN(n5074) );
  OAI222_X1 U1367 ( .A1(n14575), .A2(n13055), .B1(n14511), .B2(n13052), .C1(
        n14543), .C2(n13049), .ZN(n5082) );
  OAI222_X1 U1368 ( .A1(n14189), .A2(n13109), .B1(n14125), .B2(n13106), .C1(
        n14157), .C2(n13103), .ZN(n5037) );
  OAI222_X1 U1369 ( .A1(n14574), .A2(n13055), .B1(n14510), .B2(n13052), .C1(
        n14542), .C2(n13049), .ZN(n5045) );
  OAI222_X1 U1370 ( .A1(n14188), .A2(n13109), .B1(n14124), .B2(n13106), .C1(
        n14156), .C2(n13103), .ZN(n5000) );
  OAI222_X1 U1371 ( .A1(n14573), .A2(n13055), .B1(n14509), .B2(n13052), .C1(
        n14541), .C2(n13049), .ZN(n5008) );
  OAI222_X1 U1372 ( .A1(n14187), .A2(n13109), .B1(n14123), .B2(n13106), .C1(
        n14155), .C2(n13103), .ZN(n4963) );
  OAI222_X1 U1373 ( .A1(n14572), .A2(n13055), .B1(n14508), .B2(n13052), .C1(
        n14540), .C2(n13049), .ZN(n4971) );
  OAI222_X1 U1374 ( .A1(n14186), .A2(n13109), .B1(n14122), .B2(n13106), .C1(
        n14154), .C2(n13103), .ZN(n4926) );
  OAI222_X1 U1375 ( .A1(n14571), .A2(n13055), .B1(n14507), .B2(n13052), .C1(
        n14539), .C2(n13049), .ZN(n4934) );
  OAI222_X1 U1376 ( .A1(n14185), .A2(n13109), .B1(n14121), .B2(n13106), .C1(
        n14153), .C2(n13103), .ZN(n4889) );
  OAI222_X1 U1377 ( .A1(n14570), .A2(n13055), .B1(n14506), .B2(n13052), .C1(
        n14538), .C2(n13049), .ZN(n4897) );
  OAI222_X1 U1378 ( .A1(n14184), .A2(n13109), .B1(n14120), .B2(n13106), .C1(
        n14152), .C2(n13103), .ZN(n4852) );
  OAI222_X1 U1379 ( .A1(n14569), .A2(n13055), .B1(n14505), .B2(n13052), .C1(
        n14537), .C2(n13049), .ZN(n4860) );
  OAI222_X1 U1380 ( .A1(n14183), .A2(n13109), .B1(n14119), .B2(n13106), .C1(
        n14151), .C2(n13103), .ZN(n4815) );
  OAI222_X1 U1381 ( .A1(n14568), .A2(n13055), .B1(n14504), .B2(n13052), .C1(
        n14536), .C2(n13049), .ZN(n4823) );
  OAI222_X1 U1382 ( .A1(n14182), .A2(n13109), .B1(n14118), .B2(n13106), .C1(
        n14150), .C2(n13103), .ZN(n4778) );
  OAI222_X1 U1383 ( .A1(n14567), .A2(n13055), .B1(n14503), .B2(n13052), .C1(
        n14535), .C2(n13049), .ZN(n4786) );
  OAI222_X1 U1384 ( .A1(n14181), .A2(n13109), .B1(n14117), .B2(n13106), .C1(
        n14149), .C2(n13103), .ZN(n4741) );
  OAI222_X1 U1385 ( .A1(n14566), .A2(n13055), .B1(n14502), .B2(n13052), .C1(
        n14534), .C2(n13049), .ZN(n4749) );
  OAI222_X1 U1386 ( .A1(n14180), .A2(n13109), .B1(n14116), .B2(n13106), .C1(
        n14148), .C2(n13103), .ZN(n4704) );
  OAI222_X1 U1387 ( .A1(n14565), .A2(n13055), .B1(n14501), .B2(n13052), .C1(
        n14533), .C2(n13049), .ZN(n4712) );
  OAI222_X1 U1388 ( .A1(n14203), .A2(n13336), .B1(n14139), .B2(n13333), .C1(
        n14171), .C2(n13330), .ZN(n4281) );
  OAI222_X1 U1389 ( .A1(n14588), .A2(n13282), .B1(n14524), .B2(n13279), .C1(
        n14556), .C2(n13276), .ZN(n4292) );
  OAI222_X1 U1390 ( .A1(n14202), .A2(n13336), .B1(n14138), .B2(n13333), .C1(
        n14170), .C2(n13330), .ZN(n4234) );
  OAI222_X1 U1391 ( .A1(n14587), .A2(n13282), .B1(n14523), .B2(n13279), .C1(
        n14555), .C2(n13276), .ZN(n4242) );
  OAI222_X1 U1392 ( .A1(n14201), .A2(n13336), .B1(n14137), .B2(n13333), .C1(
        n14169), .C2(n13330), .ZN(n4197) );
  OAI222_X1 U1393 ( .A1(n14586), .A2(n13282), .B1(n14522), .B2(n13279), .C1(
        n14554), .C2(n13276), .ZN(n4205) );
  OAI222_X1 U1394 ( .A1(n14200), .A2(n13336), .B1(n14136), .B2(n13333), .C1(
        n14168), .C2(n13330), .ZN(n4160) );
  OAI222_X1 U1395 ( .A1(n14585), .A2(n13282), .B1(n14521), .B2(n13279), .C1(
        n14553), .C2(n13276), .ZN(n4168) );
  OAI222_X1 U1396 ( .A1(n14199), .A2(n13336), .B1(n14135), .B2(n13333), .C1(
        n14167), .C2(n13330), .ZN(n4123) );
  OAI222_X1 U1397 ( .A1(n14584), .A2(n13282), .B1(n14520), .B2(n13279), .C1(
        n14552), .C2(n13276), .ZN(n4131) );
  OAI222_X1 U1398 ( .A1(n14198), .A2(n13336), .B1(n14134), .B2(n13333), .C1(
        n14166), .C2(n13330), .ZN(n4086) );
  OAI222_X1 U1399 ( .A1(n14583), .A2(n13282), .B1(n14519), .B2(n13279), .C1(
        n14551), .C2(n13276), .ZN(n4094) );
  OAI222_X1 U1400 ( .A1(n14197), .A2(n13336), .B1(n14133), .B2(n13333), .C1(
        n14165), .C2(n13330), .ZN(n4049) );
  OAI222_X1 U1401 ( .A1(n14582), .A2(n13282), .B1(n14518), .B2(n13279), .C1(
        n14550), .C2(n13276), .ZN(n4057) );
  OAI222_X1 U1402 ( .A1(n14196), .A2(n13336), .B1(n14132), .B2(n13333), .C1(
        n14164), .C2(n13330), .ZN(n4012) );
  OAI222_X1 U1403 ( .A1(n14581), .A2(n13282), .B1(n14517), .B2(n13279), .C1(
        n14549), .C2(n13276), .ZN(n4020) );
  OAI222_X1 U1404 ( .A1(n14195), .A2(n13336), .B1(n14131), .B2(n13333), .C1(
        n14163), .C2(n13330), .ZN(n3975) );
  OAI222_X1 U1405 ( .A1(n14580), .A2(n13282), .B1(n14516), .B2(n13279), .C1(
        n14548), .C2(n13276), .ZN(n3983) );
  OAI222_X1 U1406 ( .A1(n14194), .A2(n13336), .B1(n14130), .B2(n13333), .C1(
        n14162), .C2(n13330), .ZN(n3938) );
  OAI222_X1 U1407 ( .A1(n14579), .A2(n13282), .B1(n14515), .B2(n13279), .C1(
        n14547), .C2(n13276), .ZN(n3946) );
  OAI222_X1 U1408 ( .A1(n14193), .A2(n13336), .B1(n14129), .B2(n13333), .C1(
        n14161), .C2(n13330), .ZN(n3901) );
  OAI222_X1 U1409 ( .A1(n14578), .A2(n13282), .B1(n14514), .B2(n13279), .C1(
        n14546), .C2(n13276), .ZN(n3909) );
  OAI222_X1 U1410 ( .A1(n14192), .A2(n13336), .B1(n14128), .B2(n13333), .C1(
        n14160), .C2(n13330), .ZN(n3864) );
  OAI222_X1 U1411 ( .A1(n14577), .A2(n13282), .B1(n14513), .B2(n13279), .C1(
        n14545), .C2(n13276), .ZN(n3872) );
  OAI222_X1 U1412 ( .A1(n14191), .A2(n13337), .B1(n14127), .B2(n13334), .C1(
        n14159), .C2(n13331), .ZN(n3827) );
  OAI222_X1 U1413 ( .A1(n14576), .A2(n13283), .B1(n14512), .B2(n13280), .C1(
        n14544), .C2(n13277), .ZN(n3835) );
  OAI222_X1 U1414 ( .A1(n14190), .A2(n13337), .B1(n14126), .B2(n13334), .C1(
        n14158), .C2(n13331), .ZN(n3790) );
  OAI222_X1 U1415 ( .A1(n14575), .A2(n13283), .B1(n14511), .B2(n13280), .C1(
        n14543), .C2(n13277), .ZN(n3798) );
  OAI222_X1 U1416 ( .A1(n14189), .A2(n13337), .B1(n14125), .B2(n13334), .C1(
        n14157), .C2(n13331), .ZN(n3753) );
  OAI222_X1 U1417 ( .A1(n14574), .A2(n13283), .B1(n14510), .B2(n13280), .C1(
        n14542), .C2(n13277), .ZN(n3761) );
  OAI222_X1 U1418 ( .A1(n14188), .A2(n13337), .B1(n14124), .B2(n13334), .C1(
        n14156), .C2(n13331), .ZN(n3716) );
  OAI222_X1 U1419 ( .A1(n14573), .A2(n13283), .B1(n14509), .B2(n13280), .C1(
        n14541), .C2(n13277), .ZN(n3724) );
  OAI222_X1 U1420 ( .A1(n14187), .A2(n13337), .B1(n14123), .B2(n13334), .C1(
        n14155), .C2(n13331), .ZN(n3679) );
  OAI222_X1 U1421 ( .A1(n14572), .A2(n13283), .B1(n14508), .B2(n13280), .C1(
        n14540), .C2(n13277), .ZN(n3687) );
  OAI222_X1 U1422 ( .A1(n14186), .A2(n13337), .B1(n14122), .B2(n13334), .C1(
        n14154), .C2(n13331), .ZN(n3642) );
  OAI222_X1 U1423 ( .A1(n14571), .A2(n13283), .B1(n14507), .B2(n13280), .C1(
        n14539), .C2(n13277), .ZN(n3650) );
  OAI222_X1 U1424 ( .A1(n14185), .A2(n13337), .B1(n14121), .B2(n13334), .C1(
        n14153), .C2(n13331), .ZN(n3605) );
  OAI222_X1 U1425 ( .A1(n14570), .A2(n13283), .B1(n14506), .B2(n13280), .C1(
        n14538), .C2(n13277), .ZN(n3613) );
  OAI222_X1 U1426 ( .A1(n14184), .A2(n13337), .B1(n14120), .B2(n13334), .C1(
        n14152), .C2(n13331), .ZN(n3568) );
  OAI222_X1 U1427 ( .A1(n14569), .A2(n13283), .B1(n14505), .B2(n13280), .C1(
        n14537), .C2(n13277), .ZN(n3576) );
  OAI222_X1 U1428 ( .A1(n14183), .A2(n13337), .B1(n14119), .B2(n13334), .C1(
        n14151), .C2(n13331), .ZN(n3531) );
  OAI222_X1 U1429 ( .A1(n14568), .A2(n13283), .B1(n14504), .B2(n13280), .C1(
        n14536), .C2(n13277), .ZN(n3539) );
  OAI222_X1 U1430 ( .A1(n14182), .A2(n13337), .B1(n14118), .B2(n13334), .C1(
        n14150), .C2(n13331), .ZN(n3494) );
  OAI222_X1 U1431 ( .A1(n14567), .A2(n13283), .B1(n14503), .B2(n13280), .C1(
        n14535), .C2(n13277), .ZN(n3502) );
  OAI222_X1 U1432 ( .A1(n14181), .A2(n13337), .B1(n14117), .B2(n13334), .C1(
        n14149), .C2(n13331), .ZN(n3457) );
  OAI222_X1 U1433 ( .A1(n14566), .A2(n13283), .B1(n14502), .B2(n13280), .C1(
        n14534), .C2(n13277), .ZN(n3465) );
  OAI222_X1 U1434 ( .A1(n14180), .A2(n13337), .B1(n14116), .B2(n13334), .C1(
        n14148), .C2(n13331), .ZN(n3420) );
  OAI222_X1 U1435 ( .A1(n14565), .A2(n13283), .B1(n14501), .B2(n13280), .C1(
        n14533), .C2(n13277), .ZN(n3428) );
  AOI221_X1 U1436 ( .B1(n13141), .B2(n14279), .C1(n13138), .C2(n15897), .A(
        n5658), .ZN(n5656) );
  OAI222_X1 U1437 ( .A1(n14375), .A2(n13135), .B1(n14311), .B2(n13132), .C1(
        n14343), .C2(n13129), .ZN(n5658) );
  AOI221_X1 U1438 ( .B1(n13033), .B2(n15013), .C1(n13030), .C2(n14981), .A(
        n5708), .ZN(n5706) );
  OAI222_X1 U1439 ( .A1(n15109), .A2(n13027), .B1(n15045), .B2(n13024), .C1(
        n15077), .C2(n13021), .ZN(n5708) );
  AOI221_X1 U1440 ( .B1(n13141), .B2(n14278), .C1(n13138), .C2(n15896), .A(
        n5596), .ZN(n5594) );
  OAI222_X1 U1441 ( .A1(n14374), .A2(n13135), .B1(n14310), .B2(n13132), .C1(
        n14342), .C2(n13129), .ZN(n5596) );
  AOI221_X1 U1442 ( .B1(n13033), .B2(n15012), .C1(n13030), .C2(n15612), .A(
        n5621), .ZN(n5620) );
  OAI222_X1 U1443 ( .A1(n15108), .A2(n13027), .B1(n15044), .B2(n13024), .C1(
        n15076), .C2(n13021), .ZN(n5621) );
  AOI221_X1 U1444 ( .B1(n13141), .B2(n14277), .C1(n13138), .C2(n15895), .A(
        n5534), .ZN(n5531) );
  OAI222_X1 U1445 ( .A1(n14373), .A2(n13135), .B1(n14309), .B2(n13132), .C1(
        n14341), .C2(n13129), .ZN(n5534) );
  AOI221_X1 U1446 ( .B1(n13033), .B2(n15011), .C1(n13030), .C2(n15611), .A(
        n5560), .ZN(n5559) );
  OAI222_X1 U1447 ( .A1(n15107), .A2(n13027), .B1(n15043), .B2(n13024), .C1(
        n15075), .C2(n13021), .ZN(n5560) );
  AOI221_X1 U1448 ( .B1(n13141), .B2(n14276), .C1(n13138), .C2(n15894), .A(
        n5471), .ZN(n5470) );
  OAI222_X1 U1449 ( .A1(n14372), .A2(n13135), .B1(n14308), .B2(n13132), .C1(
        n14340), .C2(n13129), .ZN(n5471) );
  AOI221_X1 U1450 ( .B1(n13033), .B2(n15010), .C1(n13030), .C2(n15610), .A(
        n5499), .ZN(n5498) );
  OAI222_X1 U1451 ( .A1(n15106), .A2(n13027), .B1(n15042), .B2(n13024), .C1(
        n15074), .C2(n13021), .ZN(n5499) );
  AOI221_X1 U1452 ( .B1(n13141), .B2(n14275), .C1(n13138), .C2(n15893), .A(
        n5416), .ZN(n5414) );
  OAI222_X1 U1453 ( .A1(n14371), .A2(n13135), .B1(n14307), .B2(n13132), .C1(
        n14339), .C2(n13129), .ZN(n5416) );
  AOI221_X1 U1454 ( .B1(n13033), .B2(n15009), .C1(n13030), .C2(n15609), .A(
        n5439), .ZN(n5438) );
  OAI222_X1 U1455 ( .A1(n15105), .A2(n13027), .B1(n15041), .B2(n13024), .C1(
        n15073), .C2(n13021), .ZN(n5439) );
  AOI221_X1 U1456 ( .B1(n13141), .B2(n14274), .C1(n13138), .C2(n15892), .A(
        n5368), .ZN(n5367) );
  OAI222_X1 U1457 ( .A1(n14370), .A2(n13135), .B1(n14306), .B2(n13132), .C1(
        n14338), .C2(n13129), .ZN(n5368) );
  AOI221_X1 U1458 ( .B1(n13033), .B2(n15008), .C1(n13030), .C2(n15608), .A(
        n5386), .ZN(n5384) );
  OAI222_X1 U1459 ( .A1(n15104), .A2(n13027), .B1(n15040), .B2(n13024), .C1(
        n15072), .C2(n13021), .ZN(n5386) );
  AOI221_X1 U1460 ( .B1(n13141), .B2(n14273), .C1(n13138), .C2(n15891), .A(
        n5331), .ZN(n5330) );
  OAI222_X1 U1461 ( .A1(n14369), .A2(n13135), .B1(n14305), .B2(n13132), .C1(
        n14337), .C2(n13129), .ZN(n5331) );
  AOI221_X1 U1462 ( .B1(n13033), .B2(n15007), .C1(n13030), .C2(n15607), .A(
        n5347), .ZN(n5346) );
  OAI222_X1 U1463 ( .A1(n15103), .A2(n13027), .B1(n15039), .B2(n13024), .C1(
        n15071), .C2(n13021), .ZN(n5347) );
  AOI221_X1 U1464 ( .B1(n13141), .B2(n14272), .C1(n13138), .C2(n15890), .A(
        n5294), .ZN(n5293) );
  OAI222_X1 U1465 ( .A1(n14368), .A2(n13135), .B1(n14304), .B2(n13132), .C1(
        n14336), .C2(n13129), .ZN(n5294) );
  AOI221_X1 U1466 ( .B1(n13033), .B2(n15006), .C1(n13030), .C2(n15606), .A(
        n5310), .ZN(n5309) );
  OAI222_X1 U1467 ( .A1(n15102), .A2(n13027), .B1(n15038), .B2(n13024), .C1(
        n15070), .C2(n13021), .ZN(n5310) );
  AOI221_X1 U1468 ( .B1(n13141), .B2(n14271), .C1(n13138), .C2(n15889), .A(
        n5257), .ZN(n5256) );
  OAI222_X1 U1469 ( .A1(n14367), .A2(n13135), .B1(n14303), .B2(n13132), .C1(
        n14335), .C2(n13129), .ZN(n5257) );
  AOI221_X1 U1470 ( .B1(n13033), .B2(n15005), .C1(n13030), .C2(n15657), .A(
        n5273), .ZN(n5272) );
  OAI222_X1 U1471 ( .A1(n15101), .A2(n13027), .B1(n15037), .B2(n13024), .C1(
        n15069), .C2(n13021), .ZN(n5273) );
  AOI221_X1 U1472 ( .B1(n13141), .B2(n14270), .C1(n13138), .C2(n15888), .A(
        n5220), .ZN(n5219) );
  OAI222_X1 U1473 ( .A1(n14366), .A2(n13135), .B1(n14302), .B2(n13132), .C1(
        n14334), .C2(n13129), .ZN(n5220) );
  AOI221_X1 U1474 ( .B1(n13033), .B2(n15004), .C1(n13030), .C2(n15656), .A(
        n5236), .ZN(n5235) );
  OAI222_X1 U1475 ( .A1(n15100), .A2(n13027), .B1(n15036), .B2(n13024), .C1(
        n15068), .C2(n13021), .ZN(n5236) );
  AOI221_X1 U1476 ( .B1(n13141), .B2(n14269), .C1(n13138), .C2(n15887), .A(
        n5183), .ZN(n5182) );
  OAI222_X1 U1477 ( .A1(n14365), .A2(n13135), .B1(n14301), .B2(n13132), .C1(
        n14333), .C2(n13129), .ZN(n5183) );
  AOI221_X1 U1478 ( .B1(n13033), .B2(n15003), .C1(n13030), .C2(n15655), .A(
        n5199), .ZN(n5198) );
  OAI222_X1 U1479 ( .A1(n15099), .A2(n13027), .B1(n15035), .B2(n13024), .C1(
        n15067), .C2(n13021), .ZN(n5199) );
  AOI221_X1 U1480 ( .B1(n13141), .B2(n14268), .C1(n13138), .C2(n15886), .A(
        n5146), .ZN(n5145) );
  OAI222_X1 U1481 ( .A1(n14364), .A2(n13135), .B1(n14300), .B2(n13132), .C1(
        n14332), .C2(n13129), .ZN(n5146) );
  AOI221_X1 U1482 ( .B1(n13033), .B2(n15002), .C1(n13030), .C2(n15654), .A(
        n5162), .ZN(n5161) );
  OAI222_X1 U1483 ( .A1(n15098), .A2(n13027), .B1(n15034), .B2(n13024), .C1(
        n15066), .C2(n13021), .ZN(n5162) );
  AOI221_X1 U1484 ( .B1(n12980), .B2(n15449), .C1(n12977), .C2(n15417), .A(
        n5133), .ZN(n5132) );
  OAI222_X1 U1485 ( .A1(n15545), .A2(n12974), .B1(n15481), .B2(n12971), .C1(
        n15513), .C2(n12968), .ZN(n5133) );
  AOI221_X1 U1486 ( .B1(n12980), .B2(n15448), .C1(n12977), .C2(n15416), .A(
        n5096), .ZN(n5095) );
  OAI222_X1 U1487 ( .A1(n15544), .A2(n12974), .B1(n15480), .B2(n12971), .C1(
        n15512), .C2(n12968), .ZN(n5096) );
  AOI221_X1 U1488 ( .B1(n12980), .B2(n15447), .C1(n12977), .C2(n15415), .A(
        n5059), .ZN(n5058) );
  OAI222_X1 U1489 ( .A1(n15543), .A2(n12974), .B1(n15479), .B2(n12971), .C1(
        n15511), .C2(n12968), .ZN(n5059) );
  AOI221_X1 U1490 ( .B1(n12980), .B2(n15446), .C1(n12977), .C2(n15414), .A(
        n5022), .ZN(n5021) );
  OAI222_X1 U1491 ( .A1(n15542), .A2(n12974), .B1(n15478), .B2(n12971), .C1(
        n15510), .C2(n12968), .ZN(n5022) );
  AOI221_X1 U1492 ( .B1(n12980), .B2(n15445), .C1(n12977), .C2(n15413), .A(
        n4985), .ZN(n4984) );
  OAI222_X1 U1493 ( .A1(n15541), .A2(n12974), .B1(n15477), .B2(n12971), .C1(
        n15509), .C2(n12968), .ZN(n4985) );
  AOI221_X1 U1494 ( .B1(n12980), .B2(n15444), .C1(n12977), .C2(n15412), .A(
        n4948), .ZN(n4947) );
  OAI222_X1 U1495 ( .A1(n15540), .A2(n12974), .B1(n15476), .B2(n12971), .C1(
        n15508), .C2(n12968), .ZN(n4948) );
  AOI221_X1 U1496 ( .B1(n12980), .B2(n15443), .C1(n12977), .C2(n15411), .A(
        n4911), .ZN(n4910) );
  OAI222_X1 U1497 ( .A1(n15539), .A2(n12974), .B1(n15475), .B2(n12971), .C1(
        n15507), .C2(n12968), .ZN(n4911) );
  AOI221_X1 U1498 ( .B1(n12980), .B2(n15442), .C1(n12977), .C2(n15410), .A(
        n4874), .ZN(n4873) );
  OAI222_X1 U1499 ( .A1(n15538), .A2(n12974), .B1(n15474), .B2(n12971), .C1(
        n15506), .C2(n12968), .ZN(n4874) );
  AOI221_X1 U1500 ( .B1(n13034), .B2(n14993), .C1(n13031), .C2(n15645), .A(
        n4829), .ZN(n4828) );
  OAI222_X1 U1501 ( .A1(n15089), .A2(n13028), .B1(n15025), .B2(n13025), .C1(
        n15057), .C2(n13022), .ZN(n4829) );
  AOI221_X1 U1502 ( .B1(n12980), .B2(n15441), .C1(n12977), .C2(n15409), .A(
        n4837), .ZN(n4836) );
  OAI222_X1 U1503 ( .A1(n15537), .A2(n12974), .B1(n15473), .B2(n12971), .C1(
        n15505), .C2(n12968), .ZN(n4837) );
  AOI221_X1 U1504 ( .B1(n13034), .B2(n14992), .C1(n13031), .C2(n15644), .A(
        n4792), .ZN(n4791) );
  OAI222_X1 U1505 ( .A1(n15088), .A2(n13028), .B1(n15024), .B2(n13025), .C1(
        n15056), .C2(n13022), .ZN(n4792) );
  AOI221_X1 U1506 ( .B1(n12980), .B2(n15440), .C1(n12977), .C2(n15408), .A(
        n4800), .ZN(n4799) );
  OAI222_X1 U1507 ( .A1(n15536), .A2(n12974), .B1(n15472), .B2(n12971), .C1(
        n15504), .C2(n12968), .ZN(n4800) );
  AOI221_X1 U1508 ( .B1(n13034), .B2(n14991), .C1(n13031), .C2(n15643), .A(
        n4755), .ZN(n4754) );
  OAI222_X1 U1509 ( .A1(n15087), .A2(n13028), .B1(n15023), .B2(n13025), .C1(
        n15055), .C2(n13022), .ZN(n4755) );
  AOI221_X1 U1510 ( .B1(n12980), .B2(n15439), .C1(n12977), .C2(n15407), .A(
        n4763), .ZN(n4762) );
  OAI222_X1 U1511 ( .A1(n15535), .A2(n12974), .B1(n15471), .B2(n12971), .C1(
        n15503), .C2(n12968), .ZN(n4763) );
  AOI221_X1 U1512 ( .B1(n13034), .B2(n14990), .C1(n13031), .C2(n15642), .A(
        n4718), .ZN(n4717) );
  OAI222_X1 U1513 ( .A1(n15086), .A2(n13028), .B1(n15022), .B2(n13025), .C1(
        n15054), .C2(n13022), .ZN(n4718) );
  AOI221_X1 U1514 ( .B1(n12980), .B2(n15438), .C1(n12977), .C2(n15406), .A(
        n4726), .ZN(n4725) );
  OAI222_X1 U1515 ( .A1(n15534), .A2(n12974), .B1(n15470), .B2(n12971), .C1(
        n15502), .C2(n12968), .ZN(n4726) );
  AOI221_X1 U1516 ( .B1(n13369), .B2(n14279), .C1(n13366), .C2(n15897), .A(
        n4269), .ZN(n4268) );
  OAI222_X1 U1517 ( .A1(n14375), .A2(n13363), .B1(n14311), .B2(n13360), .C1(
        n14343), .C2(n13357), .ZN(n4269) );
  AOI221_X1 U1518 ( .B1(n13261), .B2(n15013), .C1(n13258), .C2(n14981), .A(
        n4298), .ZN(n4297) );
  OAI222_X1 U1519 ( .A1(n15109), .A2(n13255), .B1(n15045), .B2(n13252), .C1(
        n15077), .C2(n13249), .ZN(n4298) );
  AOI221_X1 U1520 ( .B1(n13369), .B2(n14278), .C1(n13366), .C2(n15896), .A(
        n4232), .ZN(n4231) );
  OAI222_X1 U1521 ( .A1(n14374), .A2(n13363), .B1(n14310), .B2(n13360), .C1(
        n14342), .C2(n13357), .ZN(n4232) );
  AOI221_X1 U1522 ( .B1(n13261), .B2(n15012), .C1(n13258), .C2(n15612), .A(
        n4248), .ZN(n4247) );
  OAI222_X1 U1523 ( .A1(n15108), .A2(n13255), .B1(n15044), .B2(n13252), .C1(
        n15076), .C2(n13249), .ZN(n4248) );
  AOI221_X1 U1524 ( .B1(n13369), .B2(n14277), .C1(n13366), .C2(n15895), .A(
        n4195), .ZN(n4194) );
  OAI222_X1 U1525 ( .A1(n14373), .A2(n13363), .B1(n14309), .B2(n13360), .C1(
        n14341), .C2(n13357), .ZN(n4195) );
  AOI221_X1 U1526 ( .B1(n13261), .B2(n15011), .C1(n13258), .C2(n15611), .A(
        n4211), .ZN(n4210) );
  OAI222_X1 U1527 ( .A1(n15107), .A2(n13255), .B1(n15043), .B2(n13252), .C1(
        n15075), .C2(n13249), .ZN(n4211) );
  AOI221_X1 U1528 ( .B1(n13369), .B2(n14276), .C1(n13366), .C2(n15894), .A(
        n4158), .ZN(n4157) );
  OAI222_X1 U1529 ( .A1(n14372), .A2(n13363), .B1(n14308), .B2(n13360), .C1(
        n14340), .C2(n13357), .ZN(n4158) );
  AOI221_X1 U1530 ( .B1(n13261), .B2(n15010), .C1(n13258), .C2(n15610), .A(
        n4174), .ZN(n4173) );
  OAI222_X1 U1531 ( .A1(n15106), .A2(n13255), .B1(n15042), .B2(n13252), .C1(
        n15074), .C2(n13249), .ZN(n4174) );
  AOI221_X1 U1532 ( .B1(n13369), .B2(n14275), .C1(n13366), .C2(n15893), .A(
        n4121), .ZN(n4120) );
  OAI222_X1 U1533 ( .A1(n14371), .A2(n13363), .B1(n14307), .B2(n13360), .C1(
        n14339), .C2(n13357), .ZN(n4121) );
  AOI221_X1 U1534 ( .B1(n13261), .B2(n15009), .C1(n13258), .C2(n15609), .A(
        n4137), .ZN(n4136) );
  OAI222_X1 U1535 ( .A1(n15105), .A2(n13255), .B1(n15041), .B2(n13252), .C1(
        n15073), .C2(n13249), .ZN(n4137) );
  AOI221_X1 U1536 ( .B1(n13369), .B2(n14274), .C1(n13366), .C2(n15892), .A(
        n4084), .ZN(n4083) );
  OAI222_X1 U1537 ( .A1(n14370), .A2(n13363), .B1(n14306), .B2(n13360), .C1(
        n14338), .C2(n13357), .ZN(n4084) );
  AOI221_X1 U1538 ( .B1(n13261), .B2(n15008), .C1(n13258), .C2(n15608), .A(
        n4100), .ZN(n4099) );
  OAI222_X1 U1539 ( .A1(n15104), .A2(n13255), .B1(n15040), .B2(n13252), .C1(
        n15072), .C2(n13249), .ZN(n4100) );
  AOI221_X1 U1540 ( .B1(n13369), .B2(n14273), .C1(n13366), .C2(n15891), .A(
        n4047), .ZN(n4046) );
  OAI222_X1 U1541 ( .A1(n14369), .A2(n13363), .B1(n14305), .B2(n13360), .C1(
        n14337), .C2(n13357), .ZN(n4047) );
  AOI221_X1 U1542 ( .B1(n13261), .B2(n15007), .C1(n13258), .C2(n15607), .A(
        n4063), .ZN(n4062) );
  OAI222_X1 U1543 ( .A1(n15103), .A2(n13255), .B1(n15039), .B2(n13252), .C1(
        n15071), .C2(n13249), .ZN(n4063) );
  AOI221_X1 U1544 ( .B1(n13369), .B2(n14272), .C1(n13366), .C2(n15890), .A(
        n4010), .ZN(n4009) );
  OAI222_X1 U1545 ( .A1(n14368), .A2(n13363), .B1(n14304), .B2(n13360), .C1(
        n14336), .C2(n13357), .ZN(n4010) );
  AOI221_X1 U1546 ( .B1(n13261), .B2(n15006), .C1(n13258), .C2(n15606), .A(
        n4026), .ZN(n4025) );
  OAI222_X1 U1547 ( .A1(n15102), .A2(n13255), .B1(n15038), .B2(n13252), .C1(
        n15070), .C2(n13249), .ZN(n4026) );
  AOI221_X1 U1548 ( .B1(n13369), .B2(n14271), .C1(n13366), .C2(n15889), .A(
        n3973), .ZN(n3972) );
  OAI222_X1 U1549 ( .A1(n14367), .A2(n13363), .B1(n14303), .B2(n13360), .C1(
        n14335), .C2(n13357), .ZN(n3973) );
  AOI221_X1 U1550 ( .B1(n13261), .B2(n15005), .C1(n13258), .C2(n15657), .A(
        n3989), .ZN(n3988) );
  OAI222_X1 U1551 ( .A1(n15101), .A2(n13255), .B1(n15037), .B2(n13252), .C1(
        n15069), .C2(n13249), .ZN(n3989) );
  AOI221_X1 U1552 ( .B1(n13369), .B2(n14270), .C1(n13366), .C2(n15888), .A(
        n3936), .ZN(n3935) );
  OAI222_X1 U1553 ( .A1(n14366), .A2(n13363), .B1(n14302), .B2(n13360), .C1(
        n14334), .C2(n13357), .ZN(n3936) );
  AOI221_X1 U1554 ( .B1(n13261), .B2(n15004), .C1(n13258), .C2(n15656), .A(
        n3952), .ZN(n3951) );
  OAI222_X1 U1555 ( .A1(n15100), .A2(n13255), .B1(n15036), .B2(n13252), .C1(
        n15068), .C2(n13249), .ZN(n3952) );
  AOI221_X1 U1556 ( .B1(n13369), .B2(n14269), .C1(n13366), .C2(n15887), .A(
        n3899), .ZN(n3898) );
  OAI222_X1 U1557 ( .A1(n14365), .A2(n13363), .B1(n14301), .B2(n13360), .C1(
        n14333), .C2(n13357), .ZN(n3899) );
  AOI221_X1 U1558 ( .B1(n13261), .B2(n15003), .C1(n13258), .C2(n15655), .A(
        n3915), .ZN(n3914) );
  OAI222_X1 U1559 ( .A1(n15099), .A2(n13255), .B1(n15035), .B2(n13252), .C1(
        n15067), .C2(n13249), .ZN(n3915) );
  AOI221_X1 U1560 ( .B1(n13369), .B2(n14268), .C1(n13366), .C2(n15886), .A(
        n3862), .ZN(n3861) );
  OAI222_X1 U1561 ( .A1(n14364), .A2(n13363), .B1(n14300), .B2(n13360), .C1(
        n14332), .C2(n13357), .ZN(n3862) );
  AOI221_X1 U1562 ( .B1(n13261), .B2(n15002), .C1(n13258), .C2(n15654), .A(
        n3878), .ZN(n3877) );
  OAI222_X1 U1563 ( .A1(n15098), .A2(n13255), .B1(n15034), .B2(n13252), .C1(
        n15066), .C2(n13249), .ZN(n3878) );
  AOI221_X1 U1564 ( .B1(n13208), .B2(n15449), .C1(n13205), .C2(n15417), .A(
        n3849), .ZN(n3848) );
  OAI222_X1 U1565 ( .A1(n15545), .A2(n13202), .B1(n15481), .B2(n13199), .C1(
        n15513), .C2(n13196), .ZN(n3849) );
  AOI221_X1 U1566 ( .B1(n13208), .B2(n15448), .C1(n13205), .C2(n15416), .A(
        n3812), .ZN(n3811) );
  OAI222_X1 U1567 ( .A1(n15544), .A2(n13202), .B1(n15480), .B2(n13199), .C1(
        n15512), .C2(n13196), .ZN(n3812) );
  AOI221_X1 U1568 ( .B1(n13208), .B2(n15447), .C1(n13205), .C2(n15415), .A(
        n3775), .ZN(n3774) );
  OAI222_X1 U1569 ( .A1(n15543), .A2(n13202), .B1(n15479), .B2(n13199), .C1(
        n15511), .C2(n13196), .ZN(n3775) );
  AOI221_X1 U1570 ( .B1(n13208), .B2(n15446), .C1(n13205), .C2(n15414), .A(
        n3738), .ZN(n3737) );
  OAI222_X1 U1571 ( .A1(n15542), .A2(n13202), .B1(n15478), .B2(n13199), .C1(
        n15510), .C2(n13196), .ZN(n3738) );
  AOI221_X1 U1572 ( .B1(n13208), .B2(n15445), .C1(n13205), .C2(n15413), .A(
        n3701), .ZN(n3700) );
  OAI222_X1 U1573 ( .A1(n15541), .A2(n13202), .B1(n15477), .B2(n13199), .C1(
        n15509), .C2(n13196), .ZN(n3701) );
  AOI221_X1 U1574 ( .B1(n13208), .B2(n15444), .C1(n13205), .C2(n15412), .A(
        n3664), .ZN(n3663) );
  OAI222_X1 U1575 ( .A1(n15540), .A2(n13202), .B1(n15476), .B2(n13199), .C1(
        n15508), .C2(n13196), .ZN(n3664) );
  AOI221_X1 U1576 ( .B1(n13208), .B2(n15443), .C1(n13205), .C2(n15411), .A(
        n3627), .ZN(n3626) );
  OAI222_X1 U1577 ( .A1(n15539), .A2(n13202), .B1(n15475), .B2(n13199), .C1(
        n15507), .C2(n13196), .ZN(n3627) );
  AOI221_X1 U1578 ( .B1(n13208), .B2(n15442), .C1(n13205), .C2(n15410), .A(
        n3590), .ZN(n3589) );
  OAI222_X1 U1579 ( .A1(n15538), .A2(n13202), .B1(n15474), .B2(n13199), .C1(
        n15506), .C2(n13196), .ZN(n3590) );
  AOI221_X1 U1580 ( .B1(n13262), .B2(n14993), .C1(n13259), .C2(n15645), .A(
        n3545), .ZN(n3544) );
  OAI222_X1 U1581 ( .A1(n15089), .A2(n13256), .B1(n15025), .B2(n13253), .C1(
        n15057), .C2(n13250), .ZN(n3545) );
  AOI221_X1 U1582 ( .B1(n13208), .B2(n15441), .C1(n13205), .C2(n15409), .A(
        n3553), .ZN(n3552) );
  OAI222_X1 U1583 ( .A1(n15537), .A2(n13202), .B1(n15473), .B2(n13199), .C1(
        n15505), .C2(n13196), .ZN(n3553) );
  AOI221_X1 U1584 ( .B1(n13262), .B2(n14992), .C1(n13259), .C2(n15644), .A(
        n3508), .ZN(n3507) );
  OAI222_X1 U1585 ( .A1(n15088), .A2(n13256), .B1(n15024), .B2(n13253), .C1(
        n15056), .C2(n13250), .ZN(n3508) );
  AOI221_X1 U1586 ( .B1(n13208), .B2(n15440), .C1(n13205), .C2(n15408), .A(
        n3516), .ZN(n3515) );
  OAI222_X1 U1587 ( .A1(n15536), .A2(n13202), .B1(n15472), .B2(n13199), .C1(
        n15504), .C2(n13196), .ZN(n3516) );
  AOI221_X1 U1588 ( .B1(n13262), .B2(n14991), .C1(n13259), .C2(n15643), .A(
        n3471), .ZN(n3470) );
  OAI222_X1 U1589 ( .A1(n15087), .A2(n13256), .B1(n15023), .B2(n13253), .C1(
        n15055), .C2(n13250), .ZN(n3471) );
  AOI221_X1 U1590 ( .B1(n13208), .B2(n15439), .C1(n13205), .C2(n15407), .A(
        n3479), .ZN(n3478) );
  OAI222_X1 U1591 ( .A1(n15535), .A2(n13202), .B1(n15471), .B2(n13199), .C1(
        n15503), .C2(n13196), .ZN(n3479) );
  AOI221_X1 U1592 ( .B1(n13262), .B2(n14990), .C1(n13259), .C2(n15642), .A(
        n3434), .ZN(n3433) );
  OAI222_X1 U1593 ( .A1(n15086), .A2(n13256), .B1(n15022), .B2(n13253), .C1(
        n15054), .C2(n13250), .ZN(n3434) );
  AOI221_X1 U1594 ( .B1(n13208), .B2(n15438), .C1(n13205), .C2(n15406), .A(
        n3442), .ZN(n3441) );
  OAI222_X1 U1595 ( .A1(n15534), .A2(n13202), .B1(n15470), .B2(n13199), .C1(
        n15502), .C2(n13196), .ZN(n3442) );
  AOI221_X1 U1596 ( .B1(n13371), .B2(n14251), .C1(n13368), .C2(n15593), .A(
        n3233), .ZN(n3232) );
  OAI222_X1 U1597 ( .A1(n14347), .A2(n13365), .B1(n14283), .B2(n13362), .C1(
        n14315), .C2(n13359), .ZN(n3233) );
  AOI221_X1 U1598 ( .B1(n13317), .B2(n14663), .C1(n13314), .C2(n15569), .A(
        n3241), .ZN(n3240) );
  OAI222_X1 U1599 ( .A1(n14759), .A2(n13311), .B1(n14695), .B2(n13308), .C1(
        n14727), .C2(n13305), .ZN(n3241) );
  AOI221_X1 U1600 ( .B1(n13263), .B2(n14985), .C1(n13260), .C2(n15637), .A(
        n3249), .ZN(n3248) );
  OAI222_X1 U1601 ( .A1(n15081), .A2(n13257), .B1(n15017), .B2(n13254), .C1(
        n15049), .C2(n13251), .ZN(n3249) );
  AOI221_X1 U1602 ( .B1(n13209), .B2(n15433), .C1(n13206), .C2(n15401), .A(
        n3257), .ZN(n3256) );
  OAI222_X1 U1603 ( .A1(n15529), .A2(n13203), .B1(n15465), .B2(n13200), .C1(
        n15497), .C2(n13197), .ZN(n3257) );
  AOI221_X1 U1604 ( .B1(n13371), .B2(n14250), .C1(n13368), .C2(n15592), .A(
        n3196), .ZN(n3195) );
  OAI222_X1 U1605 ( .A1(n14346), .A2(n13365), .B1(n14282), .B2(n13362), .C1(
        n14314), .C2(n13359), .ZN(n3196) );
  AOI221_X1 U1606 ( .B1(n13317), .B2(n14662), .C1(n13314), .C2(n15568), .A(
        n3204), .ZN(n3203) );
  OAI222_X1 U1607 ( .A1(n14758), .A2(n13311), .B1(n14694), .B2(n13308), .C1(
        n14726), .C2(n13305), .ZN(n3204) );
  AOI221_X1 U1608 ( .B1(n13263), .B2(n14984), .C1(n13260), .C2(n15636), .A(
        n3212), .ZN(n3211) );
  OAI222_X1 U1609 ( .A1(n15080), .A2(n13257), .B1(n15016), .B2(n13254), .C1(
        n15048), .C2(n13251), .ZN(n3212) );
  AOI221_X1 U1610 ( .B1(n13209), .B2(n15432), .C1(n13206), .C2(n15400), .A(
        n3220), .ZN(n3219) );
  OAI222_X1 U1611 ( .A1(n15528), .A2(n13203), .B1(n15464), .B2(n13200), .C1(
        n15496), .C2(n13197), .ZN(n3220) );
  AOI221_X1 U1612 ( .B1(n13371), .B2(n14249), .C1(n13368), .C2(n15591), .A(
        n3159), .ZN(n3158) );
  OAI222_X1 U1613 ( .A1(n14345), .A2(n13365), .B1(n14281), .B2(n13362), .C1(
        n14313), .C2(n13359), .ZN(n3159) );
  AOI221_X1 U1614 ( .B1(n13317), .B2(n14661), .C1(n13314), .C2(n15567), .A(
        n3167), .ZN(n3166) );
  OAI222_X1 U1615 ( .A1(n14757), .A2(n13311), .B1(n14693), .B2(n13308), .C1(
        n14725), .C2(n13305), .ZN(n3167) );
  AOI221_X1 U1616 ( .B1(n13263), .B2(n14983), .C1(n13260), .C2(n15635), .A(
        n3175), .ZN(n3174) );
  OAI222_X1 U1617 ( .A1(n15079), .A2(n13257), .B1(n15015), .B2(n13254), .C1(
        n15047), .C2(n13251), .ZN(n3175) );
  AOI221_X1 U1618 ( .B1(n13209), .B2(n15431), .C1(n13206), .C2(n15399), .A(
        n3183), .ZN(n3182) );
  OAI222_X1 U1619 ( .A1(n15527), .A2(n13203), .B1(n15463), .B2(n13200), .C1(
        n15495), .C2(n13197), .ZN(n3183) );
  AOI221_X1 U1620 ( .B1(n13371), .B2(n14248), .C1(n13368), .C2(n15590), .A(
        n3052), .ZN(n3049) );
  OAI222_X1 U1621 ( .A1(n14344), .A2(n13365), .B1(n14280), .B2(n13362), .C1(
        n14312), .C2(n13359), .ZN(n3052) );
  AOI221_X1 U1622 ( .B1(n13317), .B2(n14660), .C1(n13314), .C2(n15566), .A(
        n3078), .ZN(n3075) );
  OAI222_X1 U1623 ( .A1(n14756), .A2(n13311), .B1(n14692), .B2(n13308), .C1(
        n14724), .C2(n13305), .ZN(n3078) );
  AOI221_X1 U1624 ( .B1(n13263), .B2(n14982), .C1(n13260), .C2(n15634), .A(
        n3104), .ZN(n3101) );
  OAI222_X1 U1625 ( .A1(n15078), .A2(n13257), .B1(n15014), .B2(n13254), .C1(
        n15046), .C2(n13251), .ZN(n3104) );
  AOI221_X1 U1626 ( .B1(n13209), .B2(n15430), .C1(n13206), .C2(n15398), .A(
        n3130), .ZN(n3127) );
  OAI222_X1 U1627 ( .A1(n15526), .A2(n13203), .B1(n15462), .B2(n13200), .C1(
        n15494), .C2(n13197), .ZN(n3130) );
  AOI221_X1 U1628 ( .B1(n13143), .B2(n14254), .C1(n13140), .C2(n15596), .A(
        n4628), .ZN(n4627) );
  OAI222_X1 U1629 ( .A1(n14350), .A2(n13137), .B1(n14286), .B2(n13134), .C1(
        n14318), .C2(n13131), .ZN(n4628) );
  AOI221_X1 U1630 ( .B1(n13089), .B2(n14666), .C1(n13086), .C2(n15572), .A(
        n4636), .ZN(n4635) );
  OAI222_X1 U1631 ( .A1(n14762), .A2(n13083), .B1(n14698), .B2(n13080), .C1(
        n14730), .C2(n13077), .ZN(n4636) );
  AOI221_X1 U1632 ( .B1(n13035), .B2(n14988), .C1(n13032), .C2(n15640), .A(
        n4644), .ZN(n4643) );
  OAI222_X1 U1633 ( .A1(n15084), .A2(n13029), .B1(n15020), .B2(n13026), .C1(
        n15052), .C2(n13023), .ZN(n4644) );
  AOI221_X1 U1634 ( .B1(n12981), .B2(n15436), .C1(n12978), .C2(n15404), .A(
        n4652), .ZN(n4651) );
  OAI222_X1 U1635 ( .A1(n15532), .A2(n12975), .B1(n15468), .B2(n12972), .C1(
        n15500), .C2(n12969), .ZN(n4652) );
  AOI221_X1 U1636 ( .B1(n13143), .B2(n14253), .C1(n13140), .C2(n15595), .A(
        n4591), .ZN(n4590) );
  OAI222_X1 U1637 ( .A1(n14349), .A2(n13137), .B1(n14285), .B2(n13134), .C1(
        n14317), .C2(n13131), .ZN(n4591) );
  AOI221_X1 U1638 ( .B1(n13089), .B2(n14665), .C1(n13086), .C2(n15571), .A(
        n4599), .ZN(n4598) );
  OAI222_X1 U1639 ( .A1(n14761), .A2(n13083), .B1(n14697), .B2(n13080), .C1(
        n14729), .C2(n13077), .ZN(n4599) );
  AOI221_X1 U1640 ( .B1(n13035), .B2(n14987), .C1(n13032), .C2(n15639), .A(
        n4607), .ZN(n4606) );
  OAI222_X1 U1641 ( .A1(n15083), .A2(n13029), .B1(n15019), .B2(n13026), .C1(
        n15051), .C2(n13023), .ZN(n4607) );
  AOI221_X1 U1642 ( .B1(n12981), .B2(n15435), .C1(n12978), .C2(n15403), .A(
        n4615), .ZN(n4614) );
  OAI222_X1 U1643 ( .A1(n15531), .A2(n12975), .B1(n15467), .B2(n12972), .C1(
        n15499), .C2(n12969), .ZN(n4615) );
  AOI221_X1 U1644 ( .B1(n13143), .B2(n14252), .C1(n13140), .C2(n15594), .A(
        n4554), .ZN(n4553) );
  OAI222_X1 U1645 ( .A1(n14348), .A2(n13137), .B1(n14284), .B2(n13134), .C1(
        n14316), .C2(n13131), .ZN(n4554) );
  AOI221_X1 U1646 ( .B1(n13089), .B2(n14664), .C1(n13086), .C2(n15570), .A(
        n4562), .ZN(n4561) );
  OAI222_X1 U1647 ( .A1(n14760), .A2(n13083), .B1(n14696), .B2(n13080), .C1(
        n14728), .C2(n13077), .ZN(n4562) );
  AOI221_X1 U1648 ( .B1(n13035), .B2(n14986), .C1(n13032), .C2(n15638), .A(
        n4570), .ZN(n4569) );
  OAI222_X1 U1649 ( .A1(n15082), .A2(n13029), .B1(n15018), .B2(n13026), .C1(
        n15050), .C2(n13023), .ZN(n4570) );
  AOI221_X1 U1650 ( .B1(n12981), .B2(n15434), .C1(n12978), .C2(n15402), .A(
        n4578), .ZN(n4577) );
  OAI222_X1 U1651 ( .A1(n15530), .A2(n12975), .B1(n15466), .B2(n12972), .C1(
        n15498), .C2(n12969), .ZN(n4578) );
  AOI221_X1 U1652 ( .B1(n13143), .B2(n14251), .C1(n13140), .C2(n15593), .A(
        n4517), .ZN(n4516) );
  OAI222_X1 U1653 ( .A1(n14347), .A2(n13137), .B1(n14283), .B2(n13134), .C1(
        n14315), .C2(n13131), .ZN(n4517) );
  AOI221_X1 U1654 ( .B1(n13089), .B2(n14663), .C1(n13086), .C2(n15569), .A(
        n4525), .ZN(n4524) );
  OAI222_X1 U1655 ( .A1(n14759), .A2(n13083), .B1(n14695), .B2(n13080), .C1(
        n14727), .C2(n13077), .ZN(n4525) );
  AOI221_X1 U1656 ( .B1(n13035), .B2(n14985), .C1(n13032), .C2(n15637), .A(
        n4533), .ZN(n4532) );
  OAI222_X1 U1657 ( .A1(n15081), .A2(n13029), .B1(n15017), .B2(n13026), .C1(
        n15049), .C2(n13023), .ZN(n4533) );
  AOI221_X1 U1658 ( .B1(n12981), .B2(n15433), .C1(n12978), .C2(n15401), .A(
        n4541), .ZN(n4540) );
  OAI222_X1 U1659 ( .A1(n15529), .A2(n12975), .B1(n15465), .B2(n12972), .C1(
        n15497), .C2(n12969), .ZN(n4541) );
  AOI221_X1 U1660 ( .B1(n13143), .B2(n14250), .C1(n13140), .C2(n15592), .A(
        n4480), .ZN(n4479) );
  OAI222_X1 U1661 ( .A1(n14346), .A2(n13137), .B1(n14282), .B2(n13134), .C1(
        n14314), .C2(n13131), .ZN(n4480) );
  AOI221_X1 U1662 ( .B1(n13089), .B2(n14662), .C1(n13086), .C2(n15568), .A(
        n4488), .ZN(n4487) );
  OAI222_X1 U1663 ( .A1(n14758), .A2(n13083), .B1(n14694), .B2(n13080), .C1(
        n14726), .C2(n13077), .ZN(n4488) );
  AOI221_X1 U1664 ( .B1(n13035), .B2(n14984), .C1(n13032), .C2(n15636), .A(
        n4496), .ZN(n4495) );
  OAI222_X1 U1665 ( .A1(n15080), .A2(n13029), .B1(n15016), .B2(n13026), .C1(
        n15048), .C2(n13023), .ZN(n4496) );
  AOI221_X1 U1666 ( .B1(n12981), .B2(n15432), .C1(n12978), .C2(n15400), .A(
        n4504), .ZN(n4503) );
  OAI222_X1 U1667 ( .A1(n15528), .A2(n12975), .B1(n15464), .B2(n12972), .C1(
        n15496), .C2(n12969), .ZN(n4504) );
  AOI221_X1 U1668 ( .B1(n13143), .B2(n14249), .C1(n13140), .C2(n15591), .A(
        n4443), .ZN(n4442) );
  OAI222_X1 U1669 ( .A1(n14345), .A2(n13137), .B1(n14281), .B2(n13134), .C1(
        n14313), .C2(n13131), .ZN(n4443) );
  AOI221_X1 U1670 ( .B1(n13089), .B2(n14661), .C1(n13086), .C2(n15567), .A(
        n4451), .ZN(n4450) );
  OAI222_X1 U1671 ( .A1(n14757), .A2(n13083), .B1(n14693), .B2(n13080), .C1(
        n14725), .C2(n13077), .ZN(n4451) );
  AOI221_X1 U1672 ( .B1(n13035), .B2(n14983), .C1(n13032), .C2(n15635), .A(
        n4459), .ZN(n4458) );
  OAI222_X1 U1673 ( .A1(n15079), .A2(n13029), .B1(n15015), .B2(n13026), .C1(
        n15047), .C2(n13023), .ZN(n4459) );
  AOI221_X1 U1674 ( .B1(n12981), .B2(n15431), .C1(n12978), .C2(n15399), .A(
        n4467), .ZN(n4466) );
  OAI222_X1 U1675 ( .A1(n15527), .A2(n12975), .B1(n15463), .B2(n12972), .C1(
        n15495), .C2(n12969), .ZN(n4467) );
  AOI221_X1 U1676 ( .B1(n13143), .B2(n14248), .C1(n13140), .C2(n15590), .A(
        n4336), .ZN(n4333) );
  OAI222_X1 U1677 ( .A1(n14344), .A2(n13137), .B1(n14280), .B2(n13134), .C1(
        n14312), .C2(n13131), .ZN(n4336) );
  AOI221_X1 U1678 ( .B1(n13089), .B2(n14660), .C1(n13086), .C2(n15566), .A(
        n4362), .ZN(n4359) );
  OAI222_X1 U1679 ( .A1(n14756), .A2(n13083), .B1(n14692), .B2(n13080), .C1(
        n14724), .C2(n13077), .ZN(n4362) );
  AOI221_X1 U1680 ( .B1(n13035), .B2(n14982), .C1(n13032), .C2(n15634), .A(
        n4388), .ZN(n4385) );
  OAI222_X1 U1681 ( .A1(n15078), .A2(n13029), .B1(n15014), .B2(n13026), .C1(
        n15046), .C2(n13023), .ZN(n4388) );
  AOI221_X1 U1682 ( .B1(n12981), .B2(n15430), .C1(n12978), .C2(n15398), .A(
        n4414), .ZN(n4411) );
  OAI222_X1 U1683 ( .A1(n15526), .A2(n12975), .B1(n15462), .B2(n12972), .C1(
        n15494), .C2(n12969), .ZN(n4414) );
  AOI221_X1 U1684 ( .B1(n13087), .B2(n14691), .C1(n13084), .C2(n15765), .A(
        n5689), .ZN(n5688) );
  OAI222_X1 U1685 ( .A1(n14787), .A2(n13081), .B1(n14723), .B2(n13078), .C1(
        n14755), .C2(n13075), .ZN(n5689) );
  AOI221_X1 U1686 ( .B1(n12979), .B2(n15461), .C1(n12976), .C2(n15429), .A(
        n5728), .ZN(n5726) );
  OAI222_X1 U1687 ( .A1(n15557), .A2(n12973), .B1(n15493), .B2(n12970), .C1(
        n15525), .C2(n12967), .ZN(n5728) );
  AOI221_X1 U1688 ( .B1(n13087), .B2(n14690), .C1(n13084), .C2(n15764), .A(
        n5609), .ZN(n5608) );
  OAI222_X1 U1689 ( .A1(n14786), .A2(n13081), .B1(n14722), .B2(n13078), .C1(
        n14754), .C2(n13075), .ZN(n5609) );
  AOI221_X1 U1690 ( .B1(n12979), .B2(n15460), .C1(n12976), .C2(n15428), .A(
        n5636), .ZN(n5634) );
  OAI222_X1 U1691 ( .A1(n15556), .A2(n12973), .B1(n15492), .B2(n12970), .C1(
        n15524), .C2(n12967), .ZN(n5636) );
  AOI221_X1 U1692 ( .B1(n13087), .B2(n14689), .C1(n13084), .C2(n15763), .A(
        n5548), .ZN(n5546) );
  OAI222_X1 U1693 ( .A1(n14785), .A2(n13081), .B1(n14721), .B2(n13078), .C1(
        n14753), .C2(n13075), .ZN(n5548) );
  AOI221_X1 U1694 ( .B1(n12979), .B2(n15459), .C1(n12976), .C2(n15427), .A(
        n5574), .ZN(n5571) );
  OAI222_X1 U1695 ( .A1(n15555), .A2(n12973), .B1(n15491), .B2(n12970), .C1(
        n15523), .C2(n12967), .ZN(n5574) );
  AOI221_X1 U1696 ( .B1(n13087), .B2(n14688), .C1(n13084), .C2(n15762), .A(
        n5486), .ZN(n5484) );
  OAI222_X1 U1697 ( .A1(n14784), .A2(n13081), .B1(n14720), .B2(n13078), .C1(
        n14752), .C2(n13075), .ZN(n5486) );
  AOI221_X1 U1698 ( .B1(n12979), .B2(n15458), .C1(n12976), .C2(n15426), .A(
        n5511), .ZN(n5510) );
  OAI222_X1 U1699 ( .A1(n15554), .A2(n12973), .B1(n15490), .B2(n12970), .C1(
        n15522), .C2(n12967), .ZN(n5511) );
  AOI221_X1 U1700 ( .B1(n13087), .B2(n14687), .C1(n13084), .C2(n15761), .A(
        n5428), .ZN(n5426) );
  OAI222_X1 U1701 ( .A1(n14783), .A2(n13081), .B1(n14719), .B2(n13078), .C1(
        n14751), .C2(n13075), .ZN(n5428) );
  AOI221_X1 U1702 ( .B1(n12979), .B2(n15457), .C1(n12976), .C2(n15425), .A(
        n5450), .ZN(n5449) );
  OAI222_X1 U1703 ( .A1(n15553), .A2(n12973), .B1(n15489), .B2(n12970), .C1(
        n15521), .C2(n12967), .ZN(n5450) );
  AOI221_X1 U1704 ( .B1(n13087), .B2(n14686), .C1(n13084), .C2(n15760), .A(
        n5376), .ZN(n5375) );
  OAI222_X1 U1705 ( .A1(n14782), .A2(n13081), .B1(n14718), .B2(n13078), .C1(
        n14750), .C2(n13075), .ZN(n5376) );
  AOI221_X1 U1706 ( .B1(n12979), .B2(n15456), .C1(n12976), .C2(n15424), .A(
        n5398), .ZN(n5396) );
  OAI222_X1 U1707 ( .A1(n15552), .A2(n12973), .B1(n15488), .B2(n12970), .C1(
        n15520), .C2(n12967), .ZN(n5398) );
  AOI221_X1 U1708 ( .B1(n13087), .B2(n14685), .C1(n13084), .C2(n15759), .A(
        n5339), .ZN(n5338) );
  OAI222_X1 U1709 ( .A1(n14781), .A2(n13081), .B1(n14717), .B2(n13078), .C1(
        n14749), .C2(n13075), .ZN(n5339) );
  AOI221_X1 U1710 ( .B1(n12979), .B2(n15455), .C1(n12976), .C2(n15423), .A(
        n5355), .ZN(n5354) );
  OAI222_X1 U1711 ( .A1(n15551), .A2(n12973), .B1(n15487), .B2(n12970), .C1(
        n15519), .C2(n12967), .ZN(n5355) );
  AOI221_X1 U1712 ( .B1(n13087), .B2(n14684), .C1(n13084), .C2(n15758), .A(
        n5302), .ZN(n5301) );
  OAI222_X1 U1713 ( .A1(n14780), .A2(n13081), .B1(n14716), .B2(n13078), .C1(
        n14748), .C2(n13075), .ZN(n5302) );
  AOI221_X1 U1714 ( .B1(n12979), .B2(n15454), .C1(n12976), .C2(n15422), .A(
        n5318), .ZN(n5317) );
  OAI222_X1 U1715 ( .A1(n15550), .A2(n12973), .B1(n15486), .B2(n12970), .C1(
        n15518), .C2(n12967), .ZN(n5318) );
  AOI221_X1 U1716 ( .B1(n13087), .B2(n14683), .C1(n13084), .C2(n15757), .A(
        n5265), .ZN(n5264) );
  OAI222_X1 U1717 ( .A1(n14779), .A2(n13081), .B1(n14715), .B2(n13078), .C1(
        n14747), .C2(n13075), .ZN(n5265) );
  AOI221_X1 U1718 ( .B1(n12979), .B2(n15453), .C1(n12976), .C2(n15421), .A(
        n5281), .ZN(n5280) );
  OAI222_X1 U1719 ( .A1(n15549), .A2(n12973), .B1(n15485), .B2(n12970), .C1(
        n15517), .C2(n12967), .ZN(n5281) );
  AOI221_X1 U1720 ( .B1(n13087), .B2(n14682), .C1(n13084), .C2(n15756), .A(
        n5228), .ZN(n5227) );
  OAI222_X1 U1721 ( .A1(n14778), .A2(n13081), .B1(n14714), .B2(n13078), .C1(
        n14746), .C2(n13075), .ZN(n5228) );
  AOI221_X1 U1722 ( .B1(n12979), .B2(n15452), .C1(n12976), .C2(n15420), .A(
        n5244), .ZN(n5243) );
  OAI222_X1 U1723 ( .A1(n15548), .A2(n12973), .B1(n15484), .B2(n12970), .C1(
        n15516), .C2(n12967), .ZN(n5244) );
  AOI221_X1 U1724 ( .B1(n13087), .B2(n14681), .C1(n13084), .C2(n15755), .A(
        n5191), .ZN(n5190) );
  OAI222_X1 U1725 ( .A1(n14777), .A2(n13081), .B1(n14713), .B2(n13078), .C1(
        n14745), .C2(n13075), .ZN(n5191) );
  AOI221_X1 U1726 ( .B1(n12979), .B2(n15451), .C1(n12976), .C2(n15419), .A(
        n5207), .ZN(n5206) );
  OAI222_X1 U1727 ( .A1(n15547), .A2(n12973), .B1(n15483), .B2(n12970), .C1(
        n15515), .C2(n12967), .ZN(n5207) );
  AOI221_X1 U1728 ( .B1(n13087), .B2(n14680), .C1(n13084), .C2(n15754), .A(
        n5154), .ZN(n5153) );
  OAI222_X1 U1729 ( .A1(n14776), .A2(n13081), .B1(n14712), .B2(n13078), .C1(
        n14744), .C2(n13075), .ZN(n5154) );
  AOI221_X1 U1730 ( .B1(n12979), .B2(n15450), .C1(n12976), .C2(n15418), .A(
        n5170), .ZN(n5169) );
  OAI222_X1 U1731 ( .A1(n15546), .A2(n12973), .B1(n15482), .B2(n12970), .C1(
        n15514), .C2(n12967), .ZN(n5170) );
  AOI221_X1 U1732 ( .B1(n13142), .B2(n14267), .C1(n13139), .C2(n15885), .A(
        n5109), .ZN(n5108) );
  OAI222_X1 U1733 ( .A1(n14363), .A2(n13136), .B1(n14299), .B2(n13133), .C1(
        n14331), .C2(n13130), .ZN(n5109) );
  AOI221_X1 U1734 ( .B1(n13088), .B2(n14679), .C1(n13085), .C2(n15753), .A(
        n5117), .ZN(n5116) );
  OAI222_X1 U1735 ( .A1(n14775), .A2(n13082), .B1(n14711), .B2(n13079), .C1(
        n14743), .C2(n13076), .ZN(n5117) );
  AOI221_X1 U1736 ( .B1(n13034), .B2(n15001), .C1(n13031), .C2(n15653), .A(
        n5125), .ZN(n5124) );
  OAI222_X1 U1737 ( .A1(n15097), .A2(n13028), .B1(n15033), .B2(n13025), .C1(
        n15065), .C2(n13022), .ZN(n5125) );
  AOI221_X1 U1738 ( .B1(n13142), .B2(n14266), .C1(n13139), .C2(n15884), .A(
        n5072), .ZN(n5071) );
  OAI222_X1 U1739 ( .A1(n14362), .A2(n13136), .B1(n14298), .B2(n13133), .C1(
        n14330), .C2(n13130), .ZN(n5072) );
  AOI221_X1 U1740 ( .B1(n13088), .B2(n14678), .C1(n13085), .C2(n15752), .A(
        n5080), .ZN(n5079) );
  OAI222_X1 U1741 ( .A1(n14774), .A2(n13082), .B1(n14710), .B2(n13079), .C1(
        n14742), .C2(n13076), .ZN(n5080) );
  AOI221_X1 U1742 ( .B1(n13034), .B2(n15000), .C1(n13031), .C2(n15652), .A(
        n5088), .ZN(n5087) );
  OAI222_X1 U1743 ( .A1(n15096), .A2(n13028), .B1(n15032), .B2(n13025), .C1(
        n15064), .C2(n13022), .ZN(n5088) );
  AOI221_X1 U1744 ( .B1(n13142), .B2(n14265), .C1(n13139), .C2(n15883), .A(
        n5035), .ZN(n5034) );
  OAI222_X1 U1745 ( .A1(n14361), .A2(n13136), .B1(n14297), .B2(n13133), .C1(
        n14329), .C2(n13130), .ZN(n5035) );
  AOI221_X1 U1746 ( .B1(n13088), .B2(n14677), .C1(n13085), .C2(n15751), .A(
        n5043), .ZN(n5042) );
  OAI222_X1 U1747 ( .A1(n14773), .A2(n13082), .B1(n14709), .B2(n13079), .C1(
        n14741), .C2(n13076), .ZN(n5043) );
  AOI221_X1 U1748 ( .B1(n13034), .B2(n14999), .C1(n13031), .C2(n15651), .A(
        n5051), .ZN(n5050) );
  OAI222_X1 U1749 ( .A1(n15095), .A2(n13028), .B1(n15031), .B2(n13025), .C1(
        n15063), .C2(n13022), .ZN(n5051) );
  AOI221_X1 U1750 ( .B1(n13142), .B2(n14264), .C1(n13139), .C2(n15882), .A(
        n4998), .ZN(n4997) );
  OAI222_X1 U1751 ( .A1(n14360), .A2(n13136), .B1(n14296), .B2(n13133), .C1(
        n14328), .C2(n13130), .ZN(n4998) );
  AOI221_X1 U1752 ( .B1(n13088), .B2(n14676), .C1(n13085), .C2(n15750), .A(
        n5006), .ZN(n5005) );
  OAI222_X1 U1753 ( .A1(n14772), .A2(n13082), .B1(n14708), .B2(n13079), .C1(
        n14740), .C2(n13076), .ZN(n5006) );
  AOI221_X1 U1754 ( .B1(n13034), .B2(n14998), .C1(n13031), .C2(n15650), .A(
        n5014), .ZN(n5013) );
  OAI222_X1 U1755 ( .A1(n15094), .A2(n13028), .B1(n15030), .B2(n13025), .C1(
        n15062), .C2(n13022), .ZN(n5014) );
  AOI221_X1 U1756 ( .B1(n13142), .B2(n14263), .C1(n13139), .C2(n15881), .A(
        n4961), .ZN(n4960) );
  OAI222_X1 U1757 ( .A1(n14359), .A2(n13136), .B1(n14295), .B2(n13133), .C1(
        n14327), .C2(n13130), .ZN(n4961) );
  AOI221_X1 U1758 ( .B1(n13088), .B2(n14675), .C1(n13085), .C2(n15749), .A(
        n4969), .ZN(n4968) );
  OAI222_X1 U1759 ( .A1(n14771), .A2(n13082), .B1(n14707), .B2(n13079), .C1(
        n14739), .C2(n13076), .ZN(n4969) );
  AOI221_X1 U1760 ( .B1(n13034), .B2(n14997), .C1(n13031), .C2(n15649), .A(
        n4977), .ZN(n4976) );
  OAI222_X1 U1761 ( .A1(n15093), .A2(n13028), .B1(n15029), .B2(n13025), .C1(
        n15061), .C2(n13022), .ZN(n4977) );
  AOI221_X1 U1762 ( .B1(n13142), .B2(n14262), .C1(n13139), .C2(n15880), .A(
        n4924), .ZN(n4923) );
  OAI222_X1 U1763 ( .A1(n14358), .A2(n13136), .B1(n14294), .B2(n13133), .C1(
        n14326), .C2(n13130), .ZN(n4924) );
  AOI221_X1 U1764 ( .B1(n13088), .B2(n14674), .C1(n13085), .C2(n15748), .A(
        n4932), .ZN(n4931) );
  OAI222_X1 U1765 ( .A1(n14770), .A2(n13082), .B1(n14706), .B2(n13079), .C1(
        n14738), .C2(n13076), .ZN(n4932) );
  AOI221_X1 U1766 ( .B1(n13034), .B2(n14996), .C1(n13031), .C2(n15648), .A(
        n4940), .ZN(n4939) );
  OAI222_X1 U1767 ( .A1(n15092), .A2(n13028), .B1(n15028), .B2(n13025), .C1(
        n15060), .C2(n13022), .ZN(n4940) );
  AOI221_X1 U1768 ( .B1(n13142), .B2(n14261), .C1(n13139), .C2(n15879), .A(
        n4887), .ZN(n4886) );
  OAI222_X1 U1769 ( .A1(n14357), .A2(n13136), .B1(n14293), .B2(n13133), .C1(
        n14325), .C2(n13130), .ZN(n4887) );
  AOI221_X1 U1770 ( .B1(n13088), .B2(n14673), .C1(n13085), .C2(n15747), .A(
        n4895), .ZN(n4894) );
  OAI222_X1 U1771 ( .A1(n14769), .A2(n13082), .B1(n14705), .B2(n13079), .C1(
        n14737), .C2(n13076), .ZN(n4895) );
  AOI221_X1 U1772 ( .B1(n13034), .B2(n14995), .C1(n13031), .C2(n15647), .A(
        n4903), .ZN(n4902) );
  OAI222_X1 U1773 ( .A1(n15091), .A2(n13028), .B1(n15027), .B2(n13025), .C1(
        n15059), .C2(n13022), .ZN(n4903) );
  AOI221_X1 U1774 ( .B1(n13142), .B2(n14260), .C1(n13139), .C2(n15878), .A(
        n4850), .ZN(n4849) );
  OAI222_X1 U1775 ( .A1(n14356), .A2(n13136), .B1(n14292), .B2(n13133), .C1(
        n14324), .C2(n13130), .ZN(n4850) );
  AOI221_X1 U1776 ( .B1(n13088), .B2(n14672), .C1(n13085), .C2(n15746), .A(
        n4858), .ZN(n4857) );
  OAI222_X1 U1777 ( .A1(n14768), .A2(n13082), .B1(n14704), .B2(n13079), .C1(
        n14736), .C2(n13076), .ZN(n4858) );
  AOI221_X1 U1778 ( .B1(n13034), .B2(n14994), .C1(n13031), .C2(n15646), .A(
        n4866), .ZN(n4865) );
  OAI222_X1 U1779 ( .A1(n15090), .A2(n13028), .B1(n15026), .B2(n13025), .C1(
        n15058), .C2(n13022), .ZN(n4866) );
  AOI221_X1 U1780 ( .B1(n13142), .B2(n14259), .C1(n13139), .C2(n15877), .A(
        n4813), .ZN(n4812) );
  OAI222_X1 U1781 ( .A1(n14355), .A2(n13136), .B1(n14291), .B2(n13133), .C1(
        n14323), .C2(n13130), .ZN(n4813) );
  AOI221_X1 U1782 ( .B1(n13088), .B2(n14671), .C1(n13085), .C2(n15745), .A(
        n4821), .ZN(n4820) );
  OAI222_X1 U1783 ( .A1(n14767), .A2(n13082), .B1(n14703), .B2(n13079), .C1(
        n14735), .C2(n13076), .ZN(n4821) );
  AOI221_X1 U1784 ( .B1(n13142), .B2(n14258), .C1(n13139), .C2(n15876), .A(
        n4776), .ZN(n4775) );
  OAI222_X1 U1785 ( .A1(n14354), .A2(n13136), .B1(n14290), .B2(n13133), .C1(
        n14322), .C2(n13130), .ZN(n4776) );
  AOI221_X1 U1786 ( .B1(n13088), .B2(n14670), .C1(n13085), .C2(n15744), .A(
        n4784), .ZN(n4783) );
  OAI222_X1 U1787 ( .A1(n14766), .A2(n13082), .B1(n14702), .B2(n13079), .C1(
        n14734), .C2(n13076), .ZN(n4784) );
  AOI221_X1 U1788 ( .B1(n13142), .B2(n14257), .C1(n13139), .C2(n15875), .A(
        n4739), .ZN(n4738) );
  OAI222_X1 U1789 ( .A1(n14353), .A2(n13136), .B1(n14289), .B2(n13133), .C1(
        n14321), .C2(n13130), .ZN(n4739) );
  AOI221_X1 U1790 ( .B1(n13088), .B2(n14669), .C1(n13085), .C2(n15743), .A(
        n4747), .ZN(n4746) );
  OAI222_X1 U1791 ( .A1(n14765), .A2(n13082), .B1(n14701), .B2(n13079), .C1(
        n14733), .C2(n13076), .ZN(n4747) );
  AOI221_X1 U1792 ( .B1(n13142), .B2(n14256), .C1(n13139), .C2(n15874), .A(
        n4702), .ZN(n4701) );
  OAI222_X1 U1793 ( .A1(n14352), .A2(n13136), .B1(n14288), .B2(n13133), .C1(
        n14320), .C2(n13130), .ZN(n4702) );
  AOI221_X1 U1794 ( .B1(n13088), .B2(n14668), .C1(n13085), .C2(n15742), .A(
        n4710), .ZN(n4709) );
  OAI222_X1 U1795 ( .A1(n14764), .A2(n13082), .B1(n14700), .B2(n13079), .C1(
        n14732), .C2(n13076), .ZN(n4710) );
  AOI221_X1 U1796 ( .B1(n13143), .B2(n14255), .C1(n13140), .C2(n15597), .A(
        n4665), .ZN(n4664) );
  OAI222_X1 U1797 ( .A1(n14351), .A2(n13137), .B1(n14287), .B2(n13134), .C1(
        n14319), .C2(n13131), .ZN(n4665) );
  AOI221_X1 U1798 ( .B1(n13089), .B2(n14667), .C1(n13086), .C2(n15573), .A(
        n4673), .ZN(n4672) );
  OAI222_X1 U1799 ( .A1(n14763), .A2(n13083), .B1(n14699), .B2(n13080), .C1(
        n14731), .C2(n13077), .ZN(n4673) );
  AOI221_X1 U1800 ( .B1(n13035), .B2(n14989), .C1(n13032), .C2(n15641), .A(
        n4681), .ZN(n4680) );
  OAI222_X1 U1801 ( .A1(n15085), .A2(n13029), .B1(n15021), .B2(n13026), .C1(
        n15053), .C2(n13023), .ZN(n4681) );
  AOI221_X1 U1802 ( .B1(n12981), .B2(n15437), .C1(n12978), .C2(n15405), .A(
        n4689), .ZN(n4688) );
  OAI222_X1 U1803 ( .A1(n15533), .A2(n12975), .B1(n15469), .B2(n12972), .C1(
        n15501), .C2(n12969), .ZN(n4689) );
  AOI221_X1 U1804 ( .B1(n13315), .B2(n14691), .C1(n13312), .C2(n15765), .A(
        n4288), .ZN(n4287) );
  OAI222_X1 U1805 ( .A1(n14787), .A2(n13309), .B1(n14723), .B2(n13306), .C1(
        n14755), .C2(n13303), .ZN(n4288) );
  AOI221_X1 U1806 ( .B1(n13207), .B2(n15461), .C1(n13204), .C2(n15429), .A(
        n4308), .ZN(n4307) );
  OAI222_X1 U1807 ( .A1(n15557), .A2(n13201), .B1(n15493), .B2(n13198), .C1(
        n15525), .C2(n13195), .ZN(n4308) );
  AOI221_X1 U1808 ( .B1(n13315), .B2(n14690), .C1(n13312), .C2(n15764), .A(
        n4240), .ZN(n4239) );
  OAI222_X1 U1809 ( .A1(n14786), .A2(n13309), .B1(n14722), .B2(n13306), .C1(
        n14754), .C2(n13303), .ZN(n4240) );
  AOI221_X1 U1810 ( .B1(n13207), .B2(n15460), .C1(n13204), .C2(n15428), .A(
        n4256), .ZN(n4255) );
  OAI222_X1 U1811 ( .A1(n15556), .A2(n13201), .B1(n15492), .B2(n13198), .C1(
        n15524), .C2(n13195), .ZN(n4256) );
  AOI221_X1 U1812 ( .B1(n13315), .B2(n14689), .C1(n13312), .C2(n15763), .A(
        n4203), .ZN(n4202) );
  OAI222_X1 U1813 ( .A1(n14785), .A2(n13309), .B1(n14721), .B2(n13306), .C1(
        n14753), .C2(n13303), .ZN(n4203) );
  AOI221_X1 U1814 ( .B1(n13207), .B2(n15459), .C1(n13204), .C2(n15427), .A(
        n4219), .ZN(n4218) );
  OAI222_X1 U1815 ( .A1(n15555), .A2(n13201), .B1(n15491), .B2(n13198), .C1(
        n15523), .C2(n13195), .ZN(n4219) );
  AOI221_X1 U1816 ( .B1(n13315), .B2(n14688), .C1(n13312), .C2(n15762), .A(
        n4166), .ZN(n4165) );
  OAI222_X1 U1817 ( .A1(n14784), .A2(n13309), .B1(n14720), .B2(n13306), .C1(
        n14752), .C2(n13303), .ZN(n4166) );
  AOI221_X1 U1818 ( .B1(n13207), .B2(n15458), .C1(n13204), .C2(n15426), .A(
        n4182), .ZN(n4181) );
  OAI222_X1 U1819 ( .A1(n15554), .A2(n13201), .B1(n15490), .B2(n13198), .C1(
        n15522), .C2(n13195), .ZN(n4182) );
  AOI221_X1 U1820 ( .B1(n13315), .B2(n14687), .C1(n13312), .C2(n15761), .A(
        n4129), .ZN(n4128) );
  OAI222_X1 U1821 ( .A1(n14783), .A2(n13309), .B1(n14719), .B2(n13306), .C1(
        n14751), .C2(n13303), .ZN(n4129) );
  AOI221_X1 U1822 ( .B1(n13207), .B2(n15457), .C1(n13204), .C2(n15425), .A(
        n4145), .ZN(n4144) );
  OAI222_X1 U1823 ( .A1(n15553), .A2(n13201), .B1(n15489), .B2(n13198), .C1(
        n15521), .C2(n13195), .ZN(n4145) );
  AOI221_X1 U1824 ( .B1(n13315), .B2(n14686), .C1(n13312), .C2(n15760), .A(
        n4092), .ZN(n4091) );
  OAI222_X1 U1825 ( .A1(n14782), .A2(n13309), .B1(n14718), .B2(n13306), .C1(
        n14750), .C2(n13303), .ZN(n4092) );
  AOI221_X1 U1826 ( .B1(n13207), .B2(n15456), .C1(n13204), .C2(n15424), .A(
        n4108), .ZN(n4107) );
  OAI222_X1 U1827 ( .A1(n15552), .A2(n13201), .B1(n15488), .B2(n13198), .C1(
        n15520), .C2(n13195), .ZN(n4108) );
  AOI221_X1 U1828 ( .B1(n13315), .B2(n14685), .C1(n13312), .C2(n15759), .A(
        n4055), .ZN(n4054) );
  OAI222_X1 U1829 ( .A1(n14781), .A2(n13309), .B1(n14717), .B2(n13306), .C1(
        n14749), .C2(n13303), .ZN(n4055) );
  AOI221_X1 U1830 ( .B1(n13207), .B2(n15455), .C1(n13204), .C2(n15423), .A(
        n4071), .ZN(n4070) );
  OAI222_X1 U1831 ( .A1(n15551), .A2(n13201), .B1(n15487), .B2(n13198), .C1(
        n15519), .C2(n13195), .ZN(n4071) );
  AOI221_X1 U1832 ( .B1(n13315), .B2(n14684), .C1(n13312), .C2(n15758), .A(
        n4018), .ZN(n4017) );
  OAI222_X1 U1833 ( .A1(n14780), .A2(n13309), .B1(n14716), .B2(n13306), .C1(
        n14748), .C2(n13303), .ZN(n4018) );
  AOI221_X1 U1834 ( .B1(n13207), .B2(n15454), .C1(n13204), .C2(n15422), .A(
        n4034), .ZN(n4033) );
  OAI222_X1 U1835 ( .A1(n15550), .A2(n13201), .B1(n15486), .B2(n13198), .C1(
        n15518), .C2(n13195), .ZN(n4034) );
  AOI221_X1 U1836 ( .B1(n13315), .B2(n14683), .C1(n13312), .C2(n15757), .A(
        n3981), .ZN(n3980) );
  OAI222_X1 U1837 ( .A1(n14779), .A2(n13309), .B1(n14715), .B2(n13306), .C1(
        n14747), .C2(n13303), .ZN(n3981) );
  AOI221_X1 U1838 ( .B1(n13207), .B2(n15453), .C1(n13204), .C2(n15421), .A(
        n3997), .ZN(n3996) );
  OAI222_X1 U1839 ( .A1(n15549), .A2(n13201), .B1(n15485), .B2(n13198), .C1(
        n15517), .C2(n13195), .ZN(n3997) );
  AOI221_X1 U1840 ( .B1(n13315), .B2(n14682), .C1(n13312), .C2(n15756), .A(
        n3944), .ZN(n3943) );
  OAI222_X1 U1841 ( .A1(n14778), .A2(n13309), .B1(n14714), .B2(n13306), .C1(
        n14746), .C2(n13303), .ZN(n3944) );
  AOI221_X1 U1842 ( .B1(n13207), .B2(n15452), .C1(n13204), .C2(n15420), .A(
        n3960), .ZN(n3959) );
  OAI222_X1 U1843 ( .A1(n15548), .A2(n13201), .B1(n15484), .B2(n13198), .C1(
        n15516), .C2(n13195), .ZN(n3960) );
  AOI221_X1 U1844 ( .B1(n13315), .B2(n14681), .C1(n13312), .C2(n15755), .A(
        n3907), .ZN(n3906) );
  OAI222_X1 U1845 ( .A1(n14777), .A2(n13309), .B1(n14713), .B2(n13306), .C1(
        n14745), .C2(n13303), .ZN(n3907) );
  AOI221_X1 U1846 ( .B1(n13207), .B2(n15451), .C1(n13204), .C2(n15419), .A(
        n3923), .ZN(n3922) );
  OAI222_X1 U1847 ( .A1(n15547), .A2(n13201), .B1(n15483), .B2(n13198), .C1(
        n15515), .C2(n13195), .ZN(n3923) );
  AOI221_X1 U1848 ( .B1(n13315), .B2(n14680), .C1(n13312), .C2(n15754), .A(
        n3870), .ZN(n3869) );
  OAI222_X1 U1849 ( .A1(n14776), .A2(n13309), .B1(n14712), .B2(n13306), .C1(
        n14744), .C2(n13303), .ZN(n3870) );
  AOI221_X1 U1850 ( .B1(n13207), .B2(n15450), .C1(n13204), .C2(n15418), .A(
        n3886), .ZN(n3885) );
  OAI222_X1 U1851 ( .A1(n15546), .A2(n13201), .B1(n15482), .B2(n13198), .C1(
        n15514), .C2(n13195), .ZN(n3886) );
  AOI221_X1 U1852 ( .B1(n13370), .B2(n14267), .C1(n13367), .C2(n15885), .A(
        n3825), .ZN(n3824) );
  OAI222_X1 U1853 ( .A1(n14363), .A2(n13364), .B1(n14299), .B2(n13361), .C1(
        n14331), .C2(n13358), .ZN(n3825) );
  AOI221_X1 U1854 ( .B1(n13316), .B2(n14679), .C1(n13313), .C2(n15753), .A(
        n3833), .ZN(n3832) );
  OAI222_X1 U1855 ( .A1(n14775), .A2(n13310), .B1(n14711), .B2(n13307), .C1(
        n14743), .C2(n13304), .ZN(n3833) );
  AOI221_X1 U1856 ( .B1(n13262), .B2(n15001), .C1(n13259), .C2(n15653), .A(
        n3841), .ZN(n3840) );
  OAI222_X1 U1857 ( .A1(n15097), .A2(n13256), .B1(n15033), .B2(n13253), .C1(
        n15065), .C2(n13250), .ZN(n3841) );
  AOI221_X1 U1858 ( .B1(n13370), .B2(n14266), .C1(n13367), .C2(n15884), .A(
        n3788), .ZN(n3787) );
  OAI222_X1 U1859 ( .A1(n14362), .A2(n13364), .B1(n14298), .B2(n13361), .C1(
        n14330), .C2(n13358), .ZN(n3788) );
  AOI221_X1 U1860 ( .B1(n13316), .B2(n14678), .C1(n13313), .C2(n15752), .A(
        n3796), .ZN(n3795) );
  OAI222_X1 U1861 ( .A1(n14774), .A2(n13310), .B1(n14710), .B2(n13307), .C1(
        n14742), .C2(n13304), .ZN(n3796) );
  AOI221_X1 U1862 ( .B1(n13262), .B2(n15000), .C1(n13259), .C2(n15652), .A(
        n3804), .ZN(n3803) );
  OAI222_X1 U1863 ( .A1(n15096), .A2(n13256), .B1(n15032), .B2(n13253), .C1(
        n15064), .C2(n13250), .ZN(n3804) );
  AOI221_X1 U1864 ( .B1(n13370), .B2(n14265), .C1(n13367), .C2(n15883), .A(
        n3751), .ZN(n3750) );
  OAI222_X1 U1865 ( .A1(n14361), .A2(n13364), .B1(n14297), .B2(n13361), .C1(
        n14329), .C2(n13358), .ZN(n3751) );
  AOI221_X1 U1866 ( .B1(n13316), .B2(n14677), .C1(n13313), .C2(n15751), .A(
        n3759), .ZN(n3758) );
  OAI222_X1 U1867 ( .A1(n14773), .A2(n13310), .B1(n14709), .B2(n13307), .C1(
        n14741), .C2(n13304), .ZN(n3759) );
  AOI221_X1 U1868 ( .B1(n13262), .B2(n14999), .C1(n13259), .C2(n15651), .A(
        n3767), .ZN(n3766) );
  OAI222_X1 U1869 ( .A1(n15095), .A2(n13256), .B1(n15031), .B2(n13253), .C1(
        n15063), .C2(n13250), .ZN(n3767) );
  AOI221_X1 U1870 ( .B1(n13370), .B2(n14264), .C1(n13367), .C2(n15882), .A(
        n3714), .ZN(n3713) );
  OAI222_X1 U1871 ( .A1(n14360), .A2(n13364), .B1(n14296), .B2(n13361), .C1(
        n14328), .C2(n13358), .ZN(n3714) );
  AOI221_X1 U1872 ( .B1(n13316), .B2(n14676), .C1(n13313), .C2(n15750), .A(
        n3722), .ZN(n3721) );
  OAI222_X1 U1873 ( .A1(n14772), .A2(n13310), .B1(n14708), .B2(n13307), .C1(
        n14740), .C2(n13304), .ZN(n3722) );
  AOI221_X1 U1874 ( .B1(n13262), .B2(n14998), .C1(n13259), .C2(n15650), .A(
        n3730), .ZN(n3729) );
  OAI222_X1 U1875 ( .A1(n15094), .A2(n13256), .B1(n15030), .B2(n13253), .C1(
        n15062), .C2(n13250), .ZN(n3730) );
  AOI221_X1 U1876 ( .B1(n13370), .B2(n14263), .C1(n13367), .C2(n15881), .A(
        n3677), .ZN(n3676) );
  OAI222_X1 U1877 ( .A1(n14359), .A2(n13364), .B1(n14295), .B2(n13361), .C1(
        n14327), .C2(n13358), .ZN(n3677) );
  AOI221_X1 U1878 ( .B1(n13316), .B2(n14675), .C1(n13313), .C2(n15749), .A(
        n3685), .ZN(n3684) );
  OAI222_X1 U1879 ( .A1(n14771), .A2(n13310), .B1(n14707), .B2(n13307), .C1(
        n14739), .C2(n13304), .ZN(n3685) );
  AOI221_X1 U1880 ( .B1(n13262), .B2(n14997), .C1(n13259), .C2(n15649), .A(
        n3693), .ZN(n3692) );
  OAI222_X1 U1881 ( .A1(n15093), .A2(n13256), .B1(n15029), .B2(n13253), .C1(
        n15061), .C2(n13250), .ZN(n3693) );
  AOI221_X1 U1882 ( .B1(n13370), .B2(n14262), .C1(n13367), .C2(n15880), .A(
        n3640), .ZN(n3639) );
  OAI222_X1 U1883 ( .A1(n14358), .A2(n13364), .B1(n14294), .B2(n13361), .C1(
        n14326), .C2(n13358), .ZN(n3640) );
  AOI221_X1 U1884 ( .B1(n13316), .B2(n14674), .C1(n13313), .C2(n15748), .A(
        n3648), .ZN(n3647) );
  OAI222_X1 U1885 ( .A1(n14770), .A2(n13310), .B1(n14706), .B2(n13307), .C1(
        n14738), .C2(n13304), .ZN(n3648) );
  AOI221_X1 U1886 ( .B1(n13262), .B2(n14996), .C1(n13259), .C2(n15648), .A(
        n3656), .ZN(n3655) );
  OAI222_X1 U1887 ( .A1(n15092), .A2(n13256), .B1(n15028), .B2(n13253), .C1(
        n15060), .C2(n13250), .ZN(n3656) );
  AOI221_X1 U1888 ( .B1(n13370), .B2(n14261), .C1(n13367), .C2(n15879), .A(
        n3603), .ZN(n3602) );
  OAI222_X1 U1889 ( .A1(n14357), .A2(n13364), .B1(n14293), .B2(n13361), .C1(
        n14325), .C2(n13358), .ZN(n3603) );
  AOI221_X1 U1890 ( .B1(n13316), .B2(n14673), .C1(n13313), .C2(n15747), .A(
        n3611), .ZN(n3610) );
  OAI222_X1 U1891 ( .A1(n14769), .A2(n13310), .B1(n14705), .B2(n13307), .C1(
        n14737), .C2(n13304), .ZN(n3611) );
  AOI221_X1 U1892 ( .B1(n13262), .B2(n14995), .C1(n13259), .C2(n15647), .A(
        n3619), .ZN(n3618) );
  OAI222_X1 U1893 ( .A1(n15091), .A2(n13256), .B1(n15027), .B2(n13253), .C1(
        n15059), .C2(n13250), .ZN(n3619) );
  AOI221_X1 U1894 ( .B1(n13370), .B2(n14260), .C1(n13367), .C2(n15878), .A(
        n3566), .ZN(n3565) );
  OAI222_X1 U1895 ( .A1(n14356), .A2(n13364), .B1(n14292), .B2(n13361), .C1(
        n14324), .C2(n13358), .ZN(n3566) );
  AOI221_X1 U1896 ( .B1(n13316), .B2(n14672), .C1(n13313), .C2(n15746), .A(
        n3574), .ZN(n3573) );
  OAI222_X1 U1897 ( .A1(n14768), .A2(n13310), .B1(n14704), .B2(n13307), .C1(
        n14736), .C2(n13304), .ZN(n3574) );
  AOI221_X1 U1898 ( .B1(n13262), .B2(n14994), .C1(n13259), .C2(n15646), .A(
        n3582), .ZN(n3581) );
  OAI222_X1 U1899 ( .A1(n15090), .A2(n13256), .B1(n15026), .B2(n13253), .C1(
        n15058), .C2(n13250), .ZN(n3582) );
  AOI221_X1 U1900 ( .B1(n13370), .B2(n14259), .C1(n13367), .C2(n15877), .A(
        n3529), .ZN(n3528) );
  OAI222_X1 U1901 ( .A1(n14355), .A2(n13364), .B1(n14291), .B2(n13361), .C1(
        n14323), .C2(n13358), .ZN(n3529) );
  AOI221_X1 U1902 ( .B1(n13316), .B2(n14671), .C1(n13313), .C2(n15745), .A(
        n3537), .ZN(n3536) );
  OAI222_X1 U1903 ( .A1(n14767), .A2(n13310), .B1(n14703), .B2(n13307), .C1(
        n14735), .C2(n13304), .ZN(n3537) );
  AOI221_X1 U1904 ( .B1(n13370), .B2(n14258), .C1(n13367), .C2(n15876), .A(
        n3492), .ZN(n3491) );
  OAI222_X1 U1905 ( .A1(n14354), .A2(n13364), .B1(n14290), .B2(n13361), .C1(
        n14322), .C2(n13358), .ZN(n3492) );
  AOI221_X1 U1906 ( .B1(n13316), .B2(n14670), .C1(n13313), .C2(n15744), .A(
        n3500), .ZN(n3499) );
  OAI222_X1 U1907 ( .A1(n14766), .A2(n13310), .B1(n14702), .B2(n13307), .C1(
        n14734), .C2(n13304), .ZN(n3500) );
  AOI221_X1 U1908 ( .B1(n13370), .B2(n14257), .C1(n13367), .C2(n15875), .A(
        n3455), .ZN(n3454) );
  OAI222_X1 U1909 ( .A1(n14353), .A2(n13364), .B1(n14289), .B2(n13361), .C1(
        n14321), .C2(n13358), .ZN(n3455) );
  AOI221_X1 U1910 ( .B1(n13316), .B2(n14669), .C1(n13313), .C2(n15743), .A(
        n3463), .ZN(n3462) );
  OAI222_X1 U1911 ( .A1(n14765), .A2(n13310), .B1(n14701), .B2(n13307), .C1(
        n14733), .C2(n13304), .ZN(n3463) );
  AOI221_X1 U1912 ( .B1(n13370), .B2(n14256), .C1(n13367), .C2(n15874), .A(
        n3418), .ZN(n3417) );
  OAI222_X1 U1913 ( .A1(n14352), .A2(n13364), .B1(n14288), .B2(n13361), .C1(
        n14320), .C2(n13358), .ZN(n3418) );
  AOI221_X1 U1914 ( .B1(n13316), .B2(n14668), .C1(n13313), .C2(n15742), .A(
        n3426), .ZN(n3425) );
  OAI222_X1 U1915 ( .A1(n14764), .A2(n13310), .B1(n14700), .B2(n13307), .C1(
        n14732), .C2(n13304), .ZN(n3426) );
  AOI221_X1 U1916 ( .B1(n13371), .B2(n14255), .C1(n13368), .C2(n15597), .A(
        n3381), .ZN(n3380) );
  OAI222_X1 U1917 ( .A1(n14351), .A2(n13365), .B1(n14287), .B2(n13362), .C1(
        n14319), .C2(n13359), .ZN(n3381) );
  AOI221_X1 U1918 ( .B1(n13317), .B2(n14667), .C1(n13314), .C2(n15573), .A(
        n3389), .ZN(n3388) );
  OAI222_X1 U1919 ( .A1(n14763), .A2(n13311), .B1(n14699), .B2(n13308), .C1(
        n14731), .C2(n13305), .ZN(n3389) );
  AOI221_X1 U1920 ( .B1(n13263), .B2(n14989), .C1(n13260), .C2(n15641), .A(
        n3397), .ZN(n3396) );
  OAI222_X1 U1921 ( .A1(n15085), .A2(n13257), .B1(n15021), .B2(n13254), .C1(
        n15053), .C2(n13251), .ZN(n3397) );
  AOI221_X1 U1922 ( .B1(n13209), .B2(n15437), .C1(n13206), .C2(n15405), .A(
        n3405), .ZN(n3404) );
  OAI222_X1 U1923 ( .A1(n15533), .A2(n13203), .B1(n15469), .B2(n13200), .C1(
        n15501), .C2(n13197), .ZN(n3405) );
  AOI221_X1 U1924 ( .B1(n13371), .B2(n14254), .C1(n13368), .C2(n15596), .A(
        n3344), .ZN(n3343) );
  OAI222_X1 U1925 ( .A1(n14350), .A2(n13365), .B1(n14286), .B2(n13362), .C1(
        n14318), .C2(n13359), .ZN(n3344) );
  AOI221_X1 U1926 ( .B1(n13317), .B2(n14666), .C1(n13314), .C2(n15572), .A(
        n3352), .ZN(n3351) );
  OAI222_X1 U1927 ( .A1(n14762), .A2(n13311), .B1(n14698), .B2(n13308), .C1(
        n14730), .C2(n13305), .ZN(n3352) );
  AOI221_X1 U1928 ( .B1(n13263), .B2(n14988), .C1(n13260), .C2(n15640), .A(
        n3360), .ZN(n3359) );
  OAI222_X1 U1929 ( .A1(n15084), .A2(n13257), .B1(n15020), .B2(n13254), .C1(
        n15052), .C2(n13251), .ZN(n3360) );
  AOI221_X1 U1930 ( .B1(n13209), .B2(n15436), .C1(n13206), .C2(n15404), .A(
        n3368), .ZN(n3367) );
  OAI222_X1 U1931 ( .A1(n15532), .A2(n13203), .B1(n15468), .B2(n13200), .C1(
        n15500), .C2(n13197), .ZN(n3368) );
  AOI221_X1 U1932 ( .B1(n13371), .B2(n14253), .C1(n13368), .C2(n15595), .A(
        n3307), .ZN(n3306) );
  OAI222_X1 U1933 ( .A1(n14349), .A2(n13365), .B1(n14285), .B2(n13362), .C1(
        n14317), .C2(n13359), .ZN(n3307) );
  AOI221_X1 U1934 ( .B1(n13317), .B2(n14665), .C1(n13314), .C2(n15571), .A(
        n3315), .ZN(n3314) );
  OAI222_X1 U1935 ( .A1(n14761), .A2(n13311), .B1(n14697), .B2(n13308), .C1(
        n14729), .C2(n13305), .ZN(n3315) );
  AOI221_X1 U1936 ( .B1(n13263), .B2(n14987), .C1(n13260), .C2(n15639), .A(
        n3323), .ZN(n3322) );
  OAI222_X1 U1937 ( .A1(n15083), .A2(n13257), .B1(n15019), .B2(n13254), .C1(
        n15051), .C2(n13251), .ZN(n3323) );
  AOI221_X1 U1938 ( .B1(n13209), .B2(n15435), .C1(n13206), .C2(n15403), .A(
        n3331), .ZN(n3330) );
  OAI222_X1 U1939 ( .A1(n15531), .A2(n13203), .B1(n15467), .B2(n13200), .C1(
        n15499), .C2(n13197), .ZN(n3331) );
  AOI221_X1 U1940 ( .B1(n13371), .B2(n14252), .C1(n13368), .C2(n15594), .A(
        n3270), .ZN(n3269) );
  OAI222_X1 U1941 ( .A1(n14348), .A2(n13365), .B1(n14284), .B2(n13362), .C1(
        n14316), .C2(n13359), .ZN(n3270) );
  AOI221_X1 U1942 ( .B1(n13317), .B2(n14664), .C1(n13314), .C2(n15570), .A(
        n3278), .ZN(n3277) );
  OAI222_X1 U1943 ( .A1(n14760), .A2(n13311), .B1(n14696), .B2(n13308), .C1(
        n14728), .C2(n13305), .ZN(n3278) );
  AOI221_X1 U1944 ( .B1(n13263), .B2(n14986), .C1(n13260), .C2(n15638), .A(
        n3286), .ZN(n3285) );
  OAI222_X1 U1945 ( .A1(n15082), .A2(n13257), .B1(n15018), .B2(n13254), .C1(
        n15050), .C2(n13251), .ZN(n3286) );
  AOI221_X1 U1946 ( .B1(n13209), .B2(n15434), .C1(n13206), .C2(n15402), .A(
        n3294), .ZN(n3293) );
  OAI222_X1 U1947 ( .A1(n15530), .A2(n13203), .B1(n15466), .B2(n13200), .C1(
        n15498), .C2(n13197), .ZN(n3294) );
  AOI221_X1 U1948 ( .B1(n13221), .B2(n15733), .C1(n13218), .C2(n15622), .A(
        n3252), .ZN(n3245) );
  OAI22_X1 U1949 ( .A1(n14823), .A2(n13215), .B1(n14791), .B2(n13212), .ZN(
        n3252) );
  AOI221_X1 U1950 ( .B1(n13221), .B2(n15732), .C1(n13218), .C2(n15621), .A(
        n3215), .ZN(n3208) );
  OAI22_X1 U1951 ( .A1(n14822), .A2(n13215), .B1(n14790), .B2(n13212), .ZN(
        n3215) );
  AOI221_X1 U1952 ( .B1(n13221), .B2(n15731), .C1(n13218), .C2(n15620), .A(
        n3178), .ZN(n3171) );
  OAI22_X1 U1953 ( .A1(n14821), .A2(n13215), .B1(n14789), .B2(n13212), .ZN(
        n3178) );
  AOI221_X1 U1954 ( .B1(n12993), .B2(n15736), .C1(n12990), .C2(n15625), .A(
        n4647), .ZN(n4640) );
  OAI22_X1 U1955 ( .A1(n14826), .A2(n12987), .B1(n14794), .B2(n12984), .ZN(
        n4647) );
  AOI221_X1 U1956 ( .B1(n12993), .B2(n15735), .C1(n12990), .C2(n15624), .A(
        n4610), .ZN(n4603) );
  OAI22_X1 U1957 ( .A1(n14825), .A2(n12987), .B1(n14793), .B2(n12984), .ZN(
        n4610) );
  AOI221_X1 U1958 ( .B1(n12993), .B2(n15734), .C1(n12990), .C2(n15623), .A(
        n4573), .ZN(n4566) );
  OAI22_X1 U1959 ( .A1(n14824), .A2(n12987), .B1(n14792), .B2(n12984), .ZN(
        n4573) );
  AOI221_X1 U1960 ( .B1(n12993), .B2(n15733), .C1(n12990), .C2(n15622), .A(
        n4536), .ZN(n4529) );
  OAI22_X1 U1961 ( .A1(n14823), .A2(n12987), .B1(n14791), .B2(n12984), .ZN(
        n4536) );
  AOI221_X1 U1962 ( .B1(n12993), .B2(n15732), .C1(n12990), .C2(n15621), .A(
        n4499), .ZN(n4492) );
  OAI22_X1 U1963 ( .A1(n14822), .A2(n12987), .B1(n14790), .B2(n12984), .ZN(
        n4499) );
  AOI221_X1 U1964 ( .B1(n12993), .B2(n15731), .C1(n12990), .C2(n15620), .A(
        n4462), .ZN(n4455) );
  OAI22_X1 U1965 ( .A1(n14821), .A2(n12987), .B1(n14789), .B2(n12984), .ZN(
        n4462) );
  AOI221_X1 U1966 ( .B1(n12993), .B2(n15737), .C1(n12990), .C2(n15626), .A(
        n4684), .ZN(n4677) );
  OAI22_X1 U1967 ( .A1(n14827), .A2(n12987), .B1(n14795), .B2(n12984), .ZN(
        n4684) );
  AOI221_X1 U1968 ( .B1(n13221), .B2(n15737), .C1(n13218), .C2(n15626), .A(
        n3400), .ZN(n3393) );
  OAI22_X1 U1969 ( .A1(n14827), .A2(n13215), .B1(n14795), .B2(n13212), .ZN(
        n3400) );
  AOI221_X1 U1970 ( .B1(n13221), .B2(n15736), .C1(n13218), .C2(n15625), .A(
        n3363), .ZN(n3356) );
  OAI22_X1 U1971 ( .A1(n14826), .A2(n13215), .B1(n14794), .B2(n13212), .ZN(
        n3363) );
  AOI221_X1 U1972 ( .B1(n13221), .B2(n15735), .C1(n13218), .C2(n15624), .A(
        n3326), .ZN(n3319) );
  OAI22_X1 U1973 ( .A1(n14825), .A2(n13215), .B1(n14793), .B2(n13212), .ZN(
        n3326) );
  AOI221_X1 U1974 ( .B1(n13221), .B2(n15734), .C1(n13218), .C2(n15623), .A(
        n3289), .ZN(n3282) );
  OAI22_X1 U1975 ( .A1(n14824), .A2(n13215), .B1(n14792), .B2(n13212), .ZN(
        n3289) );
  OAI22_X1 U1976 ( .A1(n14592), .A2(n13296), .B1(n14624), .B2(n13293), .ZN(
        n3242) );
  OAI22_X1 U1977 ( .A1(n14411), .A2(n13269), .B1(n14379), .B2(n13266), .ZN(
        n3244) );
  OAI22_X1 U1978 ( .A1(n14591), .A2(n13296), .B1(n14623), .B2(n13293), .ZN(
        n3205) );
  OAI22_X1 U1979 ( .A1(n14410), .A2(n13269), .B1(n14378), .B2(n13266), .ZN(
        n3207) );
  OAI22_X1 U1980 ( .A1(n14590), .A2(n13296), .B1(n14622), .B2(n13293), .ZN(
        n3168) );
  OAI22_X1 U1981 ( .A1(n14409), .A2(n13269), .B1(n14377), .B2(n13266), .ZN(
        n3170) );
  OAI22_X1 U1982 ( .A1(n14589), .A2(n13296), .B1(n14621), .B2(n13293), .ZN(
        n3084) );
  OAI22_X1 U1983 ( .A1(n14408), .A2(n13269), .B1(n14376), .B2(n13266), .ZN(
        n3095) );
  OAI22_X1 U1984 ( .A1(n14627), .A2(n13068), .B1(n14595), .B2(n13065), .ZN(
        n4637) );
  OAI22_X1 U1985 ( .A1(n14414), .A2(n13041), .B1(n14382), .B2(n13038), .ZN(
        n4639) );
  OAI22_X1 U1986 ( .A1(n14626), .A2(n13068), .B1(n14594), .B2(n13065), .ZN(
        n4600) );
  OAI22_X1 U1987 ( .A1(n14413), .A2(n13041), .B1(n14381), .B2(n13038), .ZN(
        n4602) );
  OAI22_X1 U1988 ( .A1(n14625), .A2(n13068), .B1(n14593), .B2(n13065), .ZN(
        n4563) );
  OAI22_X1 U1989 ( .A1(n14412), .A2(n13041), .B1(n14380), .B2(n13038), .ZN(
        n4565) );
  OAI22_X1 U1990 ( .A1(n14624), .A2(n13068), .B1(n14592), .B2(n13065), .ZN(
        n4526) );
  OAI22_X1 U1991 ( .A1(n14411), .A2(n13041), .B1(n14379), .B2(n13038), .ZN(
        n4528) );
  OAI22_X1 U1992 ( .A1(n14623), .A2(n13068), .B1(n14591), .B2(n13065), .ZN(
        n4489) );
  OAI22_X1 U1993 ( .A1(n14410), .A2(n13041), .B1(n14378), .B2(n13038), .ZN(
        n4491) );
  OAI22_X1 U1994 ( .A1(n14622), .A2(n13068), .B1(n14590), .B2(n13065), .ZN(
        n4452) );
  OAI22_X1 U1995 ( .A1(n14409), .A2(n13041), .B1(n14377), .B2(n13038), .ZN(
        n4454) );
  OAI22_X1 U1996 ( .A1(n14621), .A2(n13068), .B1(n14589), .B2(n13065), .ZN(
        n4368) );
  OAI22_X1 U1997 ( .A1(n14408), .A2(n13041), .B1(n14376), .B2(n13038), .ZN(
        n4379) );
  OAI22_X1 U1998 ( .A1(n14628), .A2(n13068), .B1(n14596), .B2(n13065), .ZN(
        n4674) );
  OAI22_X1 U1999 ( .A1(n14415), .A2(n13041), .B1(n14383), .B2(n13038), .ZN(
        n4676) );
  OAI22_X1 U2000 ( .A1(n14596), .A2(n13296), .B1(n14628), .B2(n13293), .ZN(
        n3390) );
  OAI22_X1 U2001 ( .A1(n14415), .A2(n13269), .B1(n14383), .B2(n13266), .ZN(
        n3392) );
  OAI22_X1 U2002 ( .A1(n14595), .A2(n13296), .B1(n14627), .B2(n13293), .ZN(
        n3353) );
  OAI22_X1 U2003 ( .A1(n14414), .A2(n13269), .B1(n14382), .B2(n13266), .ZN(
        n3355) );
  OAI22_X1 U2004 ( .A1(n14594), .A2(n13296), .B1(n14626), .B2(n13293), .ZN(
        n3316) );
  OAI22_X1 U2005 ( .A1(n14413), .A2(n13269), .B1(n14381), .B2(n13266), .ZN(
        n3318) );
  OAI22_X1 U2006 ( .A1(n14593), .A2(n13296), .B1(n14625), .B2(n13293), .ZN(
        n3279) );
  OAI22_X1 U2007 ( .A1(n14412), .A2(n13269), .B1(n14380), .B2(n13266), .ZN(
        n3281) );
  OAI22_X1 U2008 ( .A1(n14652), .A2(n13066), .B1(n14620), .B2(n13063), .ZN(
        n5694) );
  OAI22_X1 U2009 ( .A1(n14439), .A2(n13039), .B1(n14407), .B2(n13036), .ZN(
        n5698) );
  OAI22_X1 U2010 ( .A1(n14651), .A2(n13066), .B1(n14619), .B2(n13063), .ZN(
        n5610) );
  OAI22_X1 U2011 ( .A1(n14438), .A2(n13039), .B1(n14406), .B2(n13036), .ZN(
        n5614) );
  OAI22_X1 U2012 ( .A1(n14650), .A2(n13066), .B1(n14618), .B2(n13063), .ZN(
        n5549) );
  OAI22_X1 U2013 ( .A1(n14437), .A2(n13039), .B1(n14405), .B2(n13036), .ZN(
        n5551) );
  OAI22_X1 U2014 ( .A1(n14649), .A2(n13066), .B1(n14617), .B2(n13063), .ZN(
        n5488) );
  OAI22_X1 U2015 ( .A1(n14436), .A2(n13039), .B1(n14404), .B2(n13036), .ZN(
        n5490) );
  OAI22_X1 U2016 ( .A1(n14648), .A2(n13066), .B1(n14616), .B2(n13063), .ZN(
        n5429) );
  OAI22_X1 U2017 ( .A1(n14435), .A2(n13039), .B1(n14403), .B2(n13036), .ZN(
        n5431) );
  OAI22_X1 U2018 ( .A1(n14647), .A2(n13066), .B1(n14615), .B2(n13063), .ZN(
        n5377) );
  OAI22_X1 U2019 ( .A1(n14434), .A2(n13039), .B1(n14402), .B2(n13036), .ZN(
        n5379) );
  OAI22_X1 U2020 ( .A1(n14646), .A2(n13066), .B1(n14614), .B2(n13063), .ZN(
        n5340) );
  OAI22_X1 U2021 ( .A1(n14433), .A2(n13039), .B1(n14401), .B2(n13036), .ZN(
        n5342) );
  OAI22_X1 U2022 ( .A1(n14645), .A2(n13066), .B1(n14613), .B2(n13063), .ZN(
        n5303) );
  OAI22_X1 U2023 ( .A1(n14432), .A2(n13039), .B1(n14400), .B2(n13036), .ZN(
        n5305) );
  OAI22_X1 U2024 ( .A1(n14644), .A2(n13066), .B1(n14612), .B2(n13063), .ZN(
        n5266) );
  OAI22_X1 U2025 ( .A1(n14431), .A2(n13039), .B1(n14399), .B2(n13036), .ZN(
        n5268) );
  OAI22_X1 U2026 ( .A1(n14643), .A2(n13066), .B1(n14611), .B2(n13063), .ZN(
        n5229) );
  OAI22_X1 U2027 ( .A1(n14430), .A2(n13039), .B1(n14398), .B2(n13036), .ZN(
        n5231) );
  OAI22_X1 U2028 ( .A1(n14642), .A2(n13066), .B1(n14610), .B2(n13063), .ZN(
        n5192) );
  OAI22_X1 U2029 ( .A1(n14429), .A2(n13039), .B1(n14397), .B2(n13036), .ZN(
        n5194) );
  OAI22_X1 U2030 ( .A1(n14641), .A2(n13066), .B1(n14609), .B2(n13063), .ZN(
        n5155) );
  OAI22_X1 U2031 ( .A1(n14428), .A2(n13039), .B1(n14396), .B2(n13036), .ZN(
        n5157) );
  OAI22_X1 U2032 ( .A1(n14640), .A2(n13067), .B1(n14608), .B2(n13064), .ZN(
        n5118) );
  OAI22_X1 U2033 ( .A1(n14427), .A2(n13040), .B1(n14395), .B2(n13037), .ZN(
        n5120) );
  OAI22_X1 U2034 ( .A1(n14639), .A2(n13067), .B1(n14607), .B2(n13064), .ZN(
        n5081) );
  OAI22_X1 U2035 ( .A1(n14426), .A2(n13040), .B1(n14394), .B2(n13037), .ZN(
        n5083) );
  OAI22_X1 U2036 ( .A1(n14638), .A2(n13067), .B1(n14606), .B2(n13064), .ZN(
        n5044) );
  OAI22_X1 U2037 ( .A1(n14425), .A2(n13040), .B1(n14393), .B2(n13037), .ZN(
        n5046) );
  OAI22_X1 U2038 ( .A1(n14637), .A2(n13067), .B1(n14605), .B2(n13064), .ZN(
        n5007) );
  OAI22_X1 U2039 ( .A1(n14424), .A2(n13040), .B1(n14392), .B2(n13037), .ZN(
        n5009) );
  OAI22_X1 U2040 ( .A1(n14636), .A2(n13067), .B1(n14604), .B2(n13064), .ZN(
        n4970) );
  OAI22_X1 U2041 ( .A1(n14423), .A2(n13040), .B1(n14391), .B2(n13037), .ZN(
        n4972) );
  OAI22_X1 U2042 ( .A1(n14635), .A2(n13067), .B1(n14603), .B2(n13064), .ZN(
        n4933) );
  OAI22_X1 U2043 ( .A1(n14422), .A2(n13040), .B1(n14390), .B2(n13037), .ZN(
        n4935) );
  OAI22_X1 U2044 ( .A1(n14634), .A2(n13067), .B1(n14602), .B2(n13064), .ZN(
        n4896) );
  OAI22_X1 U2045 ( .A1(n14421), .A2(n13040), .B1(n14389), .B2(n13037), .ZN(
        n4898) );
  OAI22_X1 U2046 ( .A1(n14633), .A2(n13067), .B1(n14601), .B2(n13064), .ZN(
        n4859) );
  OAI22_X1 U2047 ( .A1(n14420), .A2(n13040), .B1(n14388), .B2(n13037), .ZN(
        n4861) );
  OAI22_X1 U2048 ( .A1(n14632), .A2(n13067), .B1(n14600), .B2(n13064), .ZN(
        n4822) );
  OAI22_X1 U2049 ( .A1(n14419), .A2(n13040), .B1(n14387), .B2(n13037), .ZN(
        n4824) );
  OAI22_X1 U2050 ( .A1(n14631), .A2(n13067), .B1(n14599), .B2(n13064), .ZN(
        n4785) );
  OAI22_X1 U2051 ( .A1(n14418), .A2(n13040), .B1(n14386), .B2(n13037), .ZN(
        n4787) );
  OAI22_X1 U2052 ( .A1(n14630), .A2(n13067), .B1(n14598), .B2(n13064), .ZN(
        n4748) );
  OAI22_X1 U2053 ( .A1(n14417), .A2(n13040), .B1(n14385), .B2(n13037), .ZN(
        n4750) );
  OAI22_X1 U2054 ( .A1(n14629), .A2(n13067), .B1(n14597), .B2(n13064), .ZN(
        n4711) );
  OAI22_X1 U2055 ( .A1(n14416), .A2(n13040), .B1(n14384), .B2(n13037), .ZN(
        n4713) );
  OAI22_X1 U2056 ( .A1(n14620), .A2(n13294), .B1(n14652), .B2(n13291), .ZN(
        n4291) );
  OAI22_X1 U2057 ( .A1(n14439), .A2(n13267), .B1(n14407), .B2(n13264), .ZN(
        n4293) );
  OAI22_X1 U2058 ( .A1(n14619), .A2(n13294), .B1(n14651), .B2(n13291), .ZN(
        n4241) );
  OAI22_X1 U2059 ( .A1(n14438), .A2(n13267), .B1(n14406), .B2(n13264), .ZN(
        n4243) );
  OAI22_X1 U2060 ( .A1(n14618), .A2(n13294), .B1(n14650), .B2(n13291), .ZN(
        n4204) );
  OAI22_X1 U2061 ( .A1(n14437), .A2(n13267), .B1(n14405), .B2(n13264), .ZN(
        n4206) );
  OAI22_X1 U2062 ( .A1(n14617), .A2(n13294), .B1(n14649), .B2(n13291), .ZN(
        n4167) );
  OAI22_X1 U2063 ( .A1(n14436), .A2(n13267), .B1(n14404), .B2(n13264), .ZN(
        n4169) );
  OAI22_X1 U2064 ( .A1(n14616), .A2(n13294), .B1(n14648), .B2(n13291), .ZN(
        n4130) );
  OAI22_X1 U2065 ( .A1(n14435), .A2(n13267), .B1(n14403), .B2(n13264), .ZN(
        n4132) );
  OAI22_X1 U2066 ( .A1(n14615), .A2(n13294), .B1(n14647), .B2(n13291), .ZN(
        n4093) );
  OAI22_X1 U2067 ( .A1(n14434), .A2(n13267), .B1(n14402), .B2(n13264), .ZN(
        n4095) );
  OAI22_X1 U2068 ( .A1(n14614), .A2(n13294), .B1(n14646), .B2(n13291), .ZN(
        n4056) );
  OAI22_X1 U2069 ( .A1(n14433), .A2(n13267), .B1(n14401), .B2(n13264), .ZN(
        n4058) );
  OAI22_X1 U2070 ( .A1(n14613), .A2(n13294), .B1(n14645), .B2(n13291), .ZN(
        n4019) );
  OAI22_X1 U2071 ( .A1(n14432), .A2(n13267), .B1(n14400), .B2(n13264), .ZN(
        n4021) );
  OAI22_X1 U2072 ( .A1(n14612), .A2(n13294), .B1(n14644), .B2(n13291), .ZN(
        n3982) );
  OAI22_X1 U2073 ( .A1(n14431), .A2(n13267), .B1(n14399), .B2(n13264), .ZN(
        n3984) );
  OAI22_X1 U2074 ( .A1(n14611), .A2(n13294), .B1(n14643), .B2(n13291), .ZN(
        n3945) );
  OAI22_X1 U2075 ( .A1(n14430), .A2(n13267), .B1(n14398), .B2(n13264), .ZN(
        n3947) );
  OAI22_X1 U2076 ( .A1(n14610), .A2(n13294), .B1(n14642), .B2(n13291), .ZN(
        n3908) );
  OAI22_X1 U2077 ( .A1(n14429), .A2(n13267), .B1(n14397), .B2(n13264), .ZN(
        n3910) );
  OAI22_X1 U2078 ( .A1(n14609), .A2(n13294), .B1(n14641), .B2(n13291), .ZN(
        n3871) );
  OAI22_X1 U2079 ( .A1(n14428), .A2(n13267), .B1(n14396), .B2(n13264), .ZN(
        n3873) );
  OAI22_X1 U2080 ( .A1(n14608), .A2(n13295), .B1(n14640), .B2(n13292), .ZN(
        n3834) );
  OAI22_X1 U2081 ( .A1(n14427), .A2(n13268), .B1(n14395), .B2(n13265), .ZN(
        n3836) );
  OAI22_X1 U2082 ( .A1(n14607), .A2(n13295), .B1(n14639), .B2(n13292), .ZN(
        n3797) );
  OAI22_X1 U2083 ( .A1(n14426), .A2(n13268), .B1(n14394), .B2(n13265), .ZN(
        n3799) );
  OAI22_X1 U2084 ( .A1(n14606), .A2(n13295), .B1(n14638), .B2(n13292), .ZN(
        n3760) );
  OAI22_X1 U2085 ( .A1(n14425), .A2(n13268), .B1(n14393), .B2(n13265), .ZN(
        n3762) );
  OAI22_X1 U2086 ( .A1(n14605), .A2(n13295), .B1(n14637), .B2(n13292), .ZN(
        n3723) );
  OAI22_X1 U2087 ( .A1(n14424), .A2(n13268), .B1(n14392), .B2(n13265), .ZN(
        n3725) );
  OAI22_X1 U2088 ( .A1(n14604), .A2(n13295), .B1(n14636), .B2(n13292), .ZN(
        n3686) );
  OAI22_X1 U2089 ( .A1(n14423), .A2(n13268), .B1(n14391), .B2(n13265), .ZN(
        n3688) );
  OAI22_X1 U2090 ( .A1(n14603), .A2(n13295), .B1(n14635), .B2(n13292), .ZN(
        n3649) );
  OAI22_X1 U2091 ( .A1(n14422), .A2(n13268), .B1(n14390), .B2(n13265), .ZN(
        n3651) );
  OAI22_X1 U2092 ( .A1(n14602), .A2(n13295), .B1(n14634), .B2(n13292), .ZN(
        n3612) );
  OAI22_X1 U2093 ( .A1(n14421), .A2(n13268), .B1(n14389), .B2(n13265), .ZN(
        n3614) );
  OAI22_X1 U2094 ( .A1(n14601), .A2(n13295), .B1(n14633), .B2(n13292), .ZN(
        n3575) );
  OAI22_X1 U2095 ( .A1(n14420), .A2(n13268), .B1(n14388), .B2(n13265), .ZN(
        n3577) );
  OAI22_X1 U2096 ( .A1(n14600), .A2(n13295), .B1(n14632), .B2(n13292), .ZN(
        n3538) );
  OAI22_X1 U2097 ( .A1(n14419), .A2(n13268), .B1(n14387), .B2(n13265), .ZN(
        n3540) );
  OAI22_X1 U2098 ( .A1(n14599), .A2(n13295), .B1(n14631), .B2(n13292), .ZN(
        n3501) );
  OAI22_X1 U2099 ( .A1(n14418), .A2(n13268), .B1(n14386), .B2(n13265), .ZN(
        n3503) );
  OAI22_X1 U2100 ( .A1(n14598), .A2(n13295), .B1(n14630), .B2(n13292), .ZN(
        n3464) );
  OAI22_X1 U2101 ( .A1(n14417), .A2(n13268), .B1(n14385), .B2(n13265), .ZN(
        n3466) );
  OAI22_X1 U2102 ( .A1(n14597), .A2(n13295), .B1(n14629), .B2(n13292), .ZN(
        n3427) );
  OAI22_X1 U2103 ( .A1(n14416), .A2(n13268), .B1(n14384), .B2(n13265), .ZN(
        n3429) );
  AOI221_X1 U2104 ( .B1(n12992), .B2(n15741), .C1(n12989), .C2(n15709), .A(
        n4832), .ZN(n4825) );
  OAI22_X1 U2105 ( .A1(n14831), .A2(n12986), .B1(n14799), .B2(n12983), .ZN(
        n4832) );
  AOI221_X1 U2106 ( .B1(n12992), .B2(n15740), .C1(n12989), .C2(n15708), .A(
        n4795), .ZN(n4788) );
  OAI22_X1 U2107 ( .A1(n14830), .A2(n12986), .B1(n14798), .B2(n12983), .ZN(
        n4795) );
  AOI221_X1 U2108 ( .B1(n12992), .B2(n15739), .C1(n12989), .C2(n15707), .A(
        n4758), .ZN(n4751) );
  OAI22_X1 U2109 ( .A1(n14829), .A2(n12986), .B1(n14797), .B2(n12983), .ZN(
        n4758) );
  AOI221_X1 U2110 ( .B1(n12992), .B2(n15738), .C1(n12989), .C2(n15706), .A(
        n4721), .ZN(n4714) );
  OAI22_X1 U2111 ( .A1(n14828), .A2(n12986), .B1(n14796), .B2(n12983), .ZN(
        n4721) );
  AOI221_X1 U2112 ( .B1(n13220), .B2(n15741), .C1(n13217), .C2(n15709), .A(
        n3548), .ZN(n3541) );
  OAI22_X1 U2113 ( .A1(n14831), .A2(n13214), .B1(n14799), .B2(n13211), .ZN(
        n3548) );
  AOI221_X1 U2114 ( .B1(n13220), .B2(n15740), .C1(n13217), .C2(n15708), .A(
        n3511), .ZN(n3504) );
  OAI22_X1 U2115 ( .A1(n14830), .A2(n13214), .B1(n14798), .B2(n13211), .ZN(
        n3511) );
  AOI221_X1 U2116 ( .B1(n13220), .B2(n15739), .C1(n13217), .C2(n15707), .A(
        n3474), .ZN(n3467) );
  OAI22_X1 U2117 ( .A1(n14829), .A2(n13214), .B1(n14797), .B2(n13211), .ZN(
        n3474) );
  AOI221_X1 U2118 ( .B1(n13220), .B2(n15738), .C1(n13217), .C2(n15706), .A(
        n3437), .ZN(n3430) );
  OAI22_X1 U2119 ( .A1(n14828), .A2(n13214), .B1(n14796), .B2(n13211), .ZN(
        n3437) );
  OAI22_X1 U2120 ( .A1(n13829), .A2(n13384), .B1(n13387), .B2(n15557), .ZN(
        n7674) );
  OAI22_X1 U2121 ( .A1(n13829), .A2(n13395), .B1(n13390), .B2(n15525), .ZN(
        n7706) );
  OAI22_X1 U2122 ( .A1(n13829), .A2(n13401), .B1(n13396), .B2(n15493), .ZN(
        n7738) );
  OAI22_X1 U2123 ( .A1(n13835), .A2(n13401), .B1(n13396), .B2(n15492), .ZN(
        n7739) );
  OAI22_X1 U2124 ( .A1(n13841), .A2(n13401), .B1(n13396), .B2(n15491), .ZN(
        n7740) );
  OAI22_X1 U2125 ( .A1(n13847), .A2(n13401), .B1(n13396), .B2(n15490), .ZN(
        n7741) );
  OAI22_X1 U2126 ( .A1(n13853), .A2(n13401), .B1(n13396), .B2(n15489), .ZN(
        n7742) );
  OAI22_X1 U2127 ( .A1(n13859), .A2(n13401), .B1(n13396), .B2(n15488), .ZN(
        n7743) );
  OAI22_X1 U2128 ( .A1(n13865), .A2(n13401), .B1(n13396), .B2(n15487), .ZN(
        n7744) );
  OAI22_X1 U2129 ( .A1(n13871), .A2(n13401), .B1(n13396), .B2(n15486), .ZN(
        n7745) );
  OAI22_X1 U2130 ( .A1(n13877), .A2(n13400), .B1(n13396), .B2(n15485), .ZN(
        n7746) );
  OAI22_X1 U2131 ( .A1(n13883), .A2(n13400), .B1(n13396), .B2(n15484), .ZN(
        n7747) );
  OAI22_X1 U2132 ( .A1(n13889), .A2(n13400), .B1(n13396), .B2(n15483), .ZN(
        n7748) );
  OAI22_X1 U2133 ( .A1(n13895), .A2(n13400), .B1(n13396), .B2(n15482), .ZN(
        n7749) );
  OAI22_X1 U2134 ( .A1(n13901), .A2(n13400), .B1(n13397), .B2(n15481), .ZN(
        n7750) );
  OAI22_X1 U2135 ( .A1(n13907), .A2(n13400), .B1(n13397), .B2(n15480), .ZN(
        n7751) );
  OAI22_X1 U2136 ( .A1(n13913), .A2(n13400), .B1(n13397), .B2(n15479), .ZN(
        n7752) );
  OAI22_X1 U2137 ( .A1(n13919), .A2(n13400), .B1(n13397), .B2(n15478), .ZN(
        n7753) );
  OAI22_X1 U2138 ( .A1(n13925), .A2(n13400), .B1(n13397), .B2(n15477), .ZN(
        n7754) );
  OAI22_X1 U2139 ( .A1(n13931), .A2(n13400), .B1(n13397), .B2(n15476), .ZN(
        n7755) );
  OAI22_X1 U2140 ( .A1(n13937), .A2(n13400), .B1(n13397), .B2(n15475), .ZN(
        n7756) );
  OAI22_X1 U2141 ( .A1(n13943), .A2(n13400), .B1(n13397), .B2(n15474), .ZN(
        n7757) );
  OAI22_X1 U2142 ( .A1(n13949), .A2(n13399), .B1(n13397), .B2(n15473), .ZN(
        n7758) );
  OAI22_X1 U2143 ( .A1(n13955), .A2(n13399), .B1(n13397), .B2(n15472), .ZN(
        n7759) );
  OAI22_X1 U2144 ( .A1(n13961), .A2(n13399), .B1(n13397), .B2(n15471), .ZN(
        n7760) );
  OAI22_X1 U2145 ( .A1(n13967), .A2(n13399), .B1(n13397), .B2(n15470), .ZN(
        n7761) );
  OAI22_X1 U2146 ( .A1(n13973), .A2(n13399), .B1(n13398), .B2(n15469), .ZN(
        n7762) );
  OAI22_X1 U2147 ( .A1(n13979), .A2(n13399), .B1(n13398), .B2(n15468), .ZN(
        n7763) );
  OAI22_X1 U2148 ( .A1(n13985), .A2(n13399), .B1(n13398), .B2(n15467), .ZN(
        n7764) );
  OAI22_X1 U2149 ( .A1(n13991), .A2(n13399), .B1(n13398), .B2(n15466), .ZN(
        n7765) );
  OAI22_X1 U2150 ( .A1(n13997), .A2(n13399), .B1(n13398), .B2(n15465), .ZN(
        n7766) );
  OAI22_X1 U2151 ( .A1(n14003), .A2(n13399), .B1(n13398), .B2(n15464), .ZN(
        n7767) );
  OAI22_X1 U2152 ( .A1(n14009), .A2(n13399), .B1(n13398), .B2(n15463), .ZN(
        n7768) );
  OAI22_X1 U2153 ( .A1(n14018), .A2(n13399), .B1(n13398), .B2(n15462), .ZN(
        n7769) );
  OAI22_X1 U2154 ( .A1(n13829), .A2(n13419), .B1(n13414), .B2(n15397), .ZN(
        n7834) );
  OAI22_X1 U2155 ( .A1(n13835), .A2(n13419), .B1(n13414), .B2(n15396), .ZN(
        n7835) );
  OAI22_X1 U2156 ( .A1(n13841), .A2(n13419), .B1(n13414), .B2(n15395), .ZN(
        n7836) );
  OAI22_X1 U2157 ( .A1(n13847), .A2(n13419), .B1(n13414), .B2(n15394), .ZN(
        n7837) );
  OAI22_X1 U2158 ( .A1(n13853), .A2(n13419), .B1(n13414), .B2(n15393), .ZN(
        n7838) );
  OAI22_X1 U2159 ( .A1(n13859), .A2(n13419), .B1(n13414), .B2(n15392), .ZN(
        n7839) );
  OAI22_X1 U2160 ( .A1(n13865), .A2(n13419), .B1(n13414), .B2(n15391), .ZN(
        n7840) );
  OAI22_X1 U2161 ( .A1(n13871), .A2(n13419), .B1(n13414), .B2(n15390), .ZN(
        n7841) );
  OAI22_X1 U2162 ( .A1(n13877), .A2(n13418), .B1(n13414), .B2(n15389), .ZN(
        n7842) );
  OAI22_X1 U2163 ( .A1(n13883), .A2(n13418), .B1(n13414), .B2(n15388), .ZN(
        n7843) );
  OAI22_X1 U2164 ( .A1(n13889), .A2(n13418), .B1(n13414), .B2(n15387), .ZN(
        n7844) );
  OAI22_X1 U2165 ( .A1(n13895), .A2(n13418), .B1(n13414), .B2(n15386), .ZN(
        n7845) );
  OAI22_X1 U2166 ( .A1(n13901), .A2(n13418), .B1(n13415), .B2(n15385), .ZN(
        n7846) );
  OAI22_X1 U2167 ( .A1(n13907), .A2(n13418), .B1(n13415), .B2(n15384), .ZN(
        n7847) );
  OAI22_X1 U2168 ( .A1(n13913), .A2(n13418), .B1(n13415), .B2(n15383), .ZN(
        n7848) );
  OAI22_X1 U2169 ( .A1(n13919), .A2(n13418), .B1(n13415), .B2(n15382), .ZN(
        n7849) );
  OAI22_X1 U2170 ( .A1(n13925), .A2(n13418), .B1(n13415), .B2(n15381), .ZN(
        n7850) );
  OAI22_X1 U2171 ( .A1(n13931), .A2(n13418), .B1(n13415), .B2(n15380), .ZN(
        n7851) );
  OAI22_X1 U2172 ( .A1(n13937), .A2(n13418), .B1(n13415), .B2(n15379), .ZN(
        n7852) );
  OAI22_X1 U2173 ( .A1(n13943), .A2(n13418), .B1(n13415), .B2(n15378), .ZN(
        n7853) );
  OAI22_X1 U2174 ( .A1(n13949), .A2(n13417), .B1(n13415), .B2(n15377), .ZN(
        n7854) );
  OAI22_X1 U2175 ( .A1(n13955), .A2(n13417), .B1(n13415), .B2(n15376), .ZN(
        n7855) );
  OAI22_X1 U2176 ( .A1(n13961), .A2(n13417), .B1(n13415), .B2(n15375), .ZN(
        n7856) );
  OAI22_X1 U2177 ( .A1(n13967), .A2(n13417), .B1(n13415), .B2(n15374), .ZN(
        n7857) );
  OAI22_X1 U2178 ( .A1(n13973), .A2(n13417), .B1(n13416), .B2(n15373), .ZN(
        n7858) );
  OAI22_X1 U2179 ( .A1(n13979), .A2(n13417), .B1(n13416), .B2(n15372), .ZN(
        n7859) );
  OAI22_X1 U2180 ( .A1(n13985), .A2(n13417), .B1(n13416), .B2(n15371), .ZN(
        n7860) );
  OAI22_X1 U2181 ( .A1(n13991), .A2(n13417), .B1(n13416), .B2(n15370), .ZN(
        n7861) );
  OAI22_X1 U2182 ( .A1(n13997), .A2(n13417), .B1(n13416), .B2(n15369), .ZN(
        n7862) );
  OAI22_X1 U2183 ( .A1(n14003), .A2(n13417), .B1(n13416), .B2(n15368), .ZN(
        n7863) );
  OAI22_X1 U2184 ( .A1(n14009), .A2(n13417), .B1(n13416), .B2(n15367), .ZN(
        n7864) );
  OAI22_X1 U2185 ( .A1(n14018), .A2(n13417), .B1(n13416), .B2(n15366), .ZN(
        n7865) );
  OAI22_X1 U2186 ( .A1(n13829), .A2(n13425), .B1(n13420), .B2(n15365), .ZN(
        n7866) );
  OAI22_X1 U2187 ( .A1(n13835), .A2(n13425), .B1(n13420), .B2(n15364), .ZN(
        n7867) );
  OAI22_X1 U2188 ( .A1(n13841), .A2(n13425), .B1(n13420), .B2(n15363), .ZN(
        n7868) );
  OAI22_X1 U2189 ( .A1(n13847), .A2(n13425), .B1(n13420), .B2(n15362), .ZN(
        n7869) );
  OAI22_X1 U2190 ( .A1(n13853), .A2(n13425), .B1(n13420), .B2(n15361), .ZN(
        n7870) );
  OAI22_X1 U2191 ( .A1(n13859), .A2(n13425), .B1(n13420), .B2(n15360), .ZN(
        n7871) );
  OAI22_X1 U2192 ( .A1(n13865), .A2(n13425), .B1(n13420), .B2(n15359), .ZN(
        n7872) );
  OAI22_X1 U2193 ( .A1(n13871), .A2(n13425), .B1(n13420), .B2(n15358), .ZN(
        n7873) );
  OAI22_X1 U2194 ( .A1(n13877), .A2(n13424), .B1(n13420), .B2(n15357), .ZN(
        n7874) );
  OAI22_X1 U2195 ( .A1(n13883), .A2(n13424), .B1(n13420), .B2(n15356), .ZN(
        n7875) );
  OAI22_X1 U2196 ( .A1(n13889), .A2(n13424), .B1(n13420), .B2(n15355), .ZN(
        n7876) );
  OAI22_X1 U2197 ( .A1(n13895), .A2(n13424), .B1(n13420), .B2(n15354), .ZN(
        n7877) );
  OAI22_X1 U2198 ( .A1(n13901), .A2(n13424), .B1(n13421), .B2(n15353), .ZN(
        n7878) );
  OAI22_X1 U2199 ( .A1(n13907), .A2(n13424), .B1(n13421), .B2(n15352), .ZN(
        n7879) );
  OAI22_X1 U2200 ( .A1(n13913), .A2(n13424), .B1(n13421), .B2(n15351), .ZN(
        n7880) );
  OAI22_X1 U2201 ( .A1(n13919), .A2(n13424), .B1(n13421), .B2(n15350), .ZN(
        n7881) );
  OAI22_X1 U2202 ( .A1(n13925), .A2(n13424), .B1(n13421), .B2(n15349), .ZN(
        n7882) );
  OAI22_X1 U2203 ( .A1(n13931), .A2(n13424), .B1(n13421), .B2(n15348), .ZN(
        n7883) );
  OAI22_X1 U2204 ( .A1(n13937), .A2(n13424), .B1(n13421), .B2(n15347), .ZN(
        n7884) );
  OAI22_X1 U2205 ( .A1(n13943), .A2(n13424), .B1(n13421), .B2(n15346), .ZN(
        n7885) );
  OAI22_X1 U2206 ( .A1(n13949), .A2(n13423), .B1(n13421), .B2(n15345), .ZN(
        n7886) );
  OAI22_X1 U2207 ( .A1(n13955), .A2(n13423), .B1(n13421), .B2(n15344), .ZN(
        n7887) );
  OAI22_X1 U2208 ( .A1(n13961), .A2(n13423), .B1(n13421), .B2(n15343), .ZN(
        n7888) );
  OAI22_X1 U2209 ( .A1(n13967), .A2(n13423), .B1(n13421), .B2(n15342), .ZN(
        n7889) );
  OAI22_X1 U2210 ( .A1(n13973), .A2(n13423), .B1(n13422), .B2(n15341), .ZN(
        n7890) );
  OAI22_X1 U2211 ( .A1(n13979), .A2(n13423), .B1(n13422), .B2(n15340), .ZN(
        n7891) );
  OAI22_X1 U2212 ( .A1(n13985), .A2(n13423), .B1(n13422), .B2(n15339), .ZN(
        n7892) );
  OAI22_X1 U2213 ( .A1(n13991), .A2(n13423), .B1(n13422), .B2(n15338), .ZN(
        n7893) );
  OAI22_X1 U2214 ( .A1(n13997), .A2(n13423), .B1(n13422), .B2(n15337), .ZN(
        n7894) );
  OAI22_X1 U2215 ( .A1(n14003), .A2(n13423), .B1(n13422), .B2(n15336), .ZN(
        n7895) );
  OAI22_X1 U2216 ( .A1(n14009), .A2(n13423), .B1(n13422), .B2(n15335), .ZN(
        n7896) );
  OAI22_X1 U2217 ( .A1(n14018), .A2(n13423), .B1(n13422), .B2(n15334), .ZN(
        n7897) );
  OAI22_X1 U2218 ( .A1(n13968), .A2(n13393), .B1(n13392), .B2(n15501), .ZN(
        n7730) );
  OAI22_X1 U2219 ( .A1(n13974), .A2(n13393), .B1(n13392), .B2(n15500), .ZN(
        n7731) );
  OAI22_X1 U2220 ( .A1(n13980), .A2(n13393), .B1(n13392), .B2(n15499), .ZN(
        n7732) );
  OAI22_X1 U2221 ( .A1(n13986), .A2(n13393), .B1(n13392), .B2(n15498), .ZN(
        n7733) );
  OAI22_X1 U2222 ( .A1(n13992), .A2(n13393), .B1(n13392), .B2(n15497), .ZN(
        n7734) );
  OAI22_X1 U2223 ( .A1(n13998), .A2(n13393), .B1(n13392), .B2(n15496), .ZN(
        n7735) );
  OAI22_X1 U2224 ( .A1(n14004), .A2(n13393), .B1(n13392), .B2(n15495), .ZN(
        n7736) );
  OAI22_X1 U2225 ( .A1(n14013), .A2(n13393), .B1(n13392), .B2(n15494), .ZN(
        n7737) );
  OAI22_X1 U2226 ( .A1(n13971), .A2(n13525), .B1(n13524), .B2(n15930), .ZN(
        n8434) );
  OAI22_X1 U2227 ( .A1(n13977), .A2(n13525), .B1(n13524), .B2(n15929), .ZN(
        n8435) );
  OAI22_X1 U2228 ( .A1(n13983), .A2(n13525), .B1(n13524), .B2(n15928), .ZN(
        n8436) );
  OAI22_X1 U2229 ( .A1(n13989), .A2(n13525), .B1(n13524), .B2(n15927), .ZN(
        n8437) );
  OAI22_X1 U2230 ( .A1(n13995), .A2(n13525), .B1(n13524), .B2(n15926), .ZN(
        n8438) );
  OAI22_X1 U2231 ( .A1(n14001), .A2(n13525), .B1(n13524), .B2(n15925), .ZN(
        n8439) );
  OAI22_X1 U2232 ( .A1(n14007), .A2(n13525), .B1(n13524), .B2(n15924), .ZN(
        n8440) );
  OAI22_X1 U2233 ( .A1(n14016), .A2(n13525), .B1(n13524), .B2(n15923), .ZN(
        n8441) );
  OAI22_X1 U2234 ( .A1(n13972), .A2(n13441), .B1(n13440), .B2(n15277), .ZN(
        n7986) );
  OAI22_X1 U2235 ( .A1(n13978), .A2(n13441), .B1(n13440), .B2(n15276), .ZN(
        n7987) );
  OAI22_X1 U2236 ( .A1(n13984), .A2(n13441), .B1(n13440), .B2(n15275), .ZN(
        n7988) );
  OAI22_X1 U2237 ( .A1(n13990), .A2(n13441), .B1(n13440), .B2(n15274), .ZN(
        n7989) );
  OAI22_X1 U2238 ( .A1(n13996), .A2(n13441), .B1(n13440), .B2(n15273), .ZN(
        n7990) );
  OAI22_X1 U2239 ( .A1(n14002), .A2(n13441), .B1(n13440), .B2(n15272), .ZN(
        n7991) );
  OAI22_X1 U2240 ( .A1(n14008), .A2(n13441), .B1(n13440), .B2(n15271), .ZN(
        n7992) );
  OAI22_X1 U2241 ( .A1(n14017), .A2(n13441), .B1(n13440), .B2(n15270), .ZN(
        n7993) );
  OAI22_X1 U2242 ( .A1(n13972), .A2(n13447), .B1(n13446), .B2(n15245), .ZN(
        n8018) );
  OAI22_X1 U2243 ( .A1(n13978), .A2(n13447), .B1(n13446), .B2(n15244), .ZN(
        n8019) );
  OAI22_X1 U2244 ( .A1(n13984), .A2(n13447), .B1(n13446), .B2(n15243), .ZN(
        n8020) );
  OAI22_X1 U2245 ( .A1(n13990), .A2(n13447), .B1(n13446), .B2(n15242), .ZN(
        n8021) );
  OAI22_X1 U2246 ( .A1(n13996), .A2(n13447), .B1(n13446), .B2(n15241), .ZN(
        n8022) );
  OAI22_X1 U2247 ( .A1(n14002), .A2(n13447), .B1(n13446), .B2(n15240), .ZN(
        n8023) );
  OAI22_X1 U2248 ( .A1(n14008), .A2(n13447), .B1(n13446), .B2(n15239), .ZN(
        n8024) );
  OAI22_X1 U2249 ( .A1(n14017), .A2(n13447), .B1(n13446), .B2(n15238), .ZN(
        n8025) );
  OAI22_X1 U2250 ( .A1(n13972), .A2(n13453), .B1(n13452), .B2(n15213), .ZN(
        n8050) );
  OAI22_X1 U2251 ( .A1(n13978), .A2(n13453), .B1(n13452), .B2(n15212), .ZN(
        n8051) );
  OAI22_X1 U2252 ( .A1(n13984), .A2(n13453), .B1(n13452), .B2(n15211), .ZN(
        n8052) );
  OAI22_X1 U2253 ( .A1(n13990), .A2(n13453), .B1(n13452), .B2(n15210), .ZN(
        n8053) );
  OAI22_X1 U2254 ( .A1(n13996), .A2(n13453), .B1(n13452), .B2(n15209), .ZN(
        n8054) );
  OAI22_X1 U2255 ( .A1(n14002), .A2(n13453), .B1(n13452), .B2(n15208), .ZN(
        n8055) );
  OAI22_X1 U2256 ( .A1(n14008), .A2(n13453), .B1(n13452), .B2(n15207), .ZN(
        n8056) );
  OAI22_X1 U2257 ( .A1(n14017), .A2(n13453), .B1(n13452), .B2(n15206), .ZN(
        n8057) );
  OAI22_X1 U2258 ( .A1(n13972), .A2(n13483), .B1(n13482), .B2(n15149), .ZN(
        n8210) );
  OAI22_X1 U2259 ( .A1(n13978), .A2(n13483), .B1(n13482), .B2(n15148), .ZN(
        n8211) );
  OAI22_X1 U2260 ( .A1(n13984), .A2(n13483), .B1(n13482), .B2(n15147), .ZN(
        n8212) );
  OAI22_X1 U2261 ( .A1(n13990), .A2(n13483), .B1(n13482), .B2(n15146), .ZN(
        n8213) );
  OAI22_X1 U2262 ( .A1(n13996), .A2(n13483), .B1(n13482), .B2(n15145), .ZN(
        n8214) );
  OAI22_X1 U2263 ( .A1(n14002), .A2(n13483), .B1(n13482), .B2(n15144), .ZN(
        n8215) );
  OAI22_X1 U2264 ( .A1(n14008), .A2(n13483), .B1(n13482), .B2(n15143), .ZN(
        n8216) );
  OAI22_X1 U2265 ( .A1(n14017), .A2(n13483), .B1(n13482), .B2(n15142), .ZN(
        n8217) );
  OAI22_X1 U2266 ( .A1(n13972), .A2(n13489), .B1(n13488), .B2(n15117), .ZN(
        n8242) );
  OAI22_X1 U2267 ( .A1(n13978), .A2(n13489), .B1(n13488), .B2(n15116), .ZN(
        n8243) );
  OAI22_X1 U2268 ( .A1(n13984), .A2(n13489), .B1(n13488), .B2(n15115), .ZN(
        n8244) );
  OAI22_X1 U2269 ( .A1(n13990), .A2(n13489), .B1(n13488), .B2(n15114), .ZN(
        n8245) );
  OAI22_X1 U2270 ( .A1(n13996), .A2(n13489), .B1(n13488), .B2(n15113), .ZN(
        n8246) );
  OAI22_X1 U2271 ( .A1(n14002), .A2(n13489), .B1(n13488), .B2(n15112), .ZN(
        n8247) );
  OAI22_X1 U2272 ( .A1(n14008), .A2(n13489), .B1(n13488), .B2(n15111), .ZN(
        n8248) );
  OAI22_X1 U2273 ( .A1(n14017), .A2(n13489), .B1(n13488), .B2(n15110), .ZN(
        n8249) );
  OAI22_X1 U2274 ( .A1(n13972), .A2(n13495), .B1(n13494), .B2(n15085), .ZN(
        n8274) );
  OAI22_X1 U2275 ( .A1(n13978), .A2(n13495), .B1(n13494), .B2(n15084), .ZN(
        n8275) );
  OAI22_X1 U2276 ( .A1(n13984), .A2(n13495), .B1(n13494), .B2(n15083), .ZN(
        n8276) );
  OAI22_X1 U2277 ( .A1(n13990), .A2(n13495), .B1(n13494), .B2(n15082), .ZN(
        n8277) );
  OAI22_X1 U2278 ( .A1(n13996), .A2(n13495), .B1(n13494), .B2(n15081), .ZN(
        n8278) );
  OAI22_X1 U2279 ( .A1(n14002), .A2(n13495), .B1(n13494), .B2(n15080), .ZN(
        n8279) );
  OAI22_X1 U2280 ( .A1(n14008), .A2(n13495), .B1(n13494), .B2(n15079), .ZN(
        n8280) );
  OAI22_X1 U2281 ( .A1(n14017), .A2(n13495), .B1(n13494), .B2(n15078), .ZN(
        n8281) );
  OAI22_X1 U2282 ( .A1(n13972), .A2(n13501), .B1(n13500), .B2(n15053), .ZN(
        n8306) );
  OAI22_X1 U2283 ( .A1(n13978), .A2(n13501), .B1(n13500), .B2(n15052), .ZN(
        n8307) );
  OAI22_X1 U2284 ( .A1(n13984), .A2(n13501), .B1(n13500), .B2(n15051), .ZN(
        n8308) );
  OAI22_X1 U2285 ( .A1(n13990), .A2(n13501), .B1(n13500), .B2(n15050), .ZN(
        n8309) );
  OAI22_X1 U2286 ( .A1(n13996), .A2(n13501), .B1(n13500), .B2(n15049), .ZN(
        n8310) );
  OAI22_X1 U2287 ( .A1(n14002), .A2(n13501), .B1(n13500), .B2(n15048), .ZN(
        n8311) );
  OAI22_X1 U2288 ( .A1(n14008), .A2(n13501), .B1(n13500), .B2(n15047), .ZN(
        n8312) );
  OAI22_X1 U2289 ( .A1(n14017), .A2(n13501), .B1(n13500), .B2(n15046), .ZN(
        n8313) );
  OAI22_X1 U2290 ( .A1(n13972), .A2(n13507), .B1(n13506), .B2(n15021), .ZN(
        n8338) );
  OAI22_X1 U2291 ( .A1(n13978), .A2(n13507), .B1(n13506), .B2(n15020), .ZN(
        n8339) );
  OAI22_X1 U2292 ( .A1(n13984), .A2(n13507), .B1(n13506), .B2(n15019), .ZN(
        n8340) );
  OAI22_X1 U2293 ( .A1(n13990), .A2(n13507), .B1(n13506), .B2(n15018), .ZN(
        n8341) );
  OAI22_X1 U2294 ( .A1(n13996), .A2(n13507), .B1(n13506), .B2(n15017), .ZN(
        n8342) );
  OAI22_X1 U2295 ( .A1(n14002), .A2(n13507), .B1(n13506), .B2(n15016), .ZN(
        n8343) );
  OAI22_X1 U2296 ( .A1(n14008), .A2(n13507), .B1(n13506), .B2(n15015), .ZN(
        n8344) );
  OAI22_X1 U2297 ( .A1(n14017), .A2(n13507), .B1(n13506), .B2(n15014), .ZN(
        n8345) );
  OAI22_X1 U2298 ( .A1(n13971), .A2(n13531), .B1(n13530), .B2(n14956), .ZN(
        n8466) );
  OAI22_X1 U2299 ( .A1(n13977), .A2(n13531), .B1(n13530), .B2(n14955), .ZN(
        n8467) );
  OAI22_X1 U2300 ( .A1(n13983), .A2(n13531), .B1(n13530), .B2(n14954), .ZN(
        n8468) );
  OAI22_X1 U2301 ( .A1(n13989), .A2(n13531), .B1(n13530), .B2(n14953), .ZN(
        n8469) );
  OAI22_X1 U2302 ( .A1(n13995), .A2(n13531), .B1(n13530), .B2(n14952), .ZN(
        n8470) );
  OAI22_X1 U2303 ( .A1(n14001), .A2(n13531), .B1(n13530), .B2(n14951), .ZN(
        n8471) );
  OAI22_X1 U2304 ( .A1(n14007), .A2(n13531), .B1(n13530), .B2(n14950), .ZN(
        n8472) );
  OAI22_X1 U2305 ( .A1(n14016), .A2(n13531), .B1(n13530), .B2(n14949), .ZN(
        n8473) );
  OAI22_X1 U2306 ( .A1(n13971), .A2(n13549), .B1(n13548), .B2(n14923), .ZN(
        n8562) );
  OAI22_X1 U2307 ( .A1(n13977), .A2(n13549), .B1(n13548), .B2(n14922), .ZN(
        n8563) );
  OAI22_X1 U2308 ( .A1(n13983), .A2(n13549), .B1(n13548), .B2(n14921), .ZN(
        n8564) );
  OAI22_X1 U2309 ( .A1(n13989), .A2(n13549), .B1(n13548), .B2(n14920), .ZN(
        n8565) );
  OAI22_X1 U2310 ( .A1(n13995), .A2(n13549), .B1(n13548), .B2(n14919), .ZN(
        n8566) );
  OAI22_X1 U2311 ( .A1(n14001), .A2(n13549), .B1(n13548), .B2(n14918), .ZN(
        n8567) );
  OAI22_X1 U2312 ( .A1(n14007), .A2(n13549), .B1(n13548), .B2(n14917), .ZN(
        n8568) );
  OAI22_X1 U2313 ( .A1(n14016), .A2(n13549), .B1(n13548), .B2(n14916), .ZN(
        n8569) );
  OAI22_X1 U2314 ( .A1(n13971), .A2(n13555), .B1(n13554), .B2(n14891), .ZN(
        n8594) );
  OAI22_X1 U2315 ( .A1(n13977), .A2(n13555), .B1(n13554), .B2(n14890), .ZN(
        n8595) );
  OAI22_X1 U2316 ( .A1(n13983), .A2(n13555), .B1(n13554), .B2(n14889), .ZN(
        n8596) );
  OAI22_X1 U2317 ( .A1(n13989), .A2(n13555), .B1(n13554), .B2(n14888), .ZN(
        n8597) );
  OAI22_X1 U2318 ( .A1(n13995), .A2(n13555), .B1(n13554), .B2(n14887), .ZN(
        n8598) );
  OAI22_X1 U2319 ( .A1(n14001), .A2(n13555), .B1(n13554), .B2(n14886), .ZN(
        n8599) );
  OAI22_X1 U2320 ( .A1(n14007), .A2(n13555), .B1(n13554), .B2(n14885), .ZN(
        n8600) );
  OAI22_X1 U2321 ( .A1(n14016), .A2(n13555), .B1(n13554), .B2(n14884), .ZN(
        n8601) );
  OAI22_X1 U2322 ( .A1(n13971), .A2(n13561), .B1(n13560), .B2(n14859), .ZN(
        n8626) );
  OAI22_X1 U2323 ( .A1(n13977), .A2(n13561), .B1(n13560), .B2(n14858), .ZN(
        n8627) );
  OAI22_X1 U2324 ( .A1(n13983), .A2(n13561), .B1(n13560), .B2(n14857), .ZN(
        n8628) );
  OAI22_X1 U2325 ( .A1(n13989), .A2(n13561), .B1(n13560), .B2(n14856), .ZN(
        n8629) );
  OAI22_X1 U2326 ( .A1(n13995), .A2(n13561), .B1(n13560), .B2(n14855), .ZN(
        n8630) );
  OAI22_X1 U2327 ( .A1(n14001), .A2(n13561), .B1(n13560), .B2(n14854), .ZN(
        n8631) );
  OAI22_X1 U2328 ( .A1(n14007), .A2(n13561), .B1(n13560), .B2(n14853), .ZN(
        n8632) );
  OAI22_X1 U2329 ( .A1(n14016), .A2(n13561), .B1(n13560), .B2(n14852), .ZN(
        n8633) );
  OAI22_X1 U2330 ( .A1(n13971), .A2(n13591), .B1(n13590), .B2(n14827), .ZN(
        n8786) );
  OAI22_X1 U2331 ( .A1(n13977), .A2(n13591), .B1(n13590), .B2(n14826), .ZN(
        n8787) );
  OAI22_X1 U2332 ( .A1(n13983), .A2(n13591), .B1(n13590), .B2(n14825), .ZN(
        n8788) );
  OAI22_X1 U2333 ( .A1(n13989), .A2(n13591), .B1(n13590), .B2(n14824), .ZN(
        n8789) );
  OAI22_X1 U2334 ( .A1(n13995), .A2(n13591), .B1(n13590), .B2(n14823), .ZN(
        n8790) );
  OAI22_X1 U2335 ( .A1(n14001), .A2(n13591), .B1(n13590), .B2(n14822), .ZN(
        n8791) );
  OAI22_X1 U2336 ( .A1(n14007), .A2(n13591), .B1(n13590), .B2(n14821), .ZN(
        n8792) );
  OAI22_X1 U2337 ( .A1(n14016), .A2(n13591), .B1(n13590), .B2(n14820), .ZN(
        n8793) );
  OAI22_X1 U2338 ( .A1(n13970), .A2(n13597), .B1(n13596), .B2(n14795), .ZN(
        n8818) );
  OAI22_X1 U2339 ( .A1(n13976), .A2(n13597), .B1(n13596), .B2(n14794), .ZN(
        n8819) );
  OAI22_X1 U2340 ( .A1(n13982), .A2(n13597), .B1(n13596), .B2(n14793), .ZN(
        n8820) );
  OAI22_X1 U2341 ( .A1(n13988), .A2(n13597), .B1(n13596), .B2(n14792), .ZN(
        n8821) );
  OAI22_X1 U2342 ( .A1(n13994), .A2(n13597), .B1(n13596), .B2(n14791), .ZN(
        n8822) );
  OAI22_X1 U2343 ( .A1(n14000), .A2(n13597), .B1(n13596), .B2(n14790), .ZN(
        n8823) );
  OAI22_X1 U2344 ( .A1(n14006), .A2(n13597), .B1(n13596), .B2(n14789), .ZN(
        n8824) );
  OAI22_X1 U2345 ( .A1(n14015), .A2(n13597), .B1(n13596), .B2(n14788), .ZN(
        n8825) );
  OAI22_X1 U2346 ( .A1(n13970), .A2(n13603), .B1(n13602), .B2(n14763), .ZN(
        n8850) );
  OAI22_X1 U2347 ( .A1(n13976), .A2(n13603), .B1(n13602), .B2(n14762), .ZN(
        n8851) );
  OAI22_X1 U2348 ( .A1(n13982), .A2(n13603), .B1(n13602), .B2(n14761), .ZN(
        n8852) );
  OAI22_X1 U2349 ( .A1(n13988), .A2(n13603), .B1(n13602), .B2(n14760), .ZN(
        n8853) );
  OAI22_X1 U2350 ( .A1(n13994), .A2(n13603), .B1(n13602), .B2(n14759), .ZN(
        n8854) );
  OAI22_X1 U2351 ( .A1(n14000), .A2(n13603), .B1(n13602), .B2(n14758), .ZN(
        n8855) );
  OAI22_X1 U2352 ( .A1(n14006), .A2(n13603), .B1(n13602), .B2(n14757), .ZN(
        n8856) );
  OAI22_X1 U2353 ( .A1(n14015), .A2(n13603), .B1(n13602), .B2(n14756), .ZN(
        n8857) );
  OAI22_X1 U2354 ( .A1(n13970), .A2(n13609), .B1(n13608), .B2(n14731), .ZN(
        n8882) );
  OAI22_X1 U2355 ( .A1(n13976), .A2(n13609), .B1(n13608), .B2(n14730), .ZN(
        n8883) );
  OAI22_X1 U2356 ( .A1(n13982), .A2(n13609), .B1(n13608), .B2(n14729), .ZN(
        n8884) );
  OAI22_X1 U2357 ( .A1(n13988), .A2(n13609), .B1(n13608), .B2(n14728), .ZN(
        n8885) );
  OAI22_X1 U2358 ( .A1(n13994), .A2(n13609), .B1(n13608), .B2(n14727), .ZN(
        n8886) );
  OAI22_X1 U2359 ( .A1(n14000), .A2(n13609), .B1(n13608), .B2(n14726), .ZN(
        n8887) );
  OAI22_X1 U2360 ( .A1(n14006), .A2(n13609), .B1(n13608), .B2(n14725), .ZN(
        n8888) );
  OAI22_X1 U2361 ( .A1(n14015), .A2(n13609), .B1(n13608), .B2(n14724), .ZN(
        n8889) );
  OAI22_X1 U2362 ( .A1(n13970), .A2(n13615), .B1(n13614), .B2(n14699), .ZN(
        n8914) );
  OAI22_X1 U2363 ( .A1(n13976), .A2(n13615), .B1(n13614), .B2(n14698), .ZN(
        n8915) );
  OAI22_X1 U2364 ( .A1(n13982), .A2(n13615), .B1(n13614), .B2(n14697), .ZN(
        n8916) );
  OAI22_X1 U2365 ( .A1(n13988), .A2(n13615), .B1(n13614), .B2(n14696), .ZN(
        n8917) );
  OAI22_X1 U2366 ( .A1(n13994), .A2(n13615), .B1(n13614), .B2(n14695), .ZN(
        n8918) );
  OAI22_X1 U2367 ( .A1(n14000), .A2(n13615), .B1(n13614), .B2(n14694), .ZN(
        n8919) );
  OAI22_X1 U2368 ( .A1(n14006), .A2(n13615), .B1(n13614), .B2(n14693), .ZN(
        n8920) );
  OAI22_X1 U2369 ( .A1(n14015), .A2(n13615), .B1(n13614), .B2(n14692), .ZN(
        n8921) );
  OAI22_X1 U2370 ( .A1(n13970), .A2(n13645), .B1(n13644), .B2(n14628), .ZN(
        n9074) );
  OAI22_X1 U2371 ( .A1(n13976), .A2(n13645), .B1(n13644), .B2(n14627), .ZN(
        n9075) );
  OAI22_X1 U2372 ( .A1(n13982), .A2(n13645), .B1(n13644), .B2(n14626), .ZN(
        n9076) );
  OAI22_X1 U2373 ( .A1(n13988), .A2(n13645), .B1(n13644), .B2(n14625), .ZN(
        n9077) );
  OAI22_X1 U2374 ( .A1(n13994), .A2(n13645), .B1(n13644), .B2(n14624), .ZN(
        n9078) );
  OAI22_X1 U2375 ( .A1(n14000), .A2(n13645), .B1(n13644), .B2(n14623), .ZN(
        n9079) );
  OAI22_X1 U2376 ( .A1(n14006), .A2(n13645), .B1(n13644), .B2(n14622), .ZN(
        n9080) );
  OAI22_X1 U2377 ( .A1(n14015), .A2(n13645), .B1(n13644), .B2(n14621), .ZN(
        n9081) );
  OAI22_X1 U2378 ( .A1(n13970), .A2(n13651), .B1(n13650), .B2(n14596), .ZN(
        n9106) );
  OAI22_X1 U2379 ( .A1(n13976), .A2(n13651), .B1(n13650), .B2(n14595), .ZN(
        n9107) );
  OAI22_X1 U2380 ( .A1(n13982), .A2(n13651), .B1(n13650), .B2(n14594), .ZN(
        n9108) );
  OAI22_X1 U2381 ( .A1(n13988), .A2(n13651), .B1(n13650), .B2(n14593), .ZN(
        n9109) );
  OAI22_X1 U2382 ( .A1(n13994), .A2(n13651), .B1(n13650), .B2(n14592), .ZN(
        n9110) );
  OAI22_X1 U2383 ( .A1(n14000), .A2(n13651), .B1(n13650), .B2(n14591), .ZN(
        n9111) );
  OAI22_X1 U2384 ( .A1(n14006), .A2(n13651), .B1(n13650), .B2(n14590), .ZN(
        n9112) );
  OAI22_X1 U2385 ( .A1(n14015), .A2(n13651), .B1(n13650), .B2(n14589), .ZN(
        n9113) );
  OAI22_X1 U2386 ( .A1(n13970), .A2(n13657), .B1(n13656), .B2(n14564), .ZN(
        n9138) );
  OAI22_X1 U2387 ( .A1(n13976), .A2(n13657), .B1(n13656), .B2(n14563), .ZN(
        n9139) );
  OAI22_X1 U2388 ( .A1(n13982), .A2(n13657), .B1(n13656), .B2(n14562), .ZN(
        n9140) );
  OAI22_X1 U2389 ( .A1(n13988), .A2(n13657), .B1(n13656), .B2(n14561), .ZN(
        n9141) );
  OAI22_X1 U2390 ( .A1(n13994), .A2(n13657), .B1(n13656), .B2(n14560), .ZN(
        n9142) );
  OAI22_X1 U2391 ( .A1(n14000), .A2(n13657), .B1(n13656), .B2(n14559), .ZN(
        n9143) );
  OAI22_X1 U2392 ( .A1(n14006), .A2(n13657), .B1(n13656), .B2(n14558), .ZN(
        n9144) );
  OAI22_X1 U2393 ( .A1(n14015), .A2(n13657), .B1(n13656), .B2(n14557), .ZN(
        n9145) );
  OAI22_X1 U2394 ( .A1(n13970), .A2(n13663), .B1(n13662), .B2(n14532), .ZN(
        n9170) );
  OAI22_X1 U2395 ( .A1(n13976), .A2(n13663), .B1(n13662), .B2(n14531), .ZN(
        n9171) );
  OAI22_X1 U2396 ( .A1(n13982), .A2(n13663), .B1(n13662), .B2(n14530), .ZN(
        n9172) );
  OAI22_X1 U2397 ( .A1(n13988), .A2(n13663), .B1(n13662), .B2(n14529), .ZN(
        n9173) );
  OAI22_X1 U2398 ( .A1(n13994), .A2(n13663), .B1(n13662), .B2(n14528), .ZN(
        n9174) );
  OAI22_X1 U2399 ( .A1(n14000), .A2(n13663), .B1(n13662), .B2(n14527), .ZN(
        n9175) );
  OAI22_X1 U2400 ( .A1(n14006), .A2(n13663), .B1(n13662), .B2(n14526), .ZN(
        n9176) );
  OAI22_X1 U2401 ( .A1(n14015), .A2(n13663), .B1(n13662), .B2(n14525), .ZN(
        n9177) );
  OAI22_X1 U2402 ( .A1(n13969), .A2(n13669), .B1(n13668), .B2(n14500), .ZN(
        n9202) );
  OAI22_X1 U2403 ( .A1(n13975), .A2(n13669), .B1(n13668), .B2(n14499), .ZN(
        n9203) );
  OAI22_X1 U2404 ( .A1(n13981), .A2(n13669), .B1(n13668), .B2(n14498), .ZN(
        n9204) );
  OAI22_X1 U2405 ( .A1(n13987), .A2(n13669), .B1(n13668), .B2(n14497), .ZN(
        n9205) );
  OAI22_X1 U2406 ( .A1(n13993), .A2(n13669), .B1(n13668), .B2(n14496), .ZN(
        n9206) );
  OAI22_X1 U2407 ( .A1(n13999), .A2(n13669), .B1(n13668), .B2(n14495), .ZN(
        n9207) );
  OAI22_X1 U2408 ( .A1(n14005), .A2(n13669), .B1(n13668), .B2(n14494), .ZN(
        n9208) );
  OAI22_X1 U2409 ( .A1(n14014), .A2(n13669), .B1(n13668), .B2(n14493), .ZN(
        n9209) );
  OAI22_X1 U2410 ( .A1(n13969), .A2(n13699), .B1(n13698), .B2(n14415), .ZN(
        n9362) );
  OAI22_X1 U2411 ( .A1(n13975), .A2(n13699), .B1(n13698), .B2(n14414), .ZN(
        n9363) );
  OAI22_X1 U2412 ( .A1(n13981), .A2(n13699), .B1(n13698), .B2(n14413), .ZN(
        n9364) );
  OAI22_X1 U2413 ( .A1(n13987), .A2(n13699), .B1(n13698), .B2(n14412), .ZN(
        n9365) );
  OAI22_X1 U2414 ( .A1(n13993), .A2(n13699), .B1(n13698), .B2(n14411), .ZN(
        n9366) );
  OAI22_X1 U2415 ( .A1(n13999), .A2(n13699), .B1(n13698), .B2(n14410), .ZN(
        n9367) );
  OAI22_X1 U2416 ( .A1(n14005), .A2(n13699), .B1(n13698), .B2(n14409), .ZN(
        n9368) );
  OAI22_X1 U2417 ( .A1(n14014), .A2(n13699), .B1(n13698), .B2(n14408), .ZN(
        n9369) );
  OAI22_X1 U2418 ( .A1(n13970), .A2(n13705), .B1(n13704), .B2(n14383), .ZN(
        n9394) );
  OAI22_X1 U2419 ( .A1(n13976), .A2(n13705), .B1(n13704), .B2(n14382), .ZN(
        n9395) );
  OAI22_X1 U2420 ( .A1(n13982), .A2(n13705), .B1(n13704), .B2(n14381), .ZN(
        n9396) );
  OAI22_X1 U2421 ( .A1(n13988), .A2(n13705), .B1(n13704), .B2(n14380), .ZN(
        n9397) );
  OAI22_X1 U2422 ( .A1(n13994), .A2(n13705), .B1(n13704), .B2(n14379), .ZN(
        n9398) );
  OAI22_X1 U2423 ( .A1(n14000), .A2(n13705), .B1(n13704), .B2(n14378), .ZN(
        n9399) );
  OAI22_X1 U2424 ( .A1(n14006), .A2(n13705), .B1(n13704), .B2(n14377), .ZN(
        n9400) );
  OAI22_X1 U2425 ( .A1(n14015), .A2(n13705), .B1(n13704), .B2(n14376), .ZN(
        n9401) );
  OAI22_X1 U2426 ( .A1(n13969), .A2(n13711), .B1(n13710), .B2(n14351), .ZN(
        n9426) );
  OAI22_X1 U2427 ( .A1(n13975), .A2(n13711), .B1(n13710), .B2(n14350), .ZN(
        n9427) );
  OAI22_X1 U2428 ( .A1(n13981), .A2(n13711), .B1(n13710), .B2(n14349), .ZN(
        n9428) );
  OAI22_X1 U2429 ( .A1(n13987), .A2(n13711), .B1(n13710), .B2(n14348), .ZN(
        n9429) );
  OAI22_X1 U2430 ( .A1(n13993), .A2(n13711), .B1(n13710), .B2(n14347), .ZN(
        n9430) );
  OAI22_X1 U2431 ( .A1(n13999), .A2(n13711), .B1(n13710), .B2(n14346), .ZN(
        n9431) );
  OAI22_X1 U2432 ( .A1(n14005), .A2(n13711), .B1(n13710), .B2(n14345), .ZN(
        n9432) );
  OAI22_X1 U2433 ( .A1(n14014), .A2(n13711), .B1(n13710), .B2(n14344), .ZN(
        n9433) );
  OAI22_X1 U2434 ( .A1(n13969), .A2(n13717), .B1(n13716), .B2(n14319), .ZN(
        n9458) );
  OAI22_X1 U2435 ( .A1(n13975), .A2(n13717), .B1(n13716), .B2(n14318), .ZN(
        n9459) );
  OAI22_X1 U2436 ( .A1(n13981), .A2(n13717), .B1(n13716), .B2(n14317), .ZN(
        n9460) );
  OAI22_X1 U2437 ( .A1(n13987), .A2(n13717), .B1(n13716), .B2(n14316), .ZN(
        n9461) );
  OAI22_X1 U2438 ( .A1(n13993), .A2(n13717), .B1(n13716), .B2(n14315), .ZN(
        n9462) );
  OAI22_X1 U2439 ( .A1(n13999), .A2(n13717), .B1(n13716), .B2(n14314), .ZN(
        n9463) );
  OAI22_X1 U2440 ( .A1(n14005), .A2(n13717), .B1(n13716), .B2(n14313), .ZN(
        n9464) );
  OAI22_X1 U2441 ( .A1(n14014), .A2(n13717), .B1(n13716), .B2(n14312), .ZN(
        n9465) );
  OAI22_X1 U2442 ( .A1(n13969), .A2(n13723), .B1(n13722), .B2(n14287), .ZN(
        n9490) );
  OAI22_X1 U2443 ( .A1(n13975), .A2(n13723), .B1(n13722), .B2(n14286), .ZN(
        n9491) );
  OAI22_X1 U2444 ( .A1(n13981), .A2(n13723), .B1(n13722), .B2(n14285), .ZN(
        n9492) );
  OAI22_X1 U2445 ( .A1(n13987), .A2(n13723), .B1(n13722), .B2(n14284), .ZN(
        n9493) );
  OAI22_X1 U2446 ( .A1(n13993), .A2(n13723), .B1(n13722), .B2(n14283), .ZN(
        n9494) );
  OAI22_X1 U2447 ( .A1(n13999), .A2(n13723), .B1(n13722), .B2(n14282), .ZN(
        n9495) );
  OAI22_X1 U2448 ( .A1(n14005), .A2(n13723), .B1(n13722), .B2(n14281), .ZN(
        n9496) );
  OAI22_X1 U2449 ( .A1(n14014), .A2(n13723), .B1(n13722), .B2(n14280), .ZN(
        n9497) );
  OAI22_X1 U2450 ( .A1(n13968), .A2(n13747), .B1(n13746), .B2(n12657), .ZN(
        n9618) );
  OAI22_X1 U2451 ( .A1(n13974), .A2(n13747), .B1(n13746), .B2(n12658), .ZN(
        n9619) );
  OAI22_X1 U2452 ( .A1(n13980), .A2(n13747), .B1(n13746), .B2(n12659), .ZN(
        n9620) );
  OAI22_X1 U2453 ( .A1(n13986), .A2(n13747), .B1(n13746), .B2(n12660), .ZN(
        n9621) );
  OAI22_X1 U2454 ( .A1(n13992), .A2(n13747), .B1(n13746), .B2(n12653), .ZN(
        n9622) );
  OAI22_X1 U2455 ( .A1(n13998), .A2(n13747), .B1(n13746), .B2(n12654), .ZN(
        n9623) );
  OAI22_X1 U2456 ( .A1(n14004), .A2(n13747), .B1(n13746), .B2(n12655), .ZN(
        n9624) );
  OAI22_X1 U2457 ( .A1(n14013), .A2(n13747), .B1(n13746), .B2(n12656), .ZN(
        n9625) );
  OAI22_X1 U2458 ( .A1(n13968), .A2(n13765), .B1(n13764), .B2(n14179), .ZN(
        n9714) );
  OAI22_X1 U2459 ( .A1(n13974), .A2(n13765), .B1(n13764), .B2(n14178), .ZN(
        n9715) );
  OAI22_X1 U2460 ( .A1(n13980), .A2(n13765), .B1(n13764), .B2(n14177), .ZN(
        n9716) );
  OAI22_X1 U2461 ( .A1(n13986), .A2(n13765), .B1(n13764), .B2(n14176), .ZN(
        n9717) );
  OAI22_X1 U2462 ( .A1(n13992), .A2(n13765), .B1(n13764), .B2(n14175), .ZN(
        n9718) );
  OAI22_X1 U2463 ( .A1(n13998), .A2(n13765), .B1(n13764), .B2(n14174), .ZN(
        n9719) );
  OAI22_X1 U2464 ( .A1(n14004), .A2(n13765), .B1(n13764), .B2(n14173), .ZN(
        n9720) );
  OAI22_X1 U2465 ( .A1(n14013), .A2(n13765), .B1(n13764), .B2(n14172), .ZN(
        n9721) );
  OAI22_X1 U2466 ( .A1(n13968), .A2(n13771), .B1(n13770), .B2(n14147), .ZN(
        n9746) );
  OAI22_X1 U2467 ( .A1(n13974), .A2(n13771), .B1(n13770), .B2(n14146), .ZN(
        n9747) );
  OAI22_X1 U2468 ( .A1(n13980), .A2(n13771), .B1(n13770), .B2(n14145), .ZN(
        n9748) );
  OAI22_X1 U2469 ( .A1(n13986), .A2(n13771), .B1(n13770), .B2(n14144), .ZN(
        n9749) );
  OAI22_X1 U2470 ( .A1(n13992), .A2(n13771), .B1(n13770), .B2(n14143), .ZN(
        n9750) );
  OAI22_X1 U2471 ( .A1(n13998), .A2(n13771), .B1(n13770), .B2(n14142), .ZN(
        n9751) );
  OAI22_X1 U2472 ( .A1(n14004), .A2(n13771), .B1(n13770), .B2(n14141), .ZN(
        n9752) );
  OAI22_X1 U2473 ( .A1(n14013), .A2(n13771), .B1(n13770), .B2(n14140), .ZN(
        n9753) );
  OAI22_X1 U2474 ( .A1(n13968), .A2(n13777), .B1(n13776), .B2(n14115), .ZN(
        n9778) );
  OAI22_X1 U2475 ( .A1(n13974), .A2(n13777), .B1(n13776), .B2(n14114), .ZN(
        n9779) );
  OAI22_X1 U2476 ( .A1(n13980), .A2(n13777), .B1(n13776), .B2(n14113), .ZN(
        n9780) );
  OAI22_X1 U2477 ( .A1(n13986), .A2(n13777), .B1(n13776), .B2(n14112), .ZN(
        n9781) );
  OAI22_X1 U2478 ( .A1(n13992), .A2(n13777), .B1(n13776), .B2(n14111), .ZN(
        n9782) );
  OAI22_X1 U2479 ( .A1(n13998), .A2(n13777), .B1(n13776), .B2(n14110), .ZN(
        n9783) );
  OAI22_X1 U2480 ( .A1(n14004), .A2(n13777), .B1(n13776), .B2(n14109), .ZN(
        n9784) );
  OAI22_X1 U2481 ( .A1(n14013), .A2(n13777), .B1(n13776), .B2(n14108), .ZN(
        n9785) );
  OAI22_X1 U2482 ( .A1(n13968), .A2(n13801), .B1(n13800), .B2(n12649), .ZN(
        n9906) );
  OAI22_X1 U2483 ( .A1(n13974), .A2(n13801), .B1(n13800), .B2(n12650), .ZN(
        n9907) );
  OAI22_X1 U2484 ( .A1(n13980), .A2(n13801), .B1(n13800), .B2(n12651), .ZN(
        n9908) );
  OAI22_X1 U2485 ( .A1(n13986), .A2(n13801), .B1(n13800), .B2(n12652), .ZN(
        n9909) );
  OAI22_X1 U2486 ( .A1(n13992), .A2(n13801), .B1(n13800), .B2(n12645), .ZN(
        n9910) );
  OAI22_X1 U2487 ( .A1(n13998), .A2(n13801), .B1(n13800), .B2(n12646), .ZN(
        n9911) );
  OAI22_X1 U2488 ( .A1(n14004), .A2(n13801), .B1(n13800), .B2(n12647), .ZN(
        n9912) );
  OAI22_X1 U2489 ( .A1(n14013), .A2(n13801), .B1(n13800), .B2(n12648), .ZN(
        n9913) );
  OAI22_X1 U2490 ( .A1(n13387), .A2(n15556), .B1(n13830), .B2(n13386), .ZN(
        n7675) );
  OAI22_X1 U2491 ( .A1(n13387), .A2(n15555), .B1(n13836), .B2(n13386), .ZN(
        n7676) );
  OAI22_X1 U2492 ( .A1(n13387), .A2(n15554), .B1(n13842), .B2(n13386), .ZN(
        n7677) );
  OAI22_X1 U2493 ( .A1(n13387), .A2(n15553), .B1(n13848), .B2(n13386), .ZN(
        n7678) );
  OAI22_X1 U2494 ( .A1(n13387), .A2(n15552), .B1(n13854), .B2(n13386), .ZN(
        n7679) );
  OAI22_X1 U2495 ( .A1(n13387), .A2(n15551), .B1(n13860), .B2(n13386), .ZN(
        n7680) );
  OAI22_X1 U2496 ( .A1(n13387), .A2(n15550), .B1(n13866), .B2(n13386), .ZN(
        n7681) );
  OAI22_X1 U2497 ( .A1(n13387), .A2(n15549), .B1(n13872), .B2(n13386), .ZN(
        n7682) );
  OAI22_X1 U2498 ( .A1(n13827), .A2(n13527), .B1(n13522), .B2(n15970), .ZN(
        n8410) );
  OAI22_X1 U2499 ( .A1(n13833), .A2(n13527), .B1(n13522), .B2(n15969), .ZN(
        n8411) );
  OAI22_X1 U2500 ( .A1(n13839), .A2(n13527), .B1(n13522), .B2(n15968), .ZN(
        n8412) );
  OAI22_X1 U2501 ( .A1(n13845), .A2(n13527), .B1(n13522), .B2(n15967), .ZN(
        n8413) );
  OAI22_X1 U2502 ( .A1(n13851), .A2(n13527), .B1(n13522), .B2(n15966), .ZN(
        n8414) );
  OAI22_X1 U2503 ( .A1(n13857), .A2(n13527), .B1(n13522), .B2(n15965), .ZN(
        n8415) );
  OAI22_X1 U2504 ( .A1(n13863), .A2(n13527), .B1(n13522), .B2(n15964), .ZN(
        n8416) );
  OAI22_X1 U2505 ( .A1(n13869), .A2(n13527), .B1(n13522), .B2(n15963), .ZN(
        n8417) );
  OAI22_X1 U2506 ( .A1(n13875), .A2(n13526), .B1(n13522), .B2(n15962), .ZN(
        n8418) );
  OAI22_X1 U2507 ( .A1(n13881), .A2(n13526), .B1(n13522), .B2(n15961), .ZN(
        n8419) );
  OAI22_X1 U2508 ( .A1(n13887), .A2(n13526), .B1(n13522), .B2(n15960), .ZN(
        n8420) );
  OAI22_X1 U2509 ( .A1(n13893), .A2(n13526), .B1(n13522), .B2(n15959), .ZN(
        n8421) );
  OAI22_X1 U2510 ( .A1(n13899), .A2(n13526), .B1(n13523), .B2(n15958), .ZN(
        n8422) );
  OAI22_X1 U2511 ( .A1(n13905), .A2(n13526), .B1(n13523), .B2(n15957), .ZN(
        n8423) );
  OAI22_X1 U2512 ( .A1(n13911), .A2(n13526), .B1(n13523), .B2(n15956), .ZN(
        n8424) );
  OAI22_X1 U2513 ( .A1(n13917), .A2(n13526), .B1(n13523), .B2(n15955), .ZN(
        n8425) );
  OAI22_X1 U2514 ( .A1(n13923), .A2(n13526), .B1(n13523), .B2(n15954), .ZN(
        n8426) );
  OAI22_X1 U2515 ( .A1(n13929), .A2(n13526), .B1(n13523), .B2(n15953), .ZN(
        n8427) );
  OAI22_X1 U2516 ( .A1(n13935), .A2(n13526), .B1(n13523), .B2(n15952), .ZN(
        n8428) );
  OAI22_X1 U2517 ( .A1(n13941), .A2(n13526), .B1(n13523), .B2(n15951), .ZN(
        n8429) );
  OAI22_X1 U2518 ( .A1(n13947), .A2(n13525), .B1(n13523), .B2(n15950), .ZN(
        n8430) );
  OAI22_X1 U2519 ( .A1(n13953), .A2(n13525), .B1(n13523), .B2(n15949), .ZN(
        n8431) );
  OAI22_X1 U2520 ( .A1(n13959), .A2(n13525), .B1(n13523), .B2(n15948), .ZN(
        n8432) );
  OAI22_X1 U2521 ( .A1(n13965), .A2(n13525), .B1(n13523), .B2(n15947), .ZN(
        n8433) );
  OAI22_X1 U2522 ( .A1(n13830), .A2(n13395), .B1(n13390), .B2(n15524), .ZN(
        n7707) );
  OAI22_X1 U2523 ( .A1(n13836), .A2(n13395), .B1(n13390), .B2(n15523), .ZN(
        n7708) );
  OAI22_X1 U2524 ( .A1(n13842), .A2(n13395), .B1(n13390), .B2(n15522), .ZN(
        n7709) );
  OAI22_X1 U2525 ( .A1(n13848), .A2(n13395), .B1(n13390), .B2(n15521), .ZN(
        n7710) );
  OAI22_X1 U2526 ( .A1(n13854), .A2(n13395), .B1(n13390), .B2(n15520), .ZN(
        n7711) );
  OAI22_X1 U2527 ( .A1(n13860), .A2(n13395), .B1(n13390), .B2(n15519), .ZN(
        n7712) );
  OAI22_X1 U2528 ( .A1(n13866), .A2(n13395), .B1(n13390), .B2(n15518), .ZN(
        n7713) );
  OAI22_X1 U2529 ( .A1(n13872), .A2(n13394), .B1(n13390), .B2(n15517), .ZN(
        n7714) );
  OAI22_X1 U2530 ( .A1(n13878), .A2(n13394), .B1(n13390), .B2(n15516), .ZN(
        n7715) );
  OAI22_X1 U2531 ( .A1(n13884), .A2(n13394), .B1(n13390), .B2(n15515), .ZN(
        n7716) );
  OAI22_X1 U2532 ( .A1(n13890), .A2(n13394), .B1(n13390), .B2(n15514), .ZN(
        n7717) );
  OAI22_X1 U2533 ( .A1(n13896), .A2(n13394), .B1(n13391), .B2(n15513), .ZN(
        n7718) );
  OAI22_X1 U2534 ( .A1(n13902), .A2(n13394), .B1(n13391), .B2(n15512), .ZN(
        n7719) );
  OAI22_X1 U2535 ( .A1(n13908), .A2(n13394), .B1(n13391), .B2(n15511), .ZN(
        n7720) );
  OAI22_X1 U2536 ( .A1(n13914), .A2(n13394), .B1(n13391), .B2(n15510), .ZN(
        n7721) );
  OAI22_X1 U2537 ( .A1(n13920), .A2(n13394), .B1(n13391), .B2(n15509), .ZN(
        n7722) );
  OAI22_X1 U2538 ( .A1(n13926), .A2(n13394), .B1(n13391), .B2(n15508), .ZN(
        n7723) );
  OAI22_X1 U2539 ( .A1(n13932), .A2(n13394), .B1(n13391), .B2(n15507), .ZN(
        n7724) );
  OAI22_X1 U2540 ( .A1(n13938), .A2(n13394), .B1(n13391), .B2(n15506), .ZN(
        n7725) );
  OAI22_X1 U2541 ( .A1(n13944), .A2(n13393), .B1(n13391), .B2(n15505), .ZN(
        n7726) );
  OAI22_X1 U2542 ( .A1(n13950), .A2(n13393), .B1(n13391), .B2(n15504), .ZN(
        n7727) );
  OAI22_X1 U2543 ( .A1(n13956), .A2(n13393), .B1(n13391), .B2(n15503), .ZN(
        n7728) );
  OAI22_X1 U2544 ( .A1(n13962), .A2(n13393), .B1(n13391), .B2(n15502), .ZN(
        n7729) );
  OAI22_X1 U2545 ( .A1(n13828), .A2(n13443), .B1(n13438), .B2(n15301), .ZN(
        n7962) );
  OAI22_X1 U2546 ( .A1(n13834), .A2(n13443), .B1(n13438), .B2(n15300), .ZN(
        n7963) );
  OAI22_X1 U2547 ( .A1(n13840), .A2(n13443), .B1(n13438), .B2(n15299), .ZN(
        n7964) );
  OAI22_X1 U2548 ( .A1(n13846), .A2(n13443), .B1(n13438), .B2(n15298), .ZN(
        n7965) );
  OAI22_X1 U2549 ( .A1(n13852), .A2(n13443), .B1(n13438), .B2(n15297), .ZN(
        n7966) );
  OAI22_X1 U2550 ( .A1(n13858), .A2(n13443), .B1(n13438), .B2(n15296), .ZN(
        n7967) );
  OAI22_X1 U2551 ( .A1(n13864), .A2(n13443), .B1(n13438), .B2(n15295), .ZN(
        n7968) );
  OAI22_X1 U2552 ( .A1(n13870), .A2(n13443), .B1(n13438), .B2(n15294), .ZN(
        n7969) );
  OAI22_X1 U2553 ( .A1(n13876), .A2(n13442), .B1(n13438), .B2(n15293), .ZN(
        n7970) );
  OAI22_X1 U2554 ( .A1(n13882), .A2(n13442), .B1(n13438), .B2(n15292), .ZN(
        n7971) );
  OAI22_X1 U2555 ( .A1(n13888), .A2(n13442), .B1(n13438), .B2(n15291), .ZN(
        n7972) );
  OAI22_X1 U2556 ( .A1(n13894), .A2(n13442), .B1(n13438), .B2(n15290), .ZN(
        n7973) );
  OAI22_X1 U2557 ( .A1(n13900), .A2(n13442), .B1(n13439), .B2(n15289), .ZN(
        n7974) );
  OAI22_X1 U2558 ( .A1(n13906), .A2(n13442), .B1(n13439), .B2(n15288), .ZN(
        n7975) );
  OAI22_X1 U2559 ( .A1(n13912), .A2(n13442), .B1(n13439), .B2(n15287), .ZN(
        n7976) );
  OAI22_X1 U2560 ( .A1(n13918), .A2(n13442), .B1(n13439), .B2(n15286), .ZN(
        n7977) );
  OAI22_X1 U2561 ( .A1(n13924), .A2(n13442), .B1(n13439), .B2(n15285), .ZN(
        n7978) );
  OAI22_X1 U2562 ( .A1(n13930), .A2(n13442), .B1(n13439), .B2(n15284), .ZN(
        n7979) );
  OAI22_X1 U2563 ( .A1(n13936), .A2(n13442), .B1(n13439), .B2(n15283), .ZN(
        n7980) );
  OAI22_X1 U2564 ( .A1(n13942), .A2(n13442), .B1(n13439), .B2(n15282), .ZN(
        n7981) );
  OAI22_X1 U2565 ( .A1(n13948), .A2(n13441), .B1(n13439), .B2(n15281), .ZN(
        n7982) );
  OAI22_X1 U2566 ( .A1(n13954), .A2(n13441), .B1(n13439), .B2(n15280), .ZN(
        n7983) );
  OAI22_X1 U2567 ( .A1(n13960), .A2(n13441), .B1(n13439), .B2(n15279), .ZN(
        n7984) );
  OAI22_X1 U2568 ( .A1(n13966), .A2(n13441), .B1(n13439), .B2(n15278), .ZN(
        n7985) );
  OAI22_X1 U2569 ( .A1(n13828), .A2(n13449), .B1(n13444), .B2(n15269), .ZN(
        n7994) );
  OAI22_X1 U2570 ( .A1(n13834), .A2(n13449), .B1(n13444), .B2(n15268), .ZN(
        n7995) );
  OAI22_X1 U2571 ( .A1(n13840), .A2(n13449), .B1(n13444), .B2(n15267), .ZN(
        n7996) );
  OAI22_X1 U2572 ( .A1(n13846), .A2(n13449), .B1(n13444), .B2(n15266), .ZN(
        n7997) );
  OAI22_X1 U2573 ( .A1(n13852), .A2(n13449), .B1(n13444), .B2(n15265), .ZN(
        n7998) );
  OAI22_X1 U2574 ( .A1(n13858), .A2(n13449), .B1(n13444), .B2(n15264), .ZN(
        n7999) );
  OAI22_X1 U2575 ( .A1(n13864), .A2(n13449), .B1(n13444), .B2(n15263), .ZN(
        n8000) );
  OAI22_X1 U2576 ( .A1(n13870), .A2(n13449), .B1(n13444), .B2(n15262), .ZN(
        n8001) );
  OAI22_X1 U2577 ( .A1(n13876), .A2(n13448), .B1(n13444), .B2(n15261), .ZN(
        n8002) );
  OAI22_X1 U2578 ( .A1(n13882), .A2(n13448), .B1(n13444), .B2(n15260), .ZN(
        n8003) );
  OAI22_X1 U2579 ( .A1(n13888), .A2(n13448), .B1(n13444), .B2(n15259), .ZN(
        n8004) );
  OAI22_X1 U2580 ( .A1(n13894), .A2(n13448), .B1(n13444), .B2(n15258), .ZN(
        n8005) );
  OAI22_X1 U2581 ( .A1(n13900), .A2(n13448), .B1(n13445), .B2(n15257), .ZN(
        n8006) );
  OAI22_X1 U2582 ( .A1(n13906), .A2(n13448), .B1(n13445), .B2(n15256), .ZN(
        n8007) );
  OAI22_X1 U2583 ( .A1(n13912), .A2(n13448), .B1(n13445), .B2(n15255), .ZN(
        n8008) );
  OAI22_X1 U2584 ( .A1(n13918), .A2(n13448), .B1(n13445), .B2(n15254), .ZN(
        n8009) );
  OAI22_X1 U2585 ( .A1(n13924), .A2(n13448), .B1(n13445), .B2(n15253), .ZN(
        n8010) );
  OAI22_X1 U2586 ( .A1(n13930), .A2(n13448), .B1(n13445), .B2(n15252), .ZN(
        n8011) );
  OAI22_X1 U2587 ( .A1(n13936), .A2(n13448), .B1(n13445), .B2(n15251), .ZN(
        n8012) );
  OAI22_X1 U2588 ( .A1(n13942), .A2(n13448), .B1(n13445), .B2(n15250), .ZN(
        n8013) );
  OAI22_X1 U2589 ( .A1(n13948), .A2(n13447), .B1(n13445), .B2(n15249), .ZN(
        n8014) );
  OAI22_X1 U2590 ( .A1(n13954), .A2(n13447), .B1(n13445), .B2(n15248), .ZN(
        n8015) );
  OAI22_X1 U2591 ( .A1(n13960), .A2(n13447), .B1(n13445), .B2(n15247), .ZN(
        n8016) );
  OAI22_X1 U2592 ( .A1(n13966), .A2(n13447), .B1(n13445), .B2(n15246), .ZN(
        n8017) );
  OAI22_X1 U2593 ( .A1(n13828), .A2(n13455), .B1(n13450), .B2(n15237), .ZN(
        n8026) );
  OAI22_X1 U2594 ( .A1(n13834), .A2(n13455), .B1(n13450), .B2(n15236), .ZN(
        n8027) );
  OAI22_X1 U2595 ( .A1(n13840), .A2(n13455), .B1(n13450), .B2(n15235), .ZN(
        n8028) );
  OAI22_X1 U2596 ( .A1(n13846), .A2(n13455), .B1(n13450), .B2(n15234), .ZN(
        n8029) );
  OAI22_X1 U2597 ( .A1(n13852), .A2(n13455), .B1(n13450), .B2(n15233), .ZN(
        n8030) );
  OAI22_X1 U2598 ( .A1(n13858), .A2(n13455), .B1(n13450), .B2(n15232), .ZN(
        n8031) );
  OAI22_X1 U2599 ( .A1(n13864), .A2(n13455), .B1(n13450), .B2(n15231), .ZN(
        n8032) );
  OAI22_X1 U2600 ( .A1(n13870), .A2(n13455), .B1(n13450), .B2(n15230), .ZN(
        n8033) );
  OAI22_X1 U2601 ( .A1(n13876), .A2(n13454), .B1(n13450), .B2(n15229), .ZN(
        n8034) );
  OAI22_X1 U2602 ( .A1(n13882), .A2(n13454), .B1(n13450), .B2(n15228), .ZN(
        n8035) );
  OAI22_X1 U2603 ( .A1(n13888), .A2(n13454), .B1(n13450), .B2(n15227), .ZN(
        n8036) );
  OAI22_X1 U2604 ( .A1(n13894), .A2(n13454), .B1(n13450), .B2(n15226), .ZN(
        n8037) );
  OAI22_X1 U2605 ( .A1(n13900), .A2(n13454), .B1(n13451), .B2(n15225), .ZN(
        n8038) );
  OAI22_X1 U2606 ( .A1(n13906), .A2(n13454), .B1(n13451), .B2(n15224), .ZN(
        n8039) );
  OAI22_X1 U2607 ( .A1(n13912), .A2(n13454), .B1(n13451), .B2(n15223), .ZN(
        n8040) );
  OAI22_X1 U2608 ( .A1(n13918), .A2(n13454), .B1(n13451), .B2(n15222), .ZN(
        n8041) );
  OAI22_X1 U2609 ( .A1(n13924), .A2(n13454), .B1(n13451), .B2(n15221), .ZN(
        n8042) );
  OAI22_X1 U2610 ( .A1(n13930), .A2(n13454), .B1(n13451), .B2(n15220), .ZN(
        n8043) );
  OAI22_X1 U2611 ( .A1(n13936), .A2(n13454), .B1(n13451), .B2(n15219), .ZN(
        n8044) );
  OAI22_X1 U2612 ( .A1(n13942), .A2(n13454), .B1(n13451), .B2(n15218), .ZN(
        n8045) );
  OAI22_X1 U2613 ( .A1(n13948), .A2(n13453), .B1(n13451), .B2(n15217), .ZN(
        n8046) );
  OAI22_X1 U2614 ( .A1(n13954), .A2(n13453), .B1(n13451), .B2(n15216), .ZN(
        n8047) );
  OAI22_X1 U2615 ( .A1(n13960), .A2(n13453), .B1(n13451), .B2(n15215), .ZN(
        n8048) );
  OAI22_X1 U2616 ( .A1(n13966), .A2(n13453), .B1(n13451), .B2(n15214), .ZN(
        n8049) );
  OAI22_X1 U2617 ( .A1(n13828), .A2(n13485), .B1(n13480), .B2(n15173), .ZN(
        n8186) );
  OAI22_X1 U2618 ( .A1(n13834), .A2(n13485), .B1(n13480), .B2(n15172), .ZN(
        n8187) );
  OAI22_X1 U2619 ( .A1(n13840), .A2(n13485), .B1(n13480), .B2(n15171), .ZN(
        n8188) );
  OAI22_X1 U2620 ( .A1(n13846), .A2(n13485), .B1(n13480), .B2(n15170), .ZN(
        n8189) );
  OAI22_X1 U2621 ( .A1(n13852), .A2(n13485), .B1(n13480), .B2(n15169), .ZN(
        n8190) );
  OAI22_X1 U2622 ( .A1(n13858), .A2(n13485), .B1(n13480), .B2(n15168), .ZN(
        n8191) );
  OAI22_X1 U2623 ( .A1(n13864), .A2(n13485), .B1(n13480), .B2(n15167), .ZN(
        n8192) );
  OAI22_X1 U2624 ( .A1(n13870), .A2(n13485), .B1(n13480), .B2(n15166), .ZN(
        n8193) );
  OAI22_X1 U2625 ( .A1(n13876), .A2(n13484), .B1(n13480), .B2(n15165), .ZN(
        n8194) );
  OAI22_X1 U2626 ( .A1(n13882), .A2(n13484), .B1(n13480), .B2(n15164), .ZN(
        n8195) );
  OAI22_X1 U2627 ( .A1(n13888), .A2(n13484), .B1(n13480), .B2(n15163), .ZN(
        n8196) );
  OAI22_X1 U2628 ( .A1(n13894), .A2(n13484), .B1(n13480), .B2(n15162), .ZN(
        n8197) );
  OAI22_X1 U2629 ( .A1(n13900), .A2(n13484), .B1(n13481), .B2(n15161), .ZN(
        n8198) );
  OAI22_X1 U2630 ( .A1(n13906), .A2(n13484), .B1(n13481), .B2(n15160), .ZN(
        n8199) );
  OAI22_X1 U2631 ( .A1(n13912), .A2(n13484), .B1(n13481), .B2(n15159), .ZN(
        n8200) );
  OAI22_X1 U2632 ( .A1(n13918), .A2(n13484), .B1(n13481), .B2(n15158), .ZN(
        n8201) );
  OAI22_X1 U2633 ( .A1(n13924), .A2(n13484), .B1(n13481), .B2(n15157), .ZN(
        n8202) );
  OAI22_X1 U2634 ( .A1(n13930), .A2(n13484), .B1(n13481), .B2(n15156), .ZN(
        n8203) );
  OAI22_X1 U2635 ( .A1(n13936), .A2(n13484), .B1(n13481), .B2(n15155), .ZN(
        n8204) );
  OAI22_X1 U2636 ( .A1(n13942), .A2(n13484), .B1(n13481), .B2(n15154), .ZN(
        n8205) );
  OAI22_X1 U2637 ( .A1(n13948), .A2(n13483), .B1(n13481), .B2(n15153), .ZN(
        n8206) );
  OAI22_X1 U2638 ( .A1(n13954), .A2(n13483), .B1(n13481), .B2(n15152), .ZN(
        n8207) );
  OAI22_X1 U2639 ( .A1(n13960), .A2(n13483), .B1(n13481), .B2(n15151), .ZN(
        n8208) );
  OAI22_X1 U2640 ( .A1(n13966), .A2(n13483), .B1(n13481), .B2(n15150), .ZN(
        n8209) );
  OAI22_X1 U2641 ( .A1(n13828), .A2(n13491), .B1(n13486), .B2(n15141), .ZN(
        n8218) );
  OAI22_X1 U2642 ( .A1(n13834), .A2(n13491), .B1(n13486), .B2(n15140), .ZN(
        n8219) );
  OAI22_X1 U2643 ( .A1(n13840), .A2(n13491), .B1(n13486), .B2(n15139), .ZN(
        n8220) );
  OAI22_X1 U2644 ( .A1(n13846), .A2(n13491), .B1(n13486), .B2(n15138), .ZN(
        n8221) );
  OAI22_X1 U2645 ( .A1(n13852), .A2(n13491), .B1(n13486), .B2(n15137), .ZN(
        n8222) );
  OAI22_X1 U2646 ( .A1(n13858), .A2(n13491), .B1(n13486), .B2(n15136), .ZN(
        n8223) );
  OAI22_X1 U2647 ( .A1(n13864), .A2(n13491), .B1(n13486), .B2(n15135), .ZN(
        n8224) );
  OAI22_X1 U2648 ( .A1(n13870), .A2(n13491), .B1(n13486), .B2(n15134), .ZN(
        n8225) );
  OAI22_X1 U2649 ( .A1(n13876), .A2(n13490), .B1(n13486), .B2(n15133), .ZN(
        n8226) );
  OAI22_X1 U2650 ( .A1(n13882), .A2(n13490), .B1(n13486), .B2(n15132), .ZN(
        n8227) );
  OAI22_X1 U2651 ( .A1(n13888), .A2(n13490), .B1(n13486), .B2(n15131), .ZN(
        n8228) );
  OAI22_X1 U2652 ( .A1(n13894), .A2(n13490), .B1(n13486), .B2(n15130), .ZN(
        n8229) );
  OAI22_X1 U2653 ( .A1(n13900), .A2(n13490), .B1(n13487), .B2(n15129), .ZN(
        n8230) );
  OAI22_X1 U2654 ( .A1(n13906), .A2(n13490), .B1(n13487), .B2(n15128), .ZN(
        n8231) );
  OAI22_X1 U2655 ( .A1(n13912), .A2(n13490), .B1(n13487), .B2(n15127), .ZN(
        n8232) );
  OAI22_X1 U2656 ( .A1(n13918), .A2(n13490), .B1(n13487), .B2(n15126), .ZN(
        n8233) );
  OAI22_X1 U2657 ( .A1(n13924), .A2(n13490), .B1(n13487), .B2(n15125), .ZN(
        n8234) );
  OAI22_X1 U2658 ( .A1(n13930), .A2(n13490), .B1(n13487), .B2(n15124), .ZN(
        n8235) );
  OAI22_X1 U2659 ( .A1(n13936), .A2(n13490), .B1(n13487), .B2(n15123), .ZN(
        n8236) );
  OAI22_X1 U2660 ( .A1(n13942), .A2(n13490), .B1(n13487), .B2(n15122), .ZN(
        n8237) );
  OAI22_X1 U2661 ( .A1(n13948), .A2(n13489), .B1(n13487), .B2(n15121), .ZN(
        n8238) );
  OAI22_X1 U2662 ( .A1(n13954), .A2(n13489), .B1(n13487), .B2(n15120), .ZN(
        n8239) );
  OAI22_X1 U2663 ( .A1(n13960), .A2(n13489), .B1(n13487), .B2(n15119), .ZN(
        n8240) );
  OAI22_X1 U2664 ( .A1(n13966), .A2(n13489), .B1(n13487), .B2(n15118), .ZN(
        n8241) );
  OAI22_X1 U2665 ( .A1(n13828), .A2(n13497), .B1(n13492), .B2(n15109), .ZN(
        n8250) );
  OAI22_X1 U2666 ( .A1(n13834), .A2(n13497), .B1(n13492), .B2(n15108), .ZN(
        n8251) );
  OAI22_X1 U2667 ( .A1(n13840), .A2(n13497), .B1(n13492), .B2(n15107), .ZN(
        n8252) );
  OAI22_X1 U2668 ( .A1(n13846), .A2(n13497), .B1(n13492), .B2(n15106), .ZN(
        n8253) );
  OAI22_X1 U2669 ( .A1(n13852), .A2(n13497), .B1(n13492), .B2(n15105), .ZN(
        n8254) );
  OAI22_X1 U2670 ( .A1(n13858), .A2(n13497), .B1(n13492), .B2(n15104), .ZN(
        n8255) );
  OAI22_X1 U2671 ( .A1(n13864), .A2(n13497), .B1(n13492), .B2(n15103), .ZN(
        n8256) );
  OAI22_X1 U2672 ( .A1(n13870), .A2(n13497), .B1(n13492), .B2(n15102), .ZN(
        n8257) );
  OAI22_X1 U2673 ( .A1(n13876), .A2(n13496), .B1(n13492), .B2(n15101), .ZN(
        n8258) );
  OAI22_X1 U2674 ( .A1(n13882), .A2(n13496), .B1(n13492), .B2(n15100), .ZN(
        n8259) );
  OAI22_X1 U2675 ( .A1(n13888), .A2(n13496), .B1(n13492), .B2(n15099), .ZN(
        n8260) );
  OAI22_X1 U2676 ( .A1(n13894), .A2(n13496), .B1(n13492), .B2(n15098), .ZN(
        n8261) );
  OAI22_X1 U2677 ( .A1(n13900), .A2(n13496), .B1(n13493), .B2(n15097), .ZN(
        n8262) );
  OAI22_X1 U2678 ( .A1(n13906), .A2(n13496), .B1(n13493), .B2(n15096), .ZN(
        n8263) );
  OAI22_X1 U2679 ( .A1(n13912), .A2(n13496), .B1(n13493), .B2(n15095), .ZN(
        n8264) );
  OAI22_X1 U2680 ( .A1(n13918), .A2(n13496), .B1(n13493), .B2(n15094), .ZN(
        n8265) );
  OAI22_X1 U2681 ( .A1(n13924), .A2(n13496), .B1(n13493), .B2(n15093), .ZN(
        n8266) );
  OAI22_X1 U2682 ( .A1(n13930), .A2(n13496), .B1(n13493), .B2(n15092), .ZN(
        n8267) );
  OAI22_X1 U2683 ( .A1(n13936), .A2(n13496), .B1(n13493), .B2(n15091), .ZN(
        n8268) );
  OAI22_X1 U2684 ( .A1(n13942), .A2(n13496), .B1(n13493), .B2(n15090), .ZN(
        n8269) );
  OAI22_X1 U2685 ( .A1(n13948), .A2(n13495), .B1(n13493), .B2(n15089), .ZN(
        n8270) );
  OAI22_X1 U2686 ( .A1(n13954), .A2(n13495), .B1(n13493), .B2(n15088), .ZN(
        n8271) );
  OAI22_X1 U2687 ( .A1(n13960), .A2(n13495), .B1(n13493), .B2(n15087), .ZN(
        n8272) );
  OAI22_X1 U2688 ( .A1(n13966), .A2(n13495), .B1(n13493), .B2(n15086), .ZN(
        n8273) );
  OAI22_X1 U2689 ( .A1(n13828), .A2(n13503), .B1(n13498), .B2(n15077), .ZN(
        n8282) );
  OAI22_X1 U2690 ( .A1(n13834), .A2(n13503), .B1(n13498), .B2(n15076), .ZN(
        n8283) );
  OAI22_X1 U2691 ( .A1(n13840), .A2(n13503), .B1(n13498), .B2(n15075), .ZN(
        n8284) );
  OAI22_X1 U2692 ( .A1(n13846), .A2(n13503), .B1(n13498), .B2(n15074), .ZN(
        n8285) );
  OAI22_X1 U2693 ( .A1(n13852), .A2(n13503), .B1(n13498), .B2(n15073), .ZN(
        n8286) );
  OAI22_X1 U2694 ( .A1(n13858), .A2(n13503), .B1(n13498), .B2(n15072), .ZN(
        n8287) );
  OAI22_X1 U2695 ( .A1(n13864), .A2(n13503), .B1(n13498), .B2(n15071), .ZN(
        n8288) );
  OAI22_X1 U2696 ( .A1(n13870), .A2(n13503), .B1(n13498), .B2(n15070), .ZN(
        n8289) );
  OAI22_X1 U2697 ( .A1(n13876), .A2(n13502), .B1(n13498), .B2(n15069), .ZN(
        n8290) );
  OAI22_X1 U2698 ( .A1(n13882), .A2(n13502), .B1(n13498), .B2(n15068), .ZN(
        n8291) );
  OAI22_X1 U2699 ( .A1(n13888), .A2(n13502), .B1(n13498), .B2(n15067), .ZN(
        n8292) );
  OAI22_X1 U2700 ( .A1(n13894), .A2(n13502), .B1(n13498), .B2(n15066), .ZN(
        n8293) );
  OAI22_X1 U2701 ( .A1(n13900), .A2(n13502), .B1(n13499), .B2(n15065), .ZN(
        n8294) );
  OAI22_X1 U2702 ( .A1(n13906), .A2(n13502), .B1(n13499), .B2(n15064), .ZN(
        n8295) );
  OAI22_X1 U2703 ( .A1(n13912), .A2(n13502), .B1(n13499), .B2(n15063), .ZN(
        n8296) );
  OAI22_X1 U2704 ( .A1(n13918), .A2(n13502), .B1(n13499), .B2(n15062), .ZN(
        n8297) );
  OAI22_X1 U2705 ( .A1(n13924), .A2(n13502), .B1(n13499), .B2(n15061), .ZN(
        n8298) );
  OAI22_X1 U2706 ( .A1(n13930), .A2(n13502), .B1(n13499), .B2(n15060), .ZN(
        n8299) );
  OAI22_X1 U2707 ( .A1(n13936), .A2(n13502), .B1(n13499), .B2(n15059), .ZN(
        n8300) );
  OAI22_X1 U2708 ( .A1(n13942), .A2(n13502), .B1(n13499), .B2(n15058), .ZN(
        n8301) );
  OAI22_X1 U2709 ( .A1(n13948), .A2(n13501), .B1(n13499), .B2(n15057), .ZN(
        n8302) );
  OAI22_X1 U2710 ( .A1(n13954), .A2(n13501), .B1(n13499), .B2(n15056), .ZN(
        n8303) );
  OAI22_X1 U2711 ( .A1(n13960), .A2(n13501), .B1(n13499), .B2(n15055), .ZN(
        n8304) );
  OAI22_X1 U2712 ( .A1(n13966), .A2(n13501), .B1(n13499), .B2(n15054), .ZN(
        n8305) );
  OAI22_X1 U2713 ( .A1(n13827), .A2(n13509), .B1(n13504), .B2(n15045), .ZN(
        n8314) );
  OAI22_X1 U2714 ( .A1(n13834), .A2(n13509), .B1(n13504), .B2(n15044), .ZN(
        n8315) );
  OAI22_X1 U2715 ( .A1(n13840), .A2(n13509), .B1(n13504), .B2(n15043), .ZN(
        n8316) );
  OAI22_X1 U2716 ( .A1(n13846), .A2(n13509), .B1(n13504), .B2(n15042), .ZN(
        n8317) );
  OAI22_X1 U2717 ( .A1(n13852), .A2(n13509), .B1(n13504), .B2(n15041), .ZN(
        n8318) );
  OAI22_X1 U2718 ( .A1(n13858), .A2(n13509), .B1(n13504), .B2(n15040), .ZN(
        n8319) );
  OAI22_X1 U2719 ( .A1(n13864), .A2(n13509), .B1(n13504), .B2(n15039), .ZN(
        n8320) );
  OAI22_X1 U2720 ( .A1(n13870), .A2(n13509), .B1(n13504), .B2(n15038), .ZN(
        n8321) );
  OAI22_X1 U2721 ( .A1(n13876), .A2(n13508), .B1(n13504), .B2(n15037), .ZN(
        n8322) );
  OAI22_X1 U2722 ( .A1(n13882), .A2(n13508), .B1(n13504), .B2(n15036), .ZN(
        n8323) );
  OAI22_X1 U2723 ( .A1(n13888), .A2(n13508), .B1(n13504), .B2(n15035), .ZN(
        n8324) );
  OAI22_X1 U2724 ( .A1(n13894), .A2(n13508), .B1(n13504), .B2(n15034), .ZN(
        n8325) );
  OAI22_X1 U2725 ( .A1(n13900), .A2(n13508), .B1(n13505), .B2(n15033), .ZN(
        n8326) );
  OAI22_X1 U2726 ( .A1(n13906), .A2(n13508), .B1(n13505), .B2(n15032), .ZN(
        n8327) );
  OAI22_X1 U2727 ( .A1(n13912), .A2(n13508), .B1(n13505), .B2(n15031), .ZN(
        n8328) );
  OAI22_X1 U2728 ( .A1(n13918), .A2(n13508), .B1(n13505), .B2(n15030), .ZN(
        n8329) );
  OAI22_X1 U2729 ( .A1(n13924), .A2(n13508), .B1(n13505), .B2(n15029), .ZN(
        n8330) );
  OAI22_X1 U2730 ( .A1(n13930), .A2(n13508), .B1(n13505), .B2(n15028), .ZN(
        n8331) );
  OAI22_X1 U2731 ( .A1(n13936), .A2(n13508), .B1(n13505), .B2(n15027), .ZN(
        n8332) );
  OAI22_X1 U2732 ( .A1(n13942), .A2(n13508), .B1(n13505), .B2(n15026), .ZN(
        n8333) );
  OAI22_X1 U2733 ( .A1(n13948), .A2(n13507), .B1(n13505), .B2(n15025), .ZN(
        n8334) );
  OAI22_X1 U2734 ( .A1(n13954), .A2(n13507), .B1(n13505), .B2(n15024), .ZN(
        n8335) );
  OAI22_X1 U2735 ( .A1(n13960), .A2(n13507), .B1(n13505), .B2(n15023), .ZN(
        n8336) );
  OAI22_X1 U2736 ( .A1(n13966), .A2(n13507), .B1(n13505), .B2(n15022), .ZN(
        n8337) );
  OAI22_X1 U2737 ( .A1(n13827), .A2(n13533), .B1(n13528), .B2(n14980), .ZN(
        n8442) );
  OAI22_X1 U2738 ( .A1(n13833), .A2(n13533), .B1(n13528), .B2(n14979), .ZN(
        n8443) );
  OAI22_X1 U2739 ( .A1(n13839), .A2(n13533), .B1(n13528), .B2(n14978), .ZN(
        n8444) );
  OAI22_X1 U2740 ( .A1(n13845), .A2(n13533), .B1(n13528), .B2(n14977), .ZN(
        n8445) );
  OAI22_X1 U2741 ( .A1(n13851), .A2(n13533), .B1(n13528), .B2(n14976), .ZN(
        n8446) );
  OAI22_X1 U2742 ( .A1(n13857), .A2(n13533), .B1(n13528), .B2(n14975), .ZN(
        n8447) );
  OAI22_X1 U2743 ( .A1(n13863), .A2(n13533), .B1(n13528), .B2(n14974), .ZN(
        n8448) );
  OAI22_X1 U2744 ( .A1(n13869), .A2(n13533), .B1(n13528), .B2(n14973), .ZN(
        n8449) );
  OAI22_X1 U2745 ( .A1(n13875), .A2(n13532), .B1(n13528), .B2(n14972), .ZN(
        n8450) );
  OAI22_X1 U2746 ( .A1(n13881), .A2(n13532), .B1(n13528), .B2(n14971), .ZN(
        n8451) );
  OAI22_X1 U2747 ( .A1(n13887), .A2(n13532), .B1(n13528), .B2(n14970), .ZN(
        n8452) );
  OAI22_X1 U2748 ( .A1(n13893), .A2(n13532), .B1(n13528), .B2(n14969), .ZN(
        n8453) );
  OAI22_X1 U2749 ( .A1(n13899), .A2(n13532), .B1(n13529), .B2(n14968), .ZN(
        n8454) );
  OAI22_X1 U2750 ( .A1(n13905), .A2(n13532), .B1(n13529), .B2(n14967), .ZN(
        n8455) );
  OAI22_X1 U2751 ( .A1(n13911), .A2(n13532), .B1(n13529), .B2(n14966), .ZN(
        n8456) );
  OAI22_X1 U2752 ( .A1(n13917), .A2(n13532), .B1(n13529), .B2(n14965), .ZN(
        n8457) );
  OAI22_X1 U2753 ( .A1(n13923), .A2(n13532), .B1(n13529), .B2(n14964), .ZN(
        n8458) );
  OAI22_X1 U2754 ( .A1(n13929), .A2(n13532), .B1(n13529), .B2(n14963), .ZN(
        n8459) );
  OAI22_X1 U2755 ( .A1(n13935), .A2(n13532), .B1(n13529), .B2(n14962), .ZN(
        n8460) );
  OAI22_X1 U2756 ( .A1(n13941), .A2(n13532), .B1(n13529), .B2(n14961), .ZN(
        n8461) );
  OAI22_X1 U2757 ( .A1(n13947), .A2(n13531), .B1(n13529), .B2(n14960), .ZN(
        n8462) );
  OAI22_X1 U2758 ( .A1(n13953), .A2(n13531), .B1(n13529), .B2(n14959), .ZN(
        n8463) );
  OAI22_X1 U2759 ( .A1(n13959), .A2(n13531), .B1(n13529), .B2(n14958), .ZN(
        n8464) );
  OAI22_X1 U2760 ( .A1(n13965), .A2(n13531), .B1(n13529), .B2(n14957), .ZN(
        n8465) );
  OAI22_X1 U2761 ( .A1(n13827), .A2(n13551), .B1(n13546), .B2(n14947), .ZN(
        n8538) );
  OAI22_X1 U2762 ( .A1(n13833), .A2(n13551), .B1(n13546), .B2(n14946), .ZN(
        n8539) );
  OAI22_X1 U2763 ( .A1(n13839), .A2(n13551), .B1(n13546), .B2(n14945), .ZN(
        n8540) );
  OAI22_X1 U2764 ( .A1(n13845), .A2(n13551), .B1(n13546), .B2(n14944), .ZN(
        n8541) );
  OAI22_X1 U2765 ( .A1(n13851), .A2(n13551), .B1(n13546), .B2(n14943), .ZN(
        n8542) );
  OAI22_X1 U2766 ( .A1(n13857), .A2(n13551), .B1(n13546), .B2(n14942), .ZN(
        n8543) );
  OAI22_X1 U2767 ( .A1(n13863), .A2(n13551), .B1(n13546), .B2(n14941), .ZN(
        n8544) );
  OAI22_X1 U2768 ( .A1(n13869), .A2(n13551), .B1(n13546), .B2(n14940), .ZN(
        n8545) );
  OAI22_X1 U2769 ( .A1(n13875), .A2(n13550), .B1(n13546), .B2(n14939), .ZN(
        n8546) );
  OAI22_X1 U2770 ( .A1(n13881), .A2(n13550), .B1(n13546), .B2(n14938), .ZN(
        n8547) );
  OAI22_X1 U2771 ( .A1(n13887), .A2(n13550), .B1(n13546), .B2(n14937), .ZN(
        n8548) );
  OAI22_X1 U2772 ( .A1(n13893), .A2(n13550), .B1(n13546), .B2(n14936), .ZN(
        n8549) );
  OAI22_X1 U2773 ( .A1(n13899), .A2(n13550), .B1(n13547), .B2(n14935), .ZN(
        n8550) );
  OAI22_X1 U2774 ( .A1(n13905), .A2(n13550), .B1(n13547), .B2(n14934), .ZN(
        n8551) );
  OAI22_X1 U2775 ( .A1(n13911), .A2(n13550), .B1(n13547), .B2(n14933), .ZN(
        n8552) );
  OAI22_X1 U2776 ( .A1(n13917), .A2(n13550), .B1(n13547), .B2(n14932), .ZN(
        n8553) );
  OAI22_X1 U2777 ( .A1(n13923), .A2(n13550), .B1(n13547), .B2(n14931), .ZN(
        n8554) );
  OAI22_X1 U2778 ( .A1(n13929), .A2(n13550), .B1(n13547), .B2(n14930), .ZN(
        n8555) );
  OAI22_X1 U2779 ( .A1(n13935), .A2(n13550), .B1(n13547), .B2(n14929), .ZN(
        n8556) );
  OAI22_X1 U2780 ( .A1(n13941), .A2(n13550), .B1(n13547), .B2(n14928), .ZN(
        n8557) );
  OAI22_X1 U2781 ( .A1(n13947), .A2(n13549), .B1(n13547), .B2(n14927), .ZN(
        n8558) );
  OAI22_X1 U2782 ( .A1(n13953), .A2(n13549), .B1(n13547), .B2(n14926), .ZN(
        n8559) );
  OAI22_X1 U2783 ( .A1(n13959), .A2(n13549), .B1(n13547), .B2(n14925), .ZN(
        n8560) );
  OAI22_X1 U2784 ( .A1(n13965), .A2(n13549), .B1(n13547), .B2(n14924), .ZN(
        n8561) );
  OAI22_X1 U2785 ( .A1(n13827), .A2(n13557), .B1(n13552), .B2(n14915), .ZN(
        n8570) );
  OAI22_X1 U2786 ( .A1(n13833), .A2(n13557), .B1(n13552), .B2(n14914), .ZN(
        n8571) );
  OAI22_X1 U2787 ( .A1(n13839), .A2(n13557), .B1(n13552), .B2(n14913), .ZN(
        n8572) );
  OAI22_X1 U2788 ( .A1(n13845), .A2(n13557), .B1(n13552), .B2(n14912), .ZN(
        n8573) );
  OAI22_X1 U2789 ( .A1(n13851), .A2(n13557), .B1(n13552), .B2(n14911), .ZN(
        n8574) );
  OAI22_X1 U2790 ( .A1(n13857), .A2(n13557), .B1(n13552), .B2(n14910), .ZN(
        n8575) );
  OAI22_X1 U2791 ( .A1(n13863), .A2(n13557), .B1(n13552), .B2(n14909), .ZN(
        n8576) );
  OAI22_X1 U2792 ( .A1(n13869), .A2(n13557), .B1(n13552), .B2(n14908), .ZN(
        n8577) );
  OAI22_X1 U2793 ( .A1(n13875), .A2(n13556), .B1(n13552), .B2(n14907), .ZN(
        n8578) );
  OAI22_X1 U2794 ( .A1(n13881), .A2(n13556), .B1(n13552), .B2(n14906), .ZN(
        n8579) );
  OAI22_X1 U2795 ( .A1(n13887), .A2(n13556), .B1(n13552), .B2(n14905), .ZN(
        n8580) );
  OAI22_X1 U2796 ( .A1(n13893), .A2(n13556), .B1(n13552), .B2(n14904), .ZN(
        n8581) );
  OAI22_X1 U2797 ( .A1(n13899), .A2(n13556), .B1(n13553), .B2(n14903), .ZN(
        n8582) );
  OAI22_X1 U2798 ( .A1(n13905), .A2(n13556), .B1(n13553), .B2(n14902), .ZN(
        n8583) );
  OAI22_X1 U2799 ( .A1(n13911), .A2(n13556), .B1(n13553), .B2(n14901), .ZN(
        n8584) );
  OAI22_X1 U2800 ( .A1(n13917), .A2(n13556), .B1(n13553), .B2(n14900), .ZN(
        n8585) );
  OAI22_X1 U2801 ( .A1(n13923), .A2(n13556), .B1(n13553), .B2(n14899), .ZN(
        n8586) );
  OAI22_X1 U2802 ( .A1(n13929), .A2(n13556), .B1(n13553), .B2(n14898), .ZN(
        n8587) );
  OAI22_X1 U2803 ( .A1(n13935), .A2(n13556), .B1(n13553), .B2(n14897), .ZN(
        n8588) );
  OAI22_X1 U2804 ( .A1(n13941), .A2(n13556), .B1(n13553), .B2(n14896), .ZN(
        n8589) );
  OAI22_X1 U2805 ( .A1(n13947), .A2(n13555), .B1(n13553), .B2(n14895), .ZN(
        n8590) );
  OAI22_X1 U2806 ( .A1(n13953), .A2(n13555), .B1(n13553), .B2(n14894), .ZN(
        n8591) );
  OAI22_X1 U2807 ( .A1(n13959), .A2(n13555), .B1(n13553), .B2(n14893), .ZN(
        n8592) );
  OAI22_X1 U2808 ( .A1(n13965), .A2(n13555), .B1(n13553), .B2(n14892), .ZN(
        n8593) );
  OAI22_X1 U2809 ( .A1(n13827), .A2(n13563), .B1(n13558), .B2(n14883), .ZN(
        n8602) );
  OAI22_X1 U2810 ( .A1(n13833), .A2(n13563), .B1(n13558), .B2(n14882), .ZN(
        n8603) );
  OAI22_X1 U2811 ( .A1(n13839), .A2(n13563), .B1(n13558), .B2(n14881), .ZN(
        n8604) );
  OAI22_X1 U2812 ( .A1(n13845), .A2(n13563), .B1(n13558), .B2(n14880), .ZN(
        n8605) );
  OAI22_X1 U2813 ( .A1(n13851), .A2(n13563), .B1(n13558), .B2(n14879), .ZN(
        n8606) );
  OAI22_X1 U2814 ( .A1(n13857), .A2(n13563), .B1(n13558), .B2(n14878), .ZN(
        n8607) );
  OAI22_X1 U2815 ( .A1(n13863), .A2(n13563), .B1(n13558), .B2(n14877), .ZN(
        n8608) );
  OAI22_X1 U2816 ( .A1(n13869), .A2(n13563), .B1(n13558), .B2(n14876), .ZN(
        n8609) );
  OAI22_X1 U2817 ( .A1(n13875), .A2(n13562), .B1(n13558), .B2(n14875), .ZN(
        n8610) );
  OAI22_X1 U2818 ( .A1(n13881), .A2(n13562), .B1(n13558), .B2(n14874), .ZN(
        n8611) );
  OAI22_X1 U2819 ( .A1(n13887), .A2(n13562), .B1(n13558), .B2(n14873), .ZN(
        n8612) );
  OAI22_X1 U2820 ( .A1(n13893), .A2(n13562), .B1(n13558), .B2(n14872), .ZN(
        n8613) );
  OAI22_X1 U2821 ( .A1(n13899), .A2(n13562), .B1(n13559), .B2(n14871), .ZN(
        n8614) );
  OAI22_X1 U2822 ( .A1(n13905), .A2(n13562), .B1(n13559), .B2(n14870), .ZN(
        n8615) );
  OAI22_X1 U2823 ( .A1(n13911), .A2(n13562), .B1(n13559), .B2(n14869), .ZN(
        n8616) );
  OAI22_X1 U2824 ( .A1(n13917), .A2(n13562), .B1(n13559), .B2(n14868), .ZN(
        n8617) );
  OAI22_X1 U2825 ( .A1(n13923), .A2(n13562), .B1(n13559), .B2(n14867), .ZN(
        n8618) );
  OAI22_X1 U2826 ( .A1(n13929), .A2(n13562), .B1(n13559), .B2(n14866), .ZN(
        n8619) );
  OAI22_X1 U2827 ( .A1(n13935), .A2(n13562), .B1(n13559), .B2(n14865), .ZN(
        n8620) );
  OAI22_X1 U2828 ( .A1(n13941), .A2(n13562), .B1(n13559), .B2(n14864), .ZN(
        n8621) );
  OAI22_X1 U2829 ( .A1(n13947), .A2(n13561), .B1(n13559), .B2(n14863), .ZN(
        n8622) );
  OAI22_X1 U2830 ( .A1(n13953), .A2(n13561), .B1(n13559), .B2(n14862), .ZN(
        n8623) );
  OAI22_X1 U2831 ( .A1(n13959), .A2(n13561), .B1(n13559), .B2(n14861), .ZN(
        n8624) );
  OAI22_X1 U2832 ( .A1(n13965), .A2(n13561), .B1(n13559), .B2(n14860), .ZN(
        n8625) );
  OAI22_X1 U2833 ( .A1(n13826), .A2(n13593), .B1(n13588), .B2(n14851), .ZN(
        n8762) );
  OAI22_X1 U2834 ( .A1(n13833), .A2(n13593), .B1(n13588), .B2(n14850), .ZN(
        n8763) );
  OAI22_X1 U2835 ( .A1(n13839), .A2(n13593), .B1(n13588), .B2(n14849), .ZN(
        n8764) );
  OAI22_X1 U2836 ( .A1(n13845), .A2(n13593), .B1(n13588), .B2(n14848), .ZN(
        n8765) );
  OAI22_X1 U2837 ( .A1(n13851), .A2(n13593), .B1(n13588), .B2(n14847), .ZN(
        n8766) );
  OAI22_X1 U2838 ( .A1(n13857), .A2(n13593), .B1(n13588), .B2(n14846), .ZN(
        n8767) );
  OAI22_X1 U2839 ( .A1(n13863), .A2(n13593), .B1(n13588), .B2(n14845), .ZN(
        n8768) );
  OAI22_X1 U2840 ( .A1(n13869), .A2(n13593), .B1(n13588), .B2(n14844), .ZN(
        n8769) );
  OAI22_X1 U2841 ( .A1(n13875), .A2(n13592), .B1(n13588), .B2(n14843), .ZN(
        n8770) );
  OAI22_X1 U2842 ( .A1(n13881), .A2(n13592), .B1(n13588), .B2(n14842), .ZN(
        n8771) );
  OAI22_X1 U2843 ( .A1(n13887), .A2(n13592), .B1(n13588), .B2(n14841), .ZN(
        n8772) );
  OAI22_X1 U2844 ( .A1(n13893), .A2(n13592), .B1(n13588), .B2(n14840), .ZN(
        n8773) );
  OAI22_X1 U2845 ( .A1(n13899), .A2(n13592), .B1(n13589), .B2(n14839), .ZN(
        n8774) );
  OAI22_X1 U2846 ( .A1(n13905), .A2(n13592), .B1(n13589), .B2(n14838), .ZN(
        n8775) );
  OAI22_X1 U2847 ( .A1(n13911), .A2(n13592), .B1(n13589), .B2(n14837), .ZN(
        n8776) );
  OAI22_X1 U2848 ( .A1(n13917), .A2(n13592), .B1(n13589), .B2(n14836), .ZN(
        n8777) );
  OAI22_X1 U2849 ( .A1(n13923), .A2(n13592), .B1(n13589), .B2(n14835), .ZN(
        n8778) );
  OAI22_X1 U2850 ( .A1(n13929), .A2(n13592), .B1(n13589), .B2(n14834), .ZN(
        n8779) );
  OAI22_X1 U2851 ( .A1(n13935), .A2(n13592), .B1(n13589), .B2(n14833), .ZN(
        n8780) );
  OAI22_X1 U2852 ( .A1(n13941), .A2(n13592), .B1(n13589), .B2(n14832), .ZN(
        n8781) );
  OAI22_X1 U2853 ( .A1(n13947), .A2(n13591), .B1(n13589), .B2(n14831), .ZN(
        n8782) );
  OAI22_X1 U2854 ( .A1(n13953), .A2(n13591), .B1(n13589), .B2(n14830), .ZN(
        n8783) );
  OAI22_X1 U2855 ( .A1(n13959), .A2(n13591), .B1(n13589), .B2(n14829), .ZN(
        n8784) );
  OAI22_X1 U2856 ( .A1(n13965), .A2(n13591), .B1(n13589), .B2(n14828), .ZN(
        n8785) );
  OAI22_X1 U2857 ( .A1(n13826), .A2(n13599), .B1(n13594), .B2(n14819), .ZN(
        n8794) );
  OAI22_X1 U2858 ( .A1(n13832), .A2(n13599), .B1(n13594), .B2(n14818), .ZN(
        n8795) );
  OAI22_X1 U2859 ( .A1(n13838), .A2(n13599), .B1(n13594), .B2(n14817), .ZN(
        n8796) );
  OAI22_X1 U2860 ( .A1(n13844), .A2(n13599), .B1(n13594), .B2(n14816), .ZN(
        n8797) );
  OAI22_X1 U2861 ( .A1(n13850), .A2(n13599), .B1(n13594), .B2(n14815), .ZN(
        n8798) );
  OAI22_X1 U2862 ( .A1(n13856), .A2(n13599), .B1(n13594), .B2(n14814), .ZN(
        n8799) );
  OAI22_X1 U2863 ( .A1(n13862), .A2(n13599), .B1(n13594), .B2(n14813), .ZN(
        n8800) );
  OAI22_X1 U2864 ( .A1(n13868), .A2(n13599), .B1(n13594), .B2(n14812), .ZN(
        n8801) );
  OAI22_X1 U2865 ( .A1(n13874), .A2(n13598), .B1(n13594), .B2(n14811), .ZN(
        n8802) );
  OAI22_X1 U2866 ( .A1(n13880), .A2(n13598), .B1(n13594), .B2(n14810), .ZN(
        n8803) );
  OAI22_X1 U2867 ( .A1(n13886), .A2(n13598), .B1(n13594), .B2(n14809), .ZN(
        n8804) );
  OAI22_X1 U2868 ( .A1(n13892), .A2(n13598), .B1(n13594), .B2(n14808), .ZN(
        n8805) );
  OAI22_X1 U2869 ( .A1(n13898), .A2(n13598), .B1(n13595), .B2(n14807), .ZN(
        n8806) );
  OAI22_X1 U2870 ( .A1(n13904), .A2(n13598), .B1(n13595), .B2(n14806), .ZN(
        n8807) );
  OAI22_X1 U2871 ( .A1(n13910), .A2(n13598), .B1(n13595), .B2(n14805), .ZN(
        n8808) );
  OAI22_X1 U2872 ( .A1(n13916), .A2(n13598), .B1(n13595), .B2(n14804), .ZN(
        n8809) );
  OAI22_X1 U2873 ( .A1(n13922), .A2(n13598), .B1(n13595), .B2(n14803), .ZN(
        n8810) );
  OAI22_X1 U2874 ( .A1(n13928), .A2(n13598), .B1(n13595), .B2(n14802), .ZN(
        n8811) );
  OAI22_X1 U2875 ( .A1(n13934), .A2(n13598), .B1(n13595), .B2(n14801), .ZN(
        n8812) );
  OAI22_X1 U2876 ( .A1(n13940), .A2(n13598), .B1(n13595), .B2(n14800), .ZN(
        n8813) );
  OAI22_X1 U2877 ( .A1(n13946), .A2(n13597), .B1(n13595), .B2(n14799), .ZN(
        n8814) );
  OAI22_X1 U2878 ( .A1(n13952), .A2(n13597), .B1(n13595), .B2(n14798), .ZN(
        n8815) );
  OAI22_X1 U2879 ( .A1(n13958), .A2(n13597), .B1(n13595), .B2(n14797), .ZN(
        n8816) );
  OAI22_X1 U2880 ( .A1(n13964), .A2(n13597), .B1(n13595), .B2(n14796), .ZN(
        n8817) );
  OAI22_X1 U2881 ( .A1(n13826), .A2(n13605), .B1(n13600), .B2(n14787), .ZN(
        n8826) );
  OAI22_X1 U2882 ( .A1(n13832), .A2(n13605), .B1(n13600), .B2(n14786), .ZN(
        n8827) );
  OAI22_X1 U2883 ( .A1(n13838), .A2(n13605), .B1(n13600), .B2(n14785), .ZN(
        n8828) );
  OAI22_X1 U2884 ( .A1(n13844), .A2(n13605), .B1(n13600), .B2(n14784), .ZN(
        n8829) );
  OAI22_X1 U2885 ( .A1(n13850), .A2(n13605), .B1(n13600), .B2(n14783), .ZN(
        n8830) );
  OAI22_X1 U2886 ( .A1(n13856), .A2(n13605), .B1(n13600), .B2(n14782), .ZN(
        n8831) );
  OAI22_X1 U2887 ( .A1(n13862), .A2(n13605), .B1(n13600), .B2(n14781), .ZN(
        n8832) );
  OAI22_X1 U2888 ( .A1(n13868), .A2(n13605), .B1(n13600), .B2(n14780), .ZN(
        n8833) );
  OAI22_X1 U2889 ( .A1(n13874), .A2(n13604), .B1(n13600), .B2(n14779), .ZN(
        n8834) );
  OAI22_X1 U2890 ( .A1(n13880), .A2(n13604), .B1(n13600), .B2(n14778), .ZN(
        n8835) );
  OAI22_X1 U2891 ( .A1(n13886), .A2(n13604), .B1(n13600), .B2(n14777), .ZN(
        n8836) );
  OAI22_X1 U2892 ( .A1(n13892), .A2(n13604), .B1(n13600), .B2(n14776), .ZN(
        n8837) );
  OAI22_X1 U2893 ( .A1(n13898), .A2(n13604), .B1(n13601), .B2(n14775), .ZN(
        n8838) );
  OAI22_X1 U2894 ( .A1(n13904), .A2(n13604), .B1(n13601), .B2(n14774), .ZN(
        n8839) );
  OAI22_X1 U2895 ( .A1(n13910), .A2(n13604), .B1(n13601), .B2(n14773), .ZN(
        n8840) );
  OAI22_X1 U2896 ( .A1(n13916), .A2(n13604), .B1(n13601), .B2(n14772), .ZN(
        n8841) );
  OAI22_X1 U2897 ( .A1(n13922), .A2(n13604), .B1(n13601), .B2(n14771), .ZN(
        n8842) );
  OAI22_X1 U2898 ( .A1(n13928), .A2(n13604), .B1(n13601), .B2(n14770), .ZN(
        n8843) );
  OAI22_X1 U2899 ( .A1(n13934), .A2(n13604), .B1(n13601), .B2(n14769), .ZN(
        n8844) );
  OAI22_X1 U2900 ( .A1(n13940), .A2(n13604), .B1(n13601), .B2(n14768), .ZN(
        n8845) );
  OAI22_X1 U2901 ( .A1(n13946), .A2(n13603), .B1(n13601), .B2(n14767), .ZN(
        n8846) );
  OAI22_X1 U2902 ( .A1(n13952), .A2(n13603), .B1(n13601), .B2(n14766), .ZN(
        n8847) );
  OAI22_X1 U2903 ( .A1(n13958), .A2(n13603), .B1(n13601), .B2(n14765), .ZN(
        n8848) );
  OAI22_X1 U2904 ( .A1(n13964), .A2(n13603), .B1(n13601), .B2(n14764), .ZN(
        n8849) );
  OAI22_X1 U2905 ( .A1(n13826), .A2(n13611), .B1(n13606), .B2(n14755), .ZN(
        n8858) );
  OAI22_X1 U2906 ( .A1(n13832), .A2(n13611), .B1(n13606), .B2(n14754), .ZN(
        n8859) );
  OAI22_X1 U2907 ( .A1(n13838), .A2(n13611), .B1(n13606), .B2(n14753), .ZN(
        n8860) );
  OAI22_X1 U2908 ( .A1(n13844), .A2(n13611), .B1(n13606), .B2(n14752), .ZN(
        n8861) );
  OAI22_X1 U2909 ( .A1(n13850), .A2(n13611), .B1(n13606), .B2(n14751), .ZN(
        n8862) );
  OAI22_X1 U2910 ( .A1(n13856), .A2(n13611), .B1(n13606), .B2(n14750), .ZN(
        n8863) );
  OAI22_X1 U2911 ( .A1(n13862), .A2(n13611), .B1(n13606), .B2(n14749), .ZN(
        n8864) );
  OAI22_X1 U2912 ( .A1(n13868), .A2(n13611), .B1(n13606), .B2(n14748), .ZN(
        n8865) );
  OAI22_X1 U2913 ( .A1(n13874), .A2(n13610), .B1(n13606), .B2(n14747), .ZN(
        n8866) );
  OAI22_X1 U2914 ( .A1(n13880), .A2(n13610), .B1(n13606), .B2(n14746), .ZN(
        n8867) );
  OAI22_X1 U2915 ( .A1(n13886), .A2(n13610), .B1(n13606), .B2(n14745), .ZN(
        n8868) );
  OAI22_X1 U2916 ( .A1(n13892), .A2(n13610), .B1(n13606), .B2(n14744), .ZN(
        n8869) );
  OAI22_X1 U2917 ( .A1(n13898), .A2(n13610), .B1(n13607), .B2(n14743), .ZN(
        n8870) );
  OAI22_X1 U2918 ( .A1(n13904), .A2(n13610), .B1(n13607), .B2(n14742), .ZN(
        n8871) );
  OAI22_X1 U2919 ( .A1(n13910), .A2(n13610), .B1(n13607), .B2(n14741), .ZN(
        n8872) );
  OAI22_X1 U2920 ( .A1(n13916), .A2(n13610), .B1(n13607), .B2(n14740), .ZN(
        n8873) );
  OAI22_X1 U2921 ( .A1(n13922), .A2(n13610), .B1(n13607), .B2(n14739), .ZN(
        n8874) );
  OAI22_X1 U2922 ( .A1(n13928), .A2(n13610), .B1(n13607), .B2(n14738), .ZN(
        n8875) );
  OAI22_X1 U2923 ( .A1(n13934), .A2(n13610), .B1(n13607), .B2(n14737), .ZN(
        n8876) );
  OAI22_X1 U2924 ( .A1(n13940), .A2(n13610), .B1(n13607), .B2(n14736), .ZN(
        n8877) );
  OAI22_X1 U2925 ( .A1(n13946), .A2(n13609), .B1(n13607), .B2(n14735), .ZN(
        n8878) );
  OAI22_X1 U2926 ( .A1(n13952), .A2(n13609), .B1(n13607), .B2(n14734), .ZN(
        n8879) );
  OAI22_X1 U2927 ( .A1(n13958), .A2(n13609), .B1(n13607), .B2(n14733), .ZN(
        n8880) );
  OAI22_X1 U2928 ( .A1(n13964), .A2(n13609), .B1(n13607), .B2(n14732), .ZN(
        n8881) );
  OAI22_X1 U2929 ( .A1(n13826), .A2(n13617), .B1(n13612), .B2(n14723), .ZN(
        n8890) );
  OAI22_X1 U2930 ( .A1(n13832), .A2(n13617), .B1(n13612), .B2(n14722), .ZN(
        n8891) );
  OAI22_X1 U2931 ( .A1(n13838), .A2(n13617), .B1(n13612), .B2(n14721), .ZN(
        n8892) );
  OAI22_X1 U2932 ( .A1(n13844), .A2(n13617), .B1(n13612), .B2(n14720), .ZN(
        n8893) );
  OAI22_X1 U2933 ( .A1(n13850), .A2(n13617), .B1(n13612), .B2(n14719), .ZN(
        n8894) );
  OAI22_X1 U2934 ( .A1(n13856), .A2(n13617), .B1(n13612), .B2(n14718), .ZN(
        n8895) );
  OAI22_X1 U2935 ( .A1(n13862), .A2(n13617), .B1(n13612), .B2(n14717), .ZN(
        n8896) );
  OAI22_X1 U2936 ( .A1(n13868), .A2(n13617), .B1(n13612), .B2(n14716), .ZN(
        n8897) );
  OAI22_X1 U2937 ( .A1(n13874), .A2(n13616), .B1(n13612), .B2(n14715), .ZN(
        n8898) );
  OAI22_X1 U2938 ( .A1(n13880), .A2(n13616), .B1(n13612), .B2(n14714), .ZN(
        n8899) );
  OAI22_X1 U2939 ( .A1(n13886), .A2(n13616), .B1(n13612), .B2(n14713), .ZN(
        n8900) );
  OAI22_X1 U2940 ( .A1(n13892), .A2(n13616), .B1(n13612), .B2(n14712), .ZN(
        n8901) );
  OAI22_X1 U2941 ( .A1(n13898), .A2(n13616), .B1(n13613), .B2(n14711), .ZN(
        n8902) );
  OAI22_X1 U2942 ( .A1(n13904), .A2(n13616), .B1(n13613), .B2(n14710), .ZN(
        n8903) );
  OAI22_X1 U2943 ( .A1(n13910), .A2(n13616), .B1(n13613), .B2(n14709), .ZN(
        n8904) );
  OAI22_X1 U2944 ( .A1(n13916), .A2(n13616), .B1(n13613), .B2(n14708), .ZN(
        n8905) );
  OAI22_X1 U2945 ( .A1(n13922), .A2(n13616), .B1(n13613), .B2(n14707), .ZN(
        n8906) );
  OAI22_X1 U2946 ( .A1(n13928), .A2(n13616), .B1(n13613), .B2(n14706), .ZN(
        n8907) );
  OAI22_X1 U2947 ( .A1(n13934), .A2(n13616), .B1(n13613), .B2(n14705), .ZN(
        n8908) );
  OAI22_X1 U2948 ( .A1(n13940), .A2(n13616), .B1(n13613), .B2(n14704), .ZN(
        n8909) );
  OAI22_X1 U2949 ( .A1(n13946), .A2(n13615), .B1(n13613), .B2(n14703), .ZN(
        n8910) );
  OAI22_X1 U2950 ( .A1(n13952), .A2(n13615), .B1(n13613), .B2(n14702), .ZN(
        n8911) );
  OAI22_X1 U2951 ( .A1(n13958), .A2(n13615), .B1(n13613), .B2(n14701), .ZN(
        n8912) );
  OAI22_X1 U2952 ( .A1(n13964), .A2(n13615), .B1(n13613), .B2(n14700), .ZN(
        n8913) );
  OAI22_X1 U2953 ( .A1(n13826), .A2(n13647), .B1(n13642), .B2(n14652), .ZN(
        n9050) );
  OAI22_X1 U2954 ( .A1(n13832), .A2(n13647), .B1(n13642), .B2(n14651), .ZN(
        n9051) );
  OAI22_X1 U2955 ( .A1(n13838), .A2(n13647), .B1(n13642), .B2(n14650), .ZN(
        n9052) );
  OAI22_X1 U2956 ( .A1(n13844), .A2(n13647), .B1(n13642), .B2(n14649), .ZN(
        n9053) );
  OAI22_X1 U2957 ( .A1(n13850), .A2(n13647), .B1(n13642), .B2(n14648), .ZN(
        n9054) );
  OAI22_X1 U2958 ( .A1(n13856), .A2(n13647), .B1(n13642), .B2(n14647), .ZN(
        n9055) );
  OAI22_X1 U2959 ( .A1(n13862), .A2(n13647), .B1(n13642), .B2(n14646), .ZN(
        n9056) );
  OAI22_X1 U2960 ( .A1(n13868), .A2(n13647), .B1(n13642), .B2(n14645), .ZN(
        n9057) );
  OAI22_X1 U2961 ( .A1(n13874), .A2(n13646), .B1(n13642), .B2(n14644), .ZN(
        n9058) );
  OAI22_X1 U2962 ( .A1(n13880), .A2(n13646), .B1(n13642), .B2(n14643), .ZN(
        n9059) );
  OAI22_X1 U2963 ( .A1(n13886), .A2(n13646), .B1(n13642), .B2(n14642), .ZN(
        n9060) );
  OAI22_X1 U2964 ( .A1(n13892), .A2(n13646), .B1(n13642), .B2(n14641), .ZN(
        n9061) );
  OAI22_X1 U2965 ( .A1(n13898), .A2(n13646), .B1(n13643), .B2(n14640), .ZN(
        n9062) );
  OAI22_X1 U2966 ( .A1(n13904), .A2(n13646), .B1(n13643), .B2(n14639), .ZN(
        n9063) );
  OAI22_X1 U2967 ( .A1(n13910), .A2(n13646), .B1(n13643), .B2(n14638), .ZN(
        n9064) );
  OAI22_X1 U2968 ( .A1(n13916), .A2(n13646), .B1(n13643), .B2(n14637), .ZN(
        n9065) );
  OAI22_X1 U2969 ( .A1(n13922), .A2(n13646), .B1(n13643), .B2(n14636), .ZN(
        n9066) );
  OAI22_X1 U2970 ( .A1(n13928), .A2(n13646), .B1(n13643), .B2(n14635), .ZN(
        n9067) );
  OAI22_X1 U2971 ( .A1(n13934), .A2(n13646), .B1(n13643), .B2(n14634), .ZN(
        n9068) );
  OAI22_X1 U2972 ( .A1(n13940), .A2(n13646), .B1(n13643), .B2(n14633), .ZN(
        n9069) );
  OAI22_X1 U2973 ( .A1(n13946), .A2(n13645), .B1(n13643), .B2(n14632), .ZN(
        n9070) );
  OAI22_X1 U2974 ( .A1(n13952), .A2(n13645), .B1(n13643), .B2(n14631), .ZN(
        n9071) );
  OAI22_X1 U2975 ( .A1(n13958), .A2(n13645), .B1(n13643), .B2(n14630), .ZN(
        n9072) );
  OAI22_X1 U2976 ( .A1(n13964), .A2(n13645), .B1(n13643), .B2(n14629), .ZN(
        n9073) );
  OAI22_X1 U2977 ( .A1(n13826), .A2(n13653), .B1(n13648), .B2(n14620), .ZN(
        n9082) );
  OAI22_X1 U2978 ( .A1(n13832), .A2(n13653), .B1(n13648), .B2(n14619), .ZN(
        n9083) );
  OAI22_X1 U2979 ( .A1(n13838), .A2(n13653), .B1(n13648), .B2(n14618), .ZN(
        n9084) );
  OAI22_X1 U2980 ( .A1(n13844), .A2(n13653), .B1(n13648), .B2(n14617), .ZN(
        n9085) );
  OAI22_X1 U2981 ( .A1(n13850), .A2(n13653), .B1(n13648), .B2(n14616), .ZN(
        n9086) );
  OAI22_X1 U2982 ( .A1(n13856), .A2(n13653), .B1(n13648), .B2(n14615), .ZN(
        n9087) );
  OAI22_X1 U2983 ( .A1(n13862), .A2(n13653), .B1(n13648), .B2(n14614), .ZN(
        n9088) );
  OAI22_X1 U2984 ( .A1(n13868), .A2(n13653), .B1(n13648), .B2(n14613), .ZN(
        n9089) );
  OAI22_X1 U2985 ( .A1(n13874), .A2(n13652), .B1(n13648), .B2(n14612), .ZN(
        n9090) );
  OAI22_X1 U2986 ( .A1(n13880), .A2(n13652), .B1(n13648), .B2(n14611), .ZN(
        n9091) );
  OAI22_X1 U2987 ( .A1(n13886), .A2(n13652), .B1(n13648), .B2(n14610), .ZN(
        n9092) );
  OAI22_X1 U2988 ( .A1(n13892), .A2(n13652), .B1(n13648), .B2(n14609), .ZN(
        n9093) );
  OAI22_X1 U2989 ( .A1(n13898), .A2(n13652), .B1(n13649), .B2(n14608), .ZN(
        n9094) );
  OAI22_X1 U2990 ( .A1(n13904), .A2(n13652), .B1(n13649), .B2(n14607), .ZN(
        n9095) );
  OAI22_X1 U2991 ( .A1(n13910), .A2(n13652), .B1(n13649), .B2(n14606), .ZN(
        n9096) );
  OAI22_X1 U2992 ( .A1(n13916), .A2(n13652), .B1(n13649), .B2(n14605), .ZN(
        n9097) );
  OAI22_X1 U2993 ( .A1(n13922), .A2(n13652), .B1(n13649), .B2(n14604), .ZN(
        n9098) );
  OAI22_X1 U2994 ( .A1(n13928), .A2(n13652), .B1(n13649), .B2(n14603), .ZN(
        n9099) );
  OAI22_X1 U2995 ( .A1(n13934), .A2(n13652), .B1(n13649), .B2(n14602), .ZN(
        n9100) );
  OAI22_X1 U2996 ( .A1(n13940), .A2(n13652), .B1(n13649), .B2(n14601), .ZN(
        n9101) );
  OAI22_X1 U2997 ( .A1(n13946), .A2(n13651), .B1(n13649), .B2(n14600), .ZN(
        n9102) );
  OAI22_X1 U2998 ( .A1(n13952), .A2(n13651), .B1(n13649), .B2(n14599), .ZN(
        n9103) );
  OAI22_X1 U2999 ( .A1(n13958), .A2(n13651), .B1(n13649), .B2(n14598), .ZN(
        n9104) );
  OAI22_X1 U3000 ( .A1(n13964), .A2(n13651), .B1(n13649), .B2(n14597), .ZN(
        n9105) );
  OAI22_X1 U3001 ( .A1(n13826), .A2(n13659), .B1(n13654), .B2(n14588), .ZN(
        n9114) );
  OAI22_X1 U3002 ( .A1(n13832), .A2(n13659), .B1(n13654), .B2(n14587), .ZN(
        n9115) );
  OAI22_X1 U3003 ( .A1(n13838), .A2(n13659), .B1(n13654), .B2(n14586), .ZN(
        n9116) );
  OAI22_X1 U3004 ( .A1(n13844), .A2(n13659), .B1(n13654), .B2(n14585), .ZN(
        n9117) );
  OAI22_X1 U3005 ( .A1(n13850), .A2(n13659), .B1(n13654), .B2(n14584), .ZN(
        n9118) );
  OAI22_X1 U3006 ( .A1(n13856), .A2(n13659), .B1(n13654), .B2(n14583), .ZN(
        n9119) );
  OAI22_X1 U3007 ( .A1(n13862), .A2(n13659), .B1(n13654), .B2(n14582), .ZN(
        n9120) );
  OAI22_X1 U3008 ( .A1(n13868), .A2(n13659), .B1(n13654), .B2(n14581), .ZN(
        n9121) );
  OAI22_X1 U3009 ( .A1(n13874), .A2(n13658), .B1(n13654), .B2(n14580), .ZN(
        n9122) );
  OAI22_X1 U3010 ( .A1(n13880), .A2(n13658), .B1(n13654), .B2(n14579), .ZN(
        n9123) );
  OAI22_X1 U3011 ( .A1(n13886), .A2(n13658), .B1(n13654), .B2(n14578), .ZN(
        n9124) );
  OAI22_X1 U3012 ( .A1(n13892), .A2(n13658), .B1(n13654), .B2(n14577), .ZN(
        n9125) );
  OAI22_X1 U3013 ( .A1(n13898), .A2(n13658), .B1(n13655), .B2(n14576), .ZN(
        n9126) );
  OAI22_X1 U3014 ( .A1(n13904), .A2(n13658), .B1(n13655), .B2(n14575), .ZN(
        n9127) );
  OAI22_X1 U3015 ( .A1(n13910), .A2(n13658), .B1(n13655), .B2(n14574), .ZN(
        n9128) );
  OAI22_X1 U3016 ( .A1(n13916), .A2(n13658), .B1(n13655), .B2(n14573), .ZN(
        n9129) );
  OAI22_X1 U3017 ( .A1(n13922), .A2(n13658), .B1(n13655), .B2(n14572), .ZN(
        n9130) );
  OAI22_X1 U3018 ( .A1(n13928), .A2(n13658), .B1(n13655), .B2(n14571), .ZN(
        n9131) );
  OAI22_X1 U3019 ( .A1(n13934), .A2(n13658), .B1(n13655), .B2(n14570), .ZN(
        n9132) );
  OAI22_X1 U3020 ( .A1(n13940), .A2(n13658), .B1(n13655), .B2(n14569), .ZN(
        n9133) );
  OAI22_X1 U3021 ( .A1(n13946), .A2(n13657), .B1(n13655), .B2(n14568), .ZN(
        n9134) );
  OAI22_X1 U3022 ( .A1(n13952), .A2(n13657), .B1(n13655), .B2(n14567), .ZN(
        n9135) );
  OAI22_X1 U3023 ( .A1(n13958), .A2(n13657), .B1(n13655), .B2(n14566), .ZN(
        n9136) );
  OAI22_X1 U3024 ( .A1(n13964), .A2(n13657), .B1(n13655), .B2(n14565), .ZN(
        n9137) );
  OAI22_X1 U3025 ( .A1(n13825), .A2(n13665), .B1(n13660), .B2(n14556), .ZN(
        n9146) );
  OAI22_X1 U3026 ( .A1(n13832), .A2(n13665), .B1(n13660), .B2(n14555), .ZN(
        n9147) );
  OAI22_X1 U3027 ( .A1(n13838), .A2(n13665), .B1(n13660), .B2(n14554), .ZN(
        n9148) );
  OAI22_X1 U3028 ( .A1(n13844), .A2(n13665), .B1(n13660), .B2(n14553), .ZN(
        n9149) );
  OAI22_X1 U3029 ( .A1(n13850), .A2(n13665), .B1(n13660), .B2(n14552), .ZN(
        n9150) );
  OAI22_X1 U3030 ( .A1(n13856), .A2(n13665), .B1(n13660), .B2(n14551), .ZN(
        n9151) );
  OAI22_X1 U3031 ( .A1(n13862), .A2(n13665), .B1(n13660), .B2(n14550), .ZN(
        n9152) );
  OAI22_X1 U3032 ( .A1(n13868), .A2(n13665), .B1(n13660), .B2(n14549), .ZN(
        n9153) );
  OAI22_X1 U3033 ( .A1(n13874), .A2(n13664), .B1(n13660), .B2(n14548), .ZN(
        n9154) );
  OAI22_X1 U3034 ( .A1(n13880), .A2(n13664), .B1(n13660), .B2(n14547), .ZN(
        n9155) );
  OAI22_X1 U3035 ( .A1(n13886), .A2(n13664), .B1(n13660), .B2(n14546), .ZN(
        n9156) );
  OAI22_X1 U3036 ( .A1(n13892), .A2(n13664), .B1(n13660), .B2(n14545), .ZN(
        n9157) );
  OAI22_X1 U3037 ( .A1(n13898), .A2(n13664), .B1(n13661), .B2(n14544), .ZN(
        n9158) );
  OAI22_X1 U3038 ( .A1(n13904), .A2(n13664), .B1(n13661), .B2(n14543), .ZN(
        n9159) );
  OAI22_X1 U3039 ( .A1(n13910), .A2(n13664), .B1(n13661), .B2(n14542), .ZN(
        n9160) );
  OAI22_X1 U3040 ( .A1(n13916), .A2(n13664), .B1(n13661), .B2(n14541), .ZN(
        n9161) );
  OAI22_X1 U3041 ( .A1(n13922), .A2(n13664), .B1(n13661), .B2(n14540), .ZN(
        n9162) );
  OAI22_X1 U3042 ( .A1(n13928), .A2(n13664), .B1(n13661), .B2(n14539), .ZN(
        n9163) );
  OAI22_X1 U3043 ( .A1(n13934), .A2(n13664), .B1(n13661), .B2(n14538), .ZN(
        n9164) );
  OAI22_X1 U3044 ( .A1(n13940), .A2(n13664), .B1(n13661), .B2(n14537), .ZN(
        n9165) );
  OAI22_X1 U3045 ( .A1(n13946), .A2(n13663), .B1(n13661), .B2(n14536), .ZN(
        n9166) );
  OAI22_X1 U3046 ( .A1(n13952), .A2(n13663), .B1(n13661), .B2(n14535), .ZN(
        n9167) );
  OAI22_X1 U3047 ( .A1(n13958), .A2(n13663), .B1(n13661), .B2(n14534), .ZN(
        n9168) );
  OAI22_X1 U3048 ( .A1(n13964), .A2(n13663), .B1(n13661), .B2(n14533), .ZN(
        n9169) );
  OAI22_X1 U3049 ( .A1(n13825), .A2(n13671), .B1(n13666), .B2(n14524), .ZN(
        n9178) );
  OAI22_X1 U3050 ( .A1(n13831), .A2(n13671), .B1(n13666), .B2(n14523), .ZN(
        n9179) );
  OAI22_X1 U3051 ( .A1(n13837), .A2(n13671), .B1(n13666), .B2(n14522), .ZN(
        n9180) );
  OAI22_X1 U3052 ( .A1(n13843), .A2(n13671), .B1(n13666), .B2(n14521), .ZN(
        n9181) );
  OAI22_X1 U3053 ( .A1(n13849), .A2(n13671), .B1(n13666), .B2(n14520), .ZN(
        n9182) );
  OAI22_X1 U3054 ( .A1(n13855), .A2(n13671), .B1(n13666), .B2(n14519), .ZN(
        n9183) );
  OAI22_X1 U3055 ( .A1(n13861), .A2(n13671), .B1(n13666), .B2(n14518), .ZN(
        n9184) );
  OAI22_X1 U3056 ( .A1(n13867), .A2(n13671), .B1(n13666), .B2(n14517), .ZN(
        n9185) );
  OAI22_X1 U3057 ( .A1(n13873), .A2(n13670), .B1(n13666), .B2(n14516), .ZN(
        n9186) );
  OAI22_X1 U3058 ( .A1(n13879), .A2(n13670), .B1(n13666), .B2(n14515), .ZN(
        n9187) );
  OAI22_X1 U3059 ( .A1(n13885), .A2(n13670), .B1(n13666), .B2(n14514), .ZN(
        n9188) );
  OAI22_X1 U3060 ( .A1(n13891), .A2(n13670), .B1(n13666), .B2(n14513), .ZN(
        n9189) );
  OAI22_X1 U3061 ( .A1(n13897), .A2(n13670), .B1(n13667), .B2(n14512), .ZN(
        n9190) );
  OAI22_X1 U3062 ( .A1(n13903), .A2(n13670), .B1(n13667), .B2(n14511), .ZN(
        n9191) );
  OAI22_X1 U3063 ( .A1(n13909), .A2(n13670), .B1(n13667), .B2(n14510), .ZN(
        n9192) );
  OAI22_X1 U3064 ( .A1(n13915), .A2(n13670), .B1(n13667), .B2(n14509), .ZN(
        n9193) );
  OAI22_X1 U3065 ( .A1(n13921), .A2(n13670), .B1(n13667), .B2(n14508), .ZN(
        n9194) );
  OAI22_X1 U3066 ( .A1(n13927), .A2(n13670), .B1(n13667), .B2(n14507), .ZN(
        n9195) );
  OAI22_X1 U3067 ( .A1(n13933), .A2(n13670), .B1(n13667), .B2(n14506), .ZN(
        n9196) );
  OAI22_X1 U3068 ( .A1(n13939), .A2(n13670), .B1(n13667), .B2(n14505), .ZN(
        n9197) );
  OAI22_X1 U3069 ( .A1(n13945), .A2(n13669), .B1(n13667), .B2(n14504), .ZN(
        n9198) );
  OAI22_X1 U3070 ( .A1(n13951), .A2(n13669), .B1(n13667), .B2(n14503), .ZN(
        n9199) );
  OAI22_X1 U3071 ( .A1(n13957), .A2(n13669), .B1(n13667), .B2(n14502), .ZN(
        n9200) );
  OAI22_X1 U3072 ( .A1(n13963), .A2(n13669), .B1(n13667), .B2(n14501), .ZN(
        n9201) );
  OAI22_X1 U3073 ( .A1(n13825), .A2(n13701), .B1(n13696), .B2(n14439), .ZN(
        n9338) );
  OAI22_X1 U3074 ( .A1(n13831), .A2(n13701), .B1(n13696), .B2(n14438), .ZN(
        n9339) );
  OAI22_X1 U3075 ( .A1(n13837), .A2(n13701), .B1(n13696), .B2(n14437), .ZN(
        n9340) );
  OAI22_X1 U3076 ( .A1(n13843), .A2(n13701), .B1(n13696), .B2(n14436), .ZN(
        n9341) );
  OAI22_X1 U3077 ( .A1(n13849), .A2(n13701), .B1(n13696), .B2(n14435), .ZN(
        n9342) );
  OAI22_X1 U3078 ( .A1(n13855), .A2(n13701), .B1(n13696), .B2(n14434), .ZN(
        n9343) );
  OAI22_X1 U3079 ( .A1(n13861), .A2(n13701), .B1(n13696), .B2(n14433), .ZN(
        n9344) );
  OAI22_X1 U3080 ( .A1(n13867), .A2(n13701), .B1(n13696), .B2(n14432), .ZN(
        n9345) );
  OAI22_X1 U3081 ( .A1(n13873), .A2(n13700), .B1(n13696), .B2(n14431), .ZN(
        n9346) );
  OAI22_X1 U3082 ( .A1(n13879), .A2(n13700), .B1(n13696), .B2(n14430), .ZN(
        n9347) );
  OAI22_X1 U3083 ( .A1(n13885), .A2(n13700), .B1(n13696), .B2(n14429), .ZN(
        n9348) );
  OAI22_X1 U3084 ( .A1(n13891), .A2(n13700), .B1(n13696), .B2(n14428), .ZN(
        n9349) );
  OAI22_X1 U3085 ( .A1(n13897), .A2(n13700), .B1(n13697), .B2(n14427), .ZN(
        n9350) );
  OAI22_X1 U3086 ( .A1(n13903), .A2(n13700), .B1(n13697), .B2(n14426), .ZN(
        n9351) );
  OAI22_X1 U3087 ( .A1(n13909), .A2(n13700), .B1(n13697), .B2(n14425), .ZN(
        n9352) );
  OAI22_X1 U3088 ( .A1(n13915), .A2(n13700), .B1(n13697), .B2(n14424), .ZN(
        n9353) );
  OAI22_X1 U3089 ( .A1(n13921), .A2(n13700), .B1(n13697), .B2(n14423), .ZN(
        n9354) );
  OAI22_X1 U3090 ( .A1(n13927), .A2(n13700), .B1(n13697), .B2(n14422), .ZN(
        n9355) );
  OAI22_X1 U3091 ( .A1(n13933), .A2(n13700), .B1(n13697), .B2(n14421), .ZN(
        n9356) );
  OAI22_X1 U3092 ( .A1(n13939), .A2(n13700), .B1(n13697), .B2(n14420), .ZN(
        n9357) );
  OAI22_X1 U3093 ( .A1(n13945), .A2(n13699), .B1(n13697), .B2(n14419), .ZN(
        n9358) );
  OAI22_X1 U3094 ( .A1(n13951), .A2(n13699), .B1(n13697), .B2(n14418), .ZN(
        n9359) );
  OAI22_X1 U3095 ( .A1(n13957), .A2(n13699), .B1(n13697), .B2(n14417), .ZN(
        n9360) );
  OAI22_X1 U3096 ( .A1(n13963), .A2(n13699), .B1(n13697), .B2(n14416), .ZN(
        n9361) );
  OAI22_X1 U3097 ( .A1(n13825), .A2(n13707), .B1(n13702), .B2(n14407), .ZN(
        n9370) );
  OAI22_X1 U3098 ( .A1(n13832), .A2(n13707), .B1(n13702), .B2(n14406), .ZN(
        n9371) );
  OAI22_X1 U3099 ( .A1(n13838), .A2(n13707), .B1(n13702), .B2(n14405), .ZN(
        n9372) );
  OAI22_X1 U3100 ( .A1(n13844), .A2(n13707), .B1(n13702), .B2(n14404), .ZN(
        n9373) );
  OAI22_X1 U3101 ( .A1(n13850), .A2(n13707), .B1(n13702), .B2(n14403), .ZN(
        n9374) );
  OAI22_X1 U3102 ( .A1(n13856), .A2(n13707), .B1(n13702), .B2(n14402), .ZN(
        n9375) );
  OAI22_X1 U3103 ( .A1(n13862), .A2(n13707), .B1(n13702), .B2(n14401), .ZN(
        n9376) );
  OAI22_X1 U3104 ( .A1(n13868), .A2(n13707), .B1(n13702), .B2(n14400), .ZN(
        n9377) );
  OAI22_X1 U3105 ( .A1(n13874), .A2(n13706), .B1(n13702), .B2(n14399), .ZN(
        n9378) );
  OAI22_X1 U3106 ( .A1(n13880), .A2(n13706), .B1(n13702), .B2(n14398), .ZN(
        n9379) );
  OAI22_X1 U3107 ( .A1(n13886), .A2(n13706), .B1(n13702), .B2(n14397), .ZN(
        n9380) );
  OAI22_X1 U3108 ( .A1(n13892), .A2(n13706), .B1(n13702), .B2(n14396), .ZN(
        n9381) );
  OAI22_X1 U3109 ( .A1(n13898), .A2(n13706), .B1(n13703), .B2(n14395), .ZN(
        n9382) );
  OAI22_X1 U3110 ( .A1(n13904), .A2(n13706), .B1(n13703), .B2(n14394), .ZN(
        n9383) );
  OAI22_X1 U3111 ( .A1(n13910), .A2(n13706), .B1(n13703), .B2(n14393), .ZN(
        n9384) );
  OAI22_X1 U3112 ( .A1(n13916), .A2(n13706), .B1(n13703), .B2(n14392), .ZN(
        n9385) );
  OAI22_X1 U3113 ( .A1(n13922), .A2(n13706), .B1(n13703), .B2(n14391), .ZN(
        n9386) );
  OAI22_X1 U3114 ( .A1(n13928), .A2(n13706), .B1(n13703), .B2(n14390), .ZN(
        n9387) );
  OAI22_X1 U3115 ( .A1(n13934), .A2(n13706), .B1(n13703), .B2(n14389), .ZN(
        n9388) );
  OAI22_X1 U3116 ( .A1(n13940), .A2(n13706), .B1(n13703), .B2(n14388), .ZN(
        n9389) );
  OAI22_X1 U3117 ( .A1(n13946), .A2(n13705), .B1(n13703), .B2(n14387), .ZN(
        n9390) );
  OAI22_X1 U3118 ( .A1(n13952), .A2(n13705), .B1(n13703), .B2(n14386), .ZN(
        n9391) );
  OAI22_X1 U3119 ( .A1(n13958), .A2(n13705), .B1(n13703), .B2(n14385), .ZN(
        n9392) );
  OAI22_X1 U3120 ( .A1(n13964), .A2(n13705), .B1(n13703), .B2(n14384), .ZN(
        n9393) );
  OAI22_X1 U3121 ( .A1(n13825), .A2(n13713), .B1(n13708), .B2(n14375), .ZN(
        n9402) );
  OAI22_X1 U3122 ( .A1(n13831), .A2(n13713), .B1(n13708), .B2(n14374), .ZN(
        n9403) );
  OAI22_X1 U3123 ( .A1(n13837), .A2(n13713), .B1(n13708), .B2(n14373), .ZN(
        n9404) );
  OAI22_X1 U3124 ( .A1(n13843), .A2(n13713), .B1(n13708), .B2(n14372), .ZN(
        n9405) );
  OAI22_X1 U3125 ( .A1(n13849), .A2(n13713), .B1(n13708), .B2(n14371), .ZN(
        n9406) );
  OAI22_X1 U3126 ( .A1(n13855), .A2(n13713), .B1(n13708), .B2(n14370), .ZN(
        n9407) );
  OAI22_X1 U3127 ( .A1(n13861), .A2(n13713), .B1(n13708), .B2(n14369), .ZN(
        n9408) );
  OAI22_X1 U3128 ( .A1(n13867), .A2(n13713), .B1(n13708), .B2(n14368), .ZN(
        n9409) );
  OAI22_X1 U3129 ( .A1(n13873), .A2(n13712), .B1(n13708), .B2(n14367), .ZN(
        n9410) );
  OAI22_X1 U3130 ( .A1(n13879), .A2(n13712), .B1(n13708), .B2(n14366), .ZN(
        n9411) );
  OAI22_X1 U3131 ( .A1(n13885), .A2(n13712), .B1(n13708), .B2(n14365), .ZN(
        n9412) );
  OAI22_X1 U3132 ( .A1(n13891), .A2(n13712), .B1(n13708), .B2(n14364), .ZN(
        n9413) );
  OAI22_X1 U3133 ( .A1(n13897), .A2(n13712), .B1(n13709), .B2(n14363), .ZN(
        n9414) );
  OAI22_X1 U3134 ( .A1(n13903), .A2(n13712), .B1(n13709), .B2(n14362), .ZN(
        n9415) );
  OAI22_X1 U3135 ( .A1(n13909), .A2(n13712), .B1(n13709), .B2(n14361), .ZN(
        n9416) );
  OAI22_X1 U3136 ( .A1(n13915), .A2(n13712), .B1(n13709), .B2(n14360), .ZN(
        n9417) );
  OAI22_X1 U3137 ( .A1(n13921), .A2(n13712), .B1(n13709), .B2(n14359), .ZN(
        n9418) );
  OAI22_X1 U3138 ( .A1(n13927), .A2(n13712), .B1(n13709), .B2(n14358), .ZN(
        n9419) );
  OAI22_X1 U3139 ( .A1(n13933), .A2(n13712), .B1(n13709), .B2(n14357), .ZN(
        n9420) );
  OAI22_X1 U3140 ( .A1(n13939), .A2(n13712), .B1(n13709), .B2(n14356), .ZN(
        n9421) );
  OAI22_X1 U3141 ( .A1(n13945), .A2(n13711), .B1(n13709), .B2(n14355), .ZN(
        n9422) );
  OAI22_X1 U3142 ( .A1(n13951), .A2(n13711), .B1(n13709), .B2(n14354), .ZN(
        n9423) );
  OAI22_X1 U3143 ( .A1(n13957), .A2(n13711), .B1(n13709), .B2(n14353), .ZN(
        n9424) );
  OAI22_X1 U3144 ( .A1(n13963), .A2(n13711), .B1(n13709), .B2(n14352), .ZN(
        n9425) );
  OAI22_X1 U3145 ( .A1(n13825), .A2(n13719), .B1(n13714), .B2(n14343), .ZN(
        n9434) );
  OAI22_X1 U3146 ( .A1(n13831), .A2(n13719), .B1(n13714), .B2(n14342), .ZN(
        n9435) );
  OAI22_X1 U3147 ( .A1(n13837), .A2(n13719), .B1(n13714), .B2(n14341), .ZN(
        n9436) );
  OAI22_X1 U3148 ( .A1(n13843), .A2(n13719), .B1(n13714), .B2(n14340), .ZN(
        n9437) );
  OAI22_X1 U3149 ( .A1(n13849), .A2(n13719), .B1(n13714), .B2(n14339), .ZN(
        n9438) );
  OAI22_X1 U3150 ( .A1(n13855), .A2(n13719), .B1(n13714), .B2(n14338), .ZN(
        n9439) );
  OAI22_X1 U3151 ( .A1(n13861), .A2(n13719), .B1(n13714), .B2(n14337), .ZN(
        n9440) );
  OAI22_X1 U3152 ( .A1(n13867), .A2(n13719), .B1(n13714), .B2(n14336), .ZN(
        n9441) );
  OAI22_X1 U3153 ( .A1(n13873), .A2(n13718), .B1(n13714), .B2(n14335), .ZN(
        n9442) );
  OAI22_X1 U3154 ( .A1(n13879), .A2(n13718), .B1(n13714), .B2(n14334), .ZN(
        n9443) );
  OAI22_X1 U3155 ( .A1(n13885), .A2(n13718), .B1(n13714), .B2(n14333), .ZN(
        n9444) );
  OAI22_X1 U3156 ( .A1(n13891), .A2(n13718), .B1(n13714), .B2(n14332), .ZN(
        n9445) );
  OAI22_X1 U3157 ( .A1(n13897), .A2(n13718), .B1(n13715), .B2(n14331), .ZN(
        n9446) );
  OAI22_X1 U3158 ( .A1(n13903), .A2(n13718), .B1(n13715), .B2(n14330), .ZN(
        n9447) );
  OAI22_X1 U3159 ( .A1(n13909), .A2(n13718), .B1(n13715), .B2(n14329), .ZN(
        n9448) );
  OAI22_X1 U3160 ( .A1(n13915), .A2(n13718), .B1(n13715), .B2(n14328), .ZN(
        n9449) );
  OAI22_X1 U3161 ( .A1(n13921), .A2(n13718), .B1(n13715), .B2(n14327), .ZN(
        n9450) );
  OAI22_X1 U3162 ( .A1(n13927), .A2(n13718), .B1(n13715), .B2(n14326), .ZN(
        n9451) );
  OAI22_X1 U3163 ( .A1(n13933), .A2(n13718), .B1(n13715), .B2(n14325), .ZN(
        n9452) );
  OAI22_X1 U3164 ( .A1(n13939), .A2(n13718), .B1(n13715), .B2(n14324), .ZN(
        n9453) );
  OAI22_X1 U3165 ( .A1(n13945), .A2(n13717), .B1(n13715), .B2(n14323), .ZN(
        n9454) );
  OAI22_X1 U3166 ( .A1(n13951), .A2(n13717), .B1(n13715), .B2(n14322), .ZN(
        n9455) );
  OAI22_X1 U3167 ( .A1(n13957), .A2(n13717), .B1(n13715), .B2(n14321), .ZN(
        n9456) );
  OAI22_X1 U3168 ( .A1(n13963), .A2(n13717), .B1(n13715), .B2(n14320), .ZN(
        n9457) );
  OAI22_X1 U3169 ( .A1(n13825), .A2(n13725), .B1(n13720), .B2(n14311), .ZN(
        n9466) );
  OAI22_X1 U3170 ( .A1(n13831), .A2(n13725), .B1(n13720), .B2(n14310), .ZN(
        n9467) );
  OAI22_X1 U3171 ( .A1(n13837), .A2(n13725), .B1(n13720), .B2(n14309), .ZN(
        n9468) );
  OAI22_X1 U3172 ( .A1(n13843), .A2(n13725), .B1(n13720), .B2(n14308), .ZN(
        n9469) );
  OAI22_X1 U3173 ( .A1(n13849), .A2(n13725), .B1(n13720), .B2(n14307), .ZN(
        n9470) );
  OAI22_X1 U3174 ( .A1(n13855), .A2(n13725), .B1(n13720), .B2(n14306), .ZN(
        n9471) );
  OAI22_X1 U3175 ( .A1(n13861), .A2(n13725), .B1(n13720), .B2(n14305), .ZN(
        n9472) );
  OAI22_X1 U3176 ( .A1(n13867), .A2(n13725), .B1(n13720), .B2(n14304), .ZN(
        n9473) );
  OAI22_X1 U3177 ( .A1(n13873), .A2(n13724), .B1(n13720), .B2(n14303), .ZN(
        n9474) );
  OAI22_X1 U3178 ( .A1(n13879), .A2(n13724), .B1(n13720), .B2(n14302), .ZN(
        n9475) );
  OAI22_X1 U3179 ( .A1(n13885), .A2(n13724), .B1(n13720), .B2(n14301), .ZN(
        n9476) );
  OAI22_X1 U3180 ( .A1(n13891), .A2(n13724), .B1(n13720), .B2(n14300), .ZN(
        n9477) );
  OAI22_X1 U3181 ( .A1(n13897), .A2(n13724), .B1(n13721), .B2(n14299), .ZN(
        n9478) );
  OAI22_X1 U3182 ( .A1(n13903), .A2(n13724), .B1(n13721), .B2(n14298), .ZN(
        n9479) );
  OAI22_X1 U3183 ( .A1(n13909), .A2(n13724), .B1(n13721), .B2(n14297), .ZN(
        n9480) );
  OAI22_X1 U3184 ( .A1(n13915), .A2(n13724), .B1(n13721), .B2(n14296), .ZN(
        n9481) );
  OAI22_X1 U3185 ( .A1(n13921), .A2(n13724), .B1(n13721), .B2(n14295), .ZN(
        n9482) );
  OAI22_X1 U3186 ( .A1(n13927), .A2(n13724), .B1(n13721), .B2(n14294), .ZN(
        n9483) );
  OAI22_X1 U3187 ( .A1(n13933), .A2(n13724), .B1(n13721), .B2(n14293), .ZN(
        n9484) );
  OAI22_X1 U3188 ( .A1(n13939), .A2(n13724), .B1(n13721), .B2(n14292), .ZN(
        n9485) );
  OAI22_X1 U3189 ( .A1(n13945), .A2(n13723), .B1(n13721), .B2(n14291), .ZN(
        n9486) );
  OAI22_X1 U3190 ( .A1(n13951), .A2(n13723), .B1(n13721), .B2(n14290), .ZN(
        n9487) );
  OAI22_X1 U3191 ( .A1(n13957), .A2(n13723), .B1(n13721), .B2(n14289), .ZN(
        n9488) );
  OAI22_X1 U3192 ( .A1(n13963), .A2(n13723), .B1(n13721), .B2(n14288), .ZN(
        n9489) );
  OAI22_X1 U3193 ( .A1(n13824), .A2(n13749), .B1(n13744), .B2(n12661), .ZN(
        n9594) );
  OAI22_X1 U3194 ( .A1(n13830), .A2(n13749), .B1(n13744), .B2(n12663), .ZN(
        n9595) );
  OAI22_X1 U3195 ( .A1(n13836), .A2(n13749), .B1(n13744), .B2(n12665), .ZN(
        n9596) );
  OAI22_X1 U3196 ( .A1(n13842), .A2(n13749), .B1(n13744), .B2(n12667), .ZN(
        n9597) );
  OAI22_X1 U3197 ( .A1(n13848), .A2(n13749), .B1(n13744), .B2(n12669), .ZN(
        n9598) );
  OAI22_X1 U3198 ( .A1(n13854), .A2(n13749), .B1(n13744), .B2(n12671), .ZN(
        n9599) );
  OAI22_X1 U3199 ( .A1(n13860), .A2(n13749), .B1(n13744), .B2(n12673), .ZN(
        n9600) );
  OAI22_X1 U3200 ( .A1(n13866), .A2(n13749), .B1(n13744), .B2(n12675), .ZN(
        n9601) );
  OAI22_X1 U3201 ( .A1(n13872), .A2(n13748), .B1(n13744), .B2(n12677), .ZN(
        n9602) );
  OAI22_X1 U3202 ( .A1(n13878), .A2(n13748), .B1(n13744), .B2(n12679), .ZN(
        n9603) );
  OAI22_X1 U3203 ( .A1(n13884), .A2(n13748), .B1(n13744), .B2(n12681), .ZN(
        n9604) );
  OAI22_X1 U3204 ( .A1(n13890), .A2(n13748), .B1(n13744), .B2(n12683), .ZN(
        n9605) );
  OAI22_X1 U3205 ( .A1(n13896), .A2(n13748), .B1(n13745), .B2(n12685), .ZN(
        n9606) );
  OAI22_X1 U3206 ( .A1(n13902), .A2(n13748), .B1(n13745), .B2(n12687), .ZN(
        n9607) );
  OAI22_X1 U3207 ( .A1(n13908), .A2(n13748), .B1(n13745), .B2(n12689), .ZN(
        n9608) );
  OAI22_X1 U3208 ( .A1(n13914), .A2(n13748), .B1(n13745), .B2(n12691), .ZN(
        n9609) );
  OAI22_X1 U3209 ( .A1(n13920), .A2(n13748), .B1(n13745), .B2(n12693), .ZN(
        n9610) );
  OAI22_X1 U3210 ( .A1(n13926), .A2(n13748), .B1(n13745), .B2(n12695), .ZN(
        n9611) );
  OAI22_X1 U3211 ( .A1(n13932), .A2(n13748), .B1(n13745), .B2(n12697), .ZN(
        n9612) );
  OAI22_X1 U3212 ( .A1(n13938), .A2(n13748), .B1(n13745), .B2(n12699), .ZN(
        n9613) );
  OAI22_X1 U3213 ( .A1(n13944), .A2(n13747), .B1(n13745), .B2(n12701), .ZN(
        n9614) );
  OAI22_X1 U3214 ( .A1(n13950), .A2(n13747), .B1(n13745), .B2(n12703), .ZN(
        n9615) );
  OAI22_X1 U3215 ( .A1(n13956), .A2(n13747), .B1(n13745), .B2(n12705), .ZN(
        n9616) );
  OAI22_X1 U3216 ( .A1(n13962), .A2(n13747), .B1(n13745), .B2(n12707), .ZN(
        n9617) );
  OAI22_X1 U3217 ( .A1(n13824), .A2(n13767), .B1(n13762), .B2(n14203), .ZN(
        n9690) );
  OAI22_X1 U3218 ( .A1(n13830), .A2(n13767), .B1(n13762), .B2(n14202), .ZN(
        n9691) );
  OAI22_X1 U3219 ( .A1(n13836), .A2(n13767), .B1(n13762), .B2(n14201), .ZN(
        n9692) );
  OAI22_X1 U3220 ( .A1(n13842), .A2(n13767), .B1(n13762), .B2(n14200), .ZN(
        n9693) );
  OAI22_X1 U3221 ( .A1(n13848), .A2(n13767), .B1(n13762), .B2(n14199), .ZN(
        n9694) );
  OAI22_X1 U3222 ( .A1(n13854), .A2(n13767), .B1(n13762), .B2(n14198), .ZN(
        n9695) );
  OAI22_X1 U3223 ( .A1(n13860), .A2(n13767), .B1(n13762), .B2(n14197), .ZN(
        n9696) );
  OAI22_X1 U3224 ( .A1(n13866), .A2(n13767), .B1(n13762), .B2(n14196), .ZN(
        n9697) );
  OAI22_X1 U3225 ( .A1(n13872), .A2(n13766), .B1(n13762), .B2(n14195), .ZN(
        n9698) );
  OAI22_X1 U3226 ( .A1(n13878), .A2(n13766), .B1(n13762), .B2(n14194), .ZN(
        n9699) );
  OAI22_X1 U3227 ( .A1(n13884), .A2(n13766), .B1(n13762), .B2(n14193), .ZN(
        n9700) );
  OAI22_X1 U3228 ( .A1(n13890), .A2(n13766), .B1(n13762), .B2(n14192), .ZN(
        n9701) );
  OAI22_X1 U3229 ( .A1(n13896), .A2(n13766), .B1(n13763), .B2(n14191), .ZN(
        n9702) );
  OAI22_X1 U3230 ( .A1(n13902), .A2(n13766), .B1(n13763), .B2(n14190), .ZN(
        n9703) );
  OAI22_X1 U3231 ( .A1(n13908), .A2(n13766), .B1(n13763), .B2(n14189), .ZN(
        n9704) );
  OAI22_X1 U3232 ( .A1(n13914), .A2(n13766), .B1(n13763), .B2(n14188), .ZN(
        n9705) );
  OAI22_X1 U3233 ( .A1(n13920), .A2(n13766), .B1(n13763), .B2(n14187), .ZN(
        n9706) );
  OAI22_X1 U3234 ( .A1(n13926), .A2(n13766), .B1(n13763), .B2(n14186), .ZN(
        n9707) );
  OAI22_X1 U3235 ( .A1(n13932), .A2(n13766), .B1(n13763), .B2(n14185), .ZN(
        n9708) );
  OAI22_X1 U3236 ( .A1(n13938), .A2(n13766), .B1(n13763), .B2(n14184), .ZN(
        n9709) );
  OAI22_X1 U3237 ( .A1(n13944), .A2(n13765), .B1(n13763), .B2(n14183), .ZN(
        n9710) );
  OAI22_X1 U3238 ( .A1(n13950), .A2(n13765), .B1(n13763), .B2(n14182), .ZN(
        n9711) );
  OAI22_X1 U3239 ( .A1(n13956), .A2(n13765), .B1(n13763), .B2(n14181), .ZN(
        n9712) );
  OAI22_X1 U3240 ( .A1(n13962), .A2(n13765), .B1(n13763), .B2(n14180), .ZN(
        n9713) );
  OAI22_X1 U3241 ( .A1(n13824), .A2(n13773), .B1(n13768), .B2(n14171), .ZN(
        n9722) );
  OAI22_X1 U3242 ( .A1(n13830), .A2(n13773), .B1(n13768), .B2(n14170), .ZN(
        n9723) );
  OAI22_X1 U3243 ( .A1(n13836), .A2(n13773), .B1(n13768), .B2(n14169), .ZN(
        n9724) );
  OAI22_X1 U3244 ( .A1(n13842), .A2(n13773), .B1(n13768), .B2(n14168), .ZN(
        n9725) );
  OAI22_X1 U3245 ( .A1(n13848), .A2(n13773), .B1(n13768), .B2(n14167), .ZN(
        n9726) );
  OAI22_X1 U3246 ( .A1(n13854), .A2(n13773), .B1(n13768), .B2(n14166), .ZN(
        n9727) );
  OAI22_X1 U3247 ( .A1(n13860), .A2(n13773), .B1(n13768), .B2(n14165), .ZN(
        n9728) );
  OAI22_X1 U3248 ( .A1(n13866), .A2(n13773), .B1(n13768), .B2(n14164), .ZN(
        n9729) );
  OAI22_X1 U3249 ( .A1(n13872), .A2(n13772), .B1(n13768), .B2(n14163), .ZN(
        n9730) );
  OAI22_X1 U3250 ( .A1(n13878), .A2(n13772), .B1(n13768), .B2(n14162), .ZN(
        n9731) );
  OAI22_X1 U3251 ( .A1(n13884), .A2(n13772), .B1(n13768), .B2(n14161), .ZN(
        n9732) );
  OAI22_X1 U3252 ( .A1(n13890), .A2(n13772), .B1(n13768), .B2(n14160), .ZN(
        n9733) );
  OAI22_X1 U3253 ( .A1(n13896), .A2(n13772), .B1(n13769), .B2(n14159), .ZN(
        n9734) );
  OAI22_X1 U3254 ( .A1(n13902), .A2(n13772), .B1(n13769), .B2(n14158), .ZN(
        n9735) );
  OAI22_X1 U3255 ( .A1(n13908), .A2(n13772), .B1(n13769), .B2(n14157), .ZN(
        n9736) );
  OAI22_X1 U3256 ( .A1(n13914), .A2(n13772), .B1(n13769), .B2(n14156), .ZN(
        n9737) );
  OAI22_X1 U3257 ( .A1(n13920), .A2(n13772), .B1(n13769), .B2(n14155), .ZN(
        n9738) );
  OAI22_X1 U3258 ( .A1(n13926), .A2(n13772), .B1(n13769), .B2(n14154), .ZN(
        n9739) );
  OAI22_X1 U3259 ( .A1(n13932), .A2(n13772), .B1(n13769), .B2(n14153), .ZN(
        n9740) );
  OAI22_X1 U3260 ( .A1(n13938), .A2(n13772), .B1(n13769), .B2(n14152), .ZN(
        n9741) );
  OAI22_X1 U3261 ( .A1(n13944), .A2(n13771), .B1(n13769), .B2(n14151), .ZN(
        n9742) );
  OAI22_X1 U3262 ( .A1(n13950), .A2(n13771), .B1(n13769), .B2(n14150), .ZN(
        n9743) );
  OAI22_X1 U3263 ( .A1(n13956), .A2(n13771), .B1(n13769), .B2(n14149), .ZN(
        n9744) );
  OAI22_X1 U3264 ( .A1(n13962), .A2(n13771), .B1(n13769), .B2(n14148), .ZN(
        n9745) );
  OAI22_X1 U3265 ( .A1(n13824), .A2(n13779), .B1(n13774), .B2(n14139), .ZN(
        n9754) );
  OAI22_X1 U3266 ( .A1(n13830), .A2(n13779), .B1(n13774), .B2(n14138), .ZN(
        n9755) );
  OAI22_X1 U3267 ( .A1(n13836), .A2(n13779), .B1(n13774), .B2(n14137), .ZN(
        n9756) );
  OAI22_X1 U3268 ( .A1(n13842), .A2(n13779), .B1(n13774), .B2(n14136), .ZN(
        n9757) );
  OAI22_X1 U3269 ( .A1(n13848), .A2(n13779), .B1(n13774), .B2(n14135), .ZN(
        n9758) );
  OAI22_X1 U3270 ( .A1(n13854), .A2(n13779), .B1(n13774), .B2(n14134), .ZN(
        n9759) );
  OAI22_X1 U3271 ( .A1(n13860), .A2(n13779), .B1(n13774), .B2(n14133), .ZN(
        n9760) );
  OAI22_X1 U3272 ( .A1(n13866), .A2(n13779), .B1(n13774), .B2(n14132), .ZN(
        n9761) );
  OAI22_X1 U3273 ( .A1(n13872), .A2(n13778), .B1(n13774), .B2(n14131), .ZN(
        n9762) );
  OAI22_X1 U3274 ( .A1(n13878), .A2(n13778), .B1(n13774), .B2(n14130), .ZN(
        n9763) );
  OAI22_X1 U3275 ( .A1(n13884), .A2(n13778), .B1(n13774), .B2(n14129), .ZN(
        n9764) );
  OAI22_X1 U3276 ( .A1(n13890), .A2(n13778), .B1(n13774), .B2(n14128), .ZN(
        n9765) );
  OAI22_X1 U3277 ( .A1(n13896), .A2(n13778), .B1(n13775), .B2(n14127), .ZN(
        n9766) );
  OAI22_X1 U3278 ( .A1(n13902), .A2(n13778), .B1(n13775), .B2(n14126), .ZN(
        n9767) );
  OAI22_X1 U3279 ( .A1(n13908), .A2(n13778), .B1(n13775), .B2(n14125), .ZN(
        n9768) );
  OAI22_X1 U3280 ( .A1(n13914), .A2(n13778), .B1(n13775), .B2(n14124), .ZN(
        n9769) );
  OAI22_X1 U3281 ( .A1(n13920), .A2(n13778), .B1(n13775), .B2(n14123), .ZN(
        n9770) );
  OAI22_X1 U3282 ( .A1(n13926), .A2(n13778), .B1(n13775), .B2(n14122), .ZN(
        n9771) );
  OAI22_X1 U3283 ( .A1(n13932), .A2(n13778), .B1(n13775), .B2(n14121), .ZN(
        n9772) );
  OAI22_X1 U3284 ( .A1(n13938), .A2(n13778), .B1(n13775), .B2(n14120), .ZN(
        n9773) );
  OAI22_X1 U3285 ( .A1(n13944), .A2(n13777), .B1(n13775), .B2(n14119), .ZN(
        n9774) );
  OAI22_X1 U3286 ( .A1(n13950), .A2(n13777), .B1(n13775), .B2(n14118), .ZN(
        n9775) );
  OAI22_X1 U3287 ( .A1(n13956), .A2(n13777), .B1(n13775), .B2(n14117), .ZN(
        n9776) );
  OAI22_X1 U3288 ( .A1(n13962), .A2(n13777), .B1(n13775), .B2(n14116), .ZN(
        n9777) );
  OAI22_X1 U3289 ( .A1(n13824), .A2(n13803), .B1(n13798), .B2(n12662), .ZN(
        n9882) );
  OAI22_X1 U3290 ( .A1(n13830), .A2(n13803), .B1(n13798), .B2(n12664), .ZN(
        n9883) );
  OAI22_X1 U3291 ( .A1(n13836), .A2(n13803), .B1(n13798), .B2(n12666), .ZN(
        n9884) );
  OAI22_X1 U3292 ( .A1(n13842), .A2(n13803), .B1(n13798), .B2(n12668), .ZN(
        n9885) );
  OAI22_X1 U3293 ( .A1(n13848), .A2(n13803), .B1(n13798), .B2(n12670), .ZN(
        n9886) );
  OAI22_X1 U3294 ( .A1(n13854), .A2(n13803), .B1(n13798), .B2(n12672), .ZN(
        n9887) );
  OAI22_X1 U3295 ( .A1(n13860), .A2(n13803), .B1(n13798), .B2(n12674), .ZN(
        n9888) );
  OAI22_X1 U3296 ( .A1(n13866), .A2(n13803), .B1(n13798), .B2(n12676), .ZN(
        n9889) );
  OAI22_X1 U3297 ( .A1(n13872), .A2(n13802), .B1(n13798), .B2(n12678), .ZN(
        n9890) );
  OAI22_X1 U3298 ( .A1(n13878), .A2(n13802), .B1(n13798), .B2(n12680), .ZN(
        n9891) );
  OAI22_X1 U3299 ( .A1(n13884), .A2(n13802), .B1(n13798), .B2(n12682), .ZN(
        n9892) );
  OAI22_X1 U3300 ( .A1(n13890), .A2(n13802), .B1(n13798), .B2(n12684), .ZN(
        n9893) );
  OAI22_X1 U3301 ( .A1(n13896), .A2(n13802), .B1(n13799), .B2(n12686), .ZN(
        n9894) );
  OAI22_X1 U3302 ( .A1(n13902), .A2(n13802), .B1(n13799), .B2(n12688), .ZN(
        n9895) );
  OAI22_X1 U3303 ( .A1(n13908), .A2(n13802), .B1(n13799), .B2(n12690), .ZN(
        n9896) );
  OAI22_X1 U3304 ( .A1(n13914), .A2(n13802), .B1(n13799), .B2(n12692), .ZN(
        n9897) );
  OAI22_X1 U3305 ( .A1(n13920), .A2(n13802), .B1(n13799), .B2(n12694), .ZN(
        n9898) );
  OAI22_X1 U3306 ( .A1(n13926), .A2(n13802), .B1(n13799), .B2(n12696), .ZN(
        n9899) );
  OAI22_X1 U3307 ( .A1(n13932), .A2(n13802), .B1(n13799), .B2(n12698), .ZN(
        n9900) );
  OAI22_X1 U3308 ( .A1(n13938), .A2(n13802), .B1(n13799), .B2(n12700), .ZN(
        n9901) );
  OAI22_X1 U3309 ( .A1(n13944), .A2(n13801), .B1(n13799), .B2(n12702), .ZN(
        n9902) );
  OAI22_X1 U3310 ( .A1(n13950), .A2(n13801), .B1(n13799), .B2(n12704), .ZN(
        n9903) );
  OAI22_X1 U3311 ( .A1(n13956), .A2(n13801), .B1(n13799), .B2(n12706), .ZN(
        n9904) );
  OAI22_X1 U3312 ( .A1(n13962), .A2(n13801), .B1(n13799), .B2(n12708), .ZN(
        n9905) );
  OAI22_X1 U3313 ( .A1(n13387), .A2(n15548), .B1(n13878), .B2(n13385), .ZN(
        n7683) );
  OAI22_X1 U3314 ( .A1(n13387), .A2(n15547), .B1(n13884), .B2(n13385), .ZN(
        n7684) );
  OAI22_X1 U3315 ( .A1(n13387), .A2(n15546), .B1(n13890), .B2(n13385), .ZN(
        n7685) );
  OAI22_X1 U3316 ( .A1(n13388), .A2(n15545), .B1(n13896), .B2(n13385), .ZN(
        n7686) );
  OAI22_X1 U3317 ( .A1(n13388), .A2(n15544), .B1(n13902), .B2(n13385), .ZN(
        n7687) );
  OAI22_X1 U3318 ( .A1(n13388), .A2(n15543), .B1(n13908), .B2(n13385), .ZN(
        n7688) );
  OAI22_X1 U3319 ( .A1(n13388), .A2(n15542), .B1(n13914), .B2(n13385), .ZN(
        n7689) );
  OAI22_X1 U3320 ( .A1(n13388), .A2(n15541), .B1(n13920), .B2(n13385), .ZN(
        n7690) );
  OAI22_X1 U3321 ( .A1(n13388), .A2(n15540), .B1(n13926), .B2(n13385), .ZN(
        n7691) );
  OAI22_X1 U3322 ( .A1(n13388), .A2(n15539), .B1(n13932), .B2(n13385), .ZN(
        n7692) );
  OAI22_X1 U3323 ( .A1(n13388), .A2(n15538), .B1(n13938), .B2(n13385), .ZN(
        n7693) );
  OAI22_X1 U3324 ( .A1(n13388), .A2(n15537), .B1(n13944), .B2(n13384), .ZN(
        n7694) );
  OAI22_X1 U3325 ( .A1(n13388), .A2(n15536), .B1(n13950), .B2(n13384), .ZN(
        n7695) );
  OAI22_X1 U3326 ( .A1(n13388), .A2(n15535), .B1(n13956), .B2(n13384), .ZN(
        n7696) );
  OAI22_X1 U3327 ( .A1(n13388), .A2(n15534), .B1(n13962), .B2(n13384), .ZN(
        n7697) );
  OAI22_X1 U3328 ( .A1(n13389), .A2(n15533), .B1(n13968), .B2(n13384), .ZN(
        n7698) );
  OAI22_X1 U3329 ( .A1(n13389), .A2(n15532), .B1(n13974), .B2(n13384), .ZN(
        n7699) );
  OAI22_X1 U3330 ( .A1(n13389), .A2(n15531), .B1(n13980), .B2(n13384), .ZN(
        n7700) );
  OAI22_X1 U3331 ( .A1(n13389), .A2(n15530), .B1(n13986), .B2(n13384), .ZN(
        n7701) );
  OAI22_X1 U3332 ( .A1(n13389), .A2(n15529), .B1(n13992), .B2(n13384), .ZN(
        n7702) );
  OAI22_X1 U3333 ( .A1(n13389), .A2(n15528), .B1(n13998), .B2(n13384), .ZN(
        n7703) );
  OAI22_X1 U3334 ( .A1(n13389), .A2(n15527), .B1(n14004), .B2(n13384), .ZN(
        n7704) );
  OAI22_X1 U3335 ( .A1(n13389), .A2(n15526), .B1(n14013), .B2(n13385), .ZN(
        n7705) );
  NAND4_X1 U3336 ( .A1(n3229), .A2(n3230), .A3(n3231), .A4(n3232), .ZN(n3228)
         );
  AOI221_X1 U3337 ( .B1(n13329), .B2(n14047), .C1(n13326), .C2(n14031), .A(
        n3236), .ZN(n3229) );
  AOI221_X1 U3338 ( .B1(n13356), .B2(n14219), .C1(n13353), .C2(n14207), .A(
        n3234), .ZN(n3231) );
  AOI221_X1 U3339 ( .B1(n13344), .B2(n14079), .C1(n13341), .C2(n15601), .A(
        n3235), .ZN(n3230) );
  NAND4_X1 U3340 ( .A1(n3192), .A2(n3193), .A3(n3194), .A4(n3195), .ZN(n3191)
         );
  AOI221_X1 U3341 ( .B1(n13329), .B2(n14046), .C1(n13326), .C2(n14030), .A(
        n3199), .ZN(n3192) );
  AOI221_X1 U3342 ( .B1(n13356), .B2(n14218), .C1(n13353), .C2(n14206), .A(
        n3197), .ZN(n3194) );
  AOI221_X1 U3343 ( .B1(n13344), .B2(n14078), .C1(n13341), .C2(n15600), .A(
        n3198), .ZN(n3193) );
  NAND4_X1 U3344 ( .A1(n3155), .A2(n3156), .A3(n3157), .A4(n3158), .ZN(n3154)
         );
  AOI221_X1 U3345 ( .B1(n13329), .B2(n14045), .C1(n13326), .C2(n14029), .A(
        n3162), .ZN(n3155) );
  AOI221_X1 U3346 ( .B1(n13356), .B2(n14217), .C1(n13353), .C2(n14205), .A(
        n3160), .ZN(n3157) );
  AOI221_X1 U3347 ( .B1(n13344), .B2(n14077), .C1(n13341), .C2(n15599), .A(
        n3161), .ZN(n3156) );
  NAND4_X1 U3348 ( .A1(n3046), .A2(n3047), .A3(n3048), .A4(n3049), .ZN(n3045)
         );
  AOI221_X1 U3349 ( .B1(n13329), .B2(n14044), .C1(n13326), .C2(n14028), .A(
        n3069), .ZN(n3046) );
  AOI221_X1 U3350 ( .B1(n13356), .B2(n14216), .C1(n13353), .C2(n14204), .A(
        n3058), .ZN(n3048) );
  AOI221_X1 U3351 ( .B1(n13344), .B2(n14076), .C1(n13341), .C2(n15598), .A(
        n3063), .ZN(n3047) );
  NAND4_X1 U3352 ( .A1(n4265), .A2(n4266), .A3(n4267), .A4(n4268), .ZN(n4264)
         );
  AOI221_X1 U3353 ( .B1(n13327), .B2(n14075), .C1(n13324), .C2(n16042), .A(
        n4283), .ZN(n4265) );
  AOI221_X1 U3354 ( .B1(n13354), .B2(n14247), .C1(n13351), .C2(n16006), .A(
        n4277), .ZN(n4267) );
  AOI221_X1 U3355 ( .B1(n13342), .B2(n14107), .C1(n13339), .C2(n15921), .A(
        n4281), .ZN(n4266) );
  NAND4_X1 U3356 ( .A1(n4228), .A2(n4229), .A3(n4230), .A4(n4231), .ZN(n4227)
         );
  AOI221_X1 U3357 ( .B1(n13327), .B2(n14074), .C1(n13324), .C2(n16041), .A(
        n4235), .ZN(n4228) );
  AOI221_X1 U3358 ( .B1(n13354), .B2(n14246), .C1(n13351), .C2(n16005), .A(
        n4233), .ZN(n4230) );
  AOI221_X1 U3359 ( .B1(n13342), .B2(n14106), .C1(n13339), .C2(n15920), .A(
        n4234), .ZN(n4229) );
  NAND4_X1 U3360 ( .A1(n4191), .A2(n4192), .A3(n4193), .A4(n4194), .ZN(n4190)
         );
  AOI221_X1 U3361 ( .B1(n13327), .B2(n14073), .C1(n13324), .C2(n16040), .A(
        n4198), .ZN(n4191) );
  AOI221_X1 U3362 ( .B1(n13354), .B2(n14245), .C1(n13351), .C2(n16004), .A(
        n4196), .ZN(n4193) );
  AOI221_X1 U3363 ( .B1(n13342), .B2(n14105), .C1(n13339), .C2(n15919), .A(
        n4197), .ZN(n4192) );
  NAND4_X1 U3364 ( .A1(n4154), .A2(n4155), .A3(n4156), .A4(n4157), .ZN(n4153)
         );
  AOI221_X1 U3365 ( .B1(n13327), .B2(n14072), .C1(n13324), .C2(n16039), .A(
        n4161), .ZN(n4154) );
  AOI221_X1 U3366 ( .B1(n13354), .B2(n14244), .C1(n13351), .C2(n16003), .A(
        n4159), .ZN(n4156) );
  AOI221_X1 U3367 ( .B1(n13342), .B2(n14104), .C1(n13339), .C2(n15918), .A(
        n4160), .ZN(n4155) );
  NAND4_X1 U3368 ( .A1(n4117), .A2(n4118), .A3(n4119), .A4(n4120), .ZN(n4116)
         );
  AOI221_X1 U3369 ( .B1(n13327), .B2(n14071), .C1(n13324), .C2(n16038), .A(
        n4124), .ZN(n4117) );
  AOI221_X1 U3370 ( .B1(n13354), .B2(n14243), .C1(n13351), .C2(n16002), .A(
        n4122), .ZN(n4119) );
  AOI221_X1 U3371 ( .B1(n13342), .B2(n14103), .C1(n13339), .C2(n15917), .A(
        n4123), .ZN(n4118) );
  NAND4_X1 U3372 ( .A1(n4080), .A2(n4081), .A3(n4082), .A4(n4083), .ZN(n4079)
         );
  AOI221_X1 U3373 ( .B1(n13327), .B2(n14070), .C1(n13324), .C2(n16037), .A(
        n4087), .ZN(n4080) );
  AOI221_X1 U3374 ( .B1(n13354), .B2(n14242), .C1(n13351), .C2(n16001), .A(
        n4085), .ZN(n4082) );
  AOI221_X1 U3375 ( .B1(n13342), .B2(n14102), .C1(n13339), .C2(n15916), .A(
        n4086), .ZN(n4081) );
  NAND4_X1 U3376 ( .A1(n4043), .A2(n4044), .A3(n4045), .A4(n4046), .ZN(n4042)
         );
  AOI221_X1 U3377 ( .B1(n13327), .B2(n14069), .C1(n13324), .C2(n16036), .A(
        n4050), .ZN(n4043) );
  AOI221_X1 U3378 ( .B1(n13354), .B2(n14241), .C1(n13351), .C2(n16000), .A(
        n4048), .ZN(n4045) );
  AOI221_X1 U3379 ( .B1(n13342), .B2(n14101), .C1(n13339), .C2(n15915), .A(
        n4049), .ZN(n4044) );
  NAND4_X1 U3380 ( .A1(n4006), .A2(n4007), .A3(n4008), .A4(n4009), .ZN(n4005)
         );
  AOI221_X1 U3381 ( .B1(n13327), .B2(n14068), .C1(n13324), .C2(n16035), .A(
        n4013), .ZN(n4006) );
  AOI221_X1 U3382 ( .B1(n13354), .B2(n14240), .C1(n13351), .C2(n15999), .A(
        n4011), .ZN(n4008) );
  AOI221_X1 U3383 ( .B1(n13342), .B2(n14100), .C1(n13339), .C2(n15914), .A(
        n4012), .ZN(n4007) );
  NAND4_X1 U3384 ( .A1(n3969), .A2(n3970), .A3(n3971), .A4(n3972), .ZN(n3968)
         );
  AOI221_X1 U3385 ( .B1(n13327), .B2(n14067), .C1(n13324), .C2(n16034), .A(
        n3976), .ZN(n3969) );
  AOI221_X1 U3386 ( .B1(n13354), .B2(n14239), .C1(n13351), .C2(n15998), .A(
        n3974), .ZN(n3971) );
  AOI221_X1 U3387 ( .B1(n13342), .B2(n14099), .C1(n13339), .C2(n15913), .A(
        n3975), .ZN(n3970) );
  NAND4_X1 U3388 ( .A1(n3932), .A2(n3933), .A3(n3934), .A4(n3935), .ZN(n3931)
         );
  AOI221_X1 U3389 ( .B1(n13327), .B2(n14066), .C1(n13324), .C2(n16033), .A(
        n3939), .ZN(n3932) );
  AOI221_X1 U3390 ( .B1(n13354), .B2(n14238), .C1(n13351), .C2(n15997), .A(
        n3937), .ZN(n3934) );
  AOI221_X1 U3391 ( .B1(n13342), .B2(n14098), .C1(n13339), .C2(n15912), .A(
        n3938), .ZN(n3933) );
  NAND4_X1 U3392 ( .A1(n3895), .A2(n3896), .A3(n3897), .A4(n3898), .ZN(n3894)
         );
  AOI221_X1 U3393 ( .B1(n13327), .B2(n14065), .C1(n13324), .C2(n16032), .A(
        n3902), .ZN(n3895) );
  AOI221_X1 U3394 ( .B1(n13354), .B2(n14237), .C1(n13351), .C2(n15996), .A(
        n3900), .ZN(n3897) );
  AOI221_X1 U3395 ( .B1(n13342), .B2(n14097), .C1(n13339), .C2(n15911), .A(
        n3901), .ZN(n3896) );
  NAND4_X1 U3396 ( .A1(n3858), .A2(n3859), .A3(n3860), .A4(n3861), .ZN(n3857)
         );
  AOI221_X1 U3397 ( .B1(n13327), .B2(n14064), .C1(n13324), .C2(n16031), .A(
        n3865), .ZN(n3858) );
  AOI221_X1 U3398 ( .B1(n13354), .B2(n14236), .C1(n13351), .C2(n15995), .A(
        n3863), .ZN(n3860) );
  AOI221_X1 U3399 ( .B1(n13342), .B2(n14096), .C1(n13339), .C2(n15910), .A(
        n3864), .ZN(n3859) );
  NAND4_X1 U3400 ( .A1(n3821), .A2(n3822), .A3(n3823), .A4(n3824), .ZN(n3820)
         );
  AOI221_X1 U3401 ( .B1(n13328), .B2(n14063), .C1(n13325), .C2(n16054), .A(
        n3828), .ZN(n3821) );
  AOI221_X1 U3402 ( .B1(n13355), .B2(n14235), .C1(n13352), .C2(n16050), .A(
        n3826), .ZN(n3823) );
  AOI221_X1 U3403 ( .B1(n13343), .B2(n14095), .C1(n13340), .C2(n15909), .A(
        n3827), .ZN(n3822) );
  NAND4_X1 U3404 ( .A1(n3784), .A2(n3785), .A3(n3786), .A4(n3787), .ZN(n3783)
         );
  AOI221_X1 U3405 ( .B1(n13328), .B2(n14062), .C1(n13325), .C2(n16053), .A(
        n3791), .ZN(n3784) );
  AOI221_X1 U3406 ( .B1(n13355), .B2(n14234), .C1(n13352), .C2(n16049), .A(
        n3789), .ZN(n3786) );
  AOI221_X1 U3407 ( .B1(n13343), .B2(n14094), .C1(n13340), .C2(n15908), .A(
        n3790), .ZN(n3785) );
  NAND4_X1 U3408 ( .A1(n3747), .A2(n3748), .A3(n3749), .A4(n3750), .ZN(n3746)
         );
  AOI221_X1 U3409 ( .B1(n13328), .B2(n14061), .C1(n13325), .C2(n16052), .A(
        n3754), .ZN(n3747) );
  AOI221_X1 U3410 ( .B1(n13355), .B2(n14233), .C1(n13352), .C2(n16048), .A(
        n3752), .ZN(n3749) );
  AOI221_X1 U3411 ( .B1(n13343), .B2(n14093), .C1(n13340), .C2(n15907), .A(
        n3753), .ZN(n3748) );
  NAND4_X1 U3412 ( .A1(n3710), .A2(n3711), .A3(n3712), .A4(n3713), .ZN(n3709)
         );
  AOI221_X1 U3413 ( .B1(n13328), .B2(n14060), .C1(n13325), .C2(n16051), .A(
        n3717), .ZN(n3710) );
  AOI221_X1 U3414 ( .B1(n13355), .B2(n14232), .C1(n13352), .C2(n16047), .A(
        n3715), .ZN(n3712) );
  AOI221_X1 U3415 ( .B1(n13343), .B2(n14092), .C1(n13340), .C2(n15906), .A(
        n3716), .ZN(n3711) );
  NAND4_X1 U3416 ( .A1(n3673), .A2(n3674), .A3(n3675), .A4(n3676), .ZN(n3672)
         );
  AOI221_X1 U3417 ( .B1(n13328), .B2(n14059), .C1(n13325), .C2(n14043), .A(
        n3680), .ZN(n3673) );
  AOI221_X1 U3418 ( .B1(n13355), .B2(n14231), .C1(n13352), .C2(n16046), .A(
        n3678), .ZN(n3675) );
  AOI221_X1 U3419 ( .B1(n13343), .B2(n14091), .C1(n13340), .C2(n15905), .A(
        n3679), .ZN(n3674) );
  NAND4_X1 U3420 ( .A1(n3636), .A2(n3637), .A3(n3638), .A4(n3639), .ZN(n3635)
         );
  AOI221_X1 U3421 ( .B1(n13328), .B2(n14058), .C1(n13325), .C2(n14042), .A(
        n3643), .ZN(n3636) );
  AOI221_X1 U3422 ( .B1(n13355), .B2(n14230), .C1(n13352), .C2(n16045), .A(
        n3641), .ZN(n3638) );
  AOI221_X1 U3423 ( .B1(n13343), .B2(n14090), .C1(n13340), .C2(n15904), .A(
        n3642), .ZN(n3637) );
  NAND4_X1 U3424 ( .A1(n3599), .A2(n3600), .A3(n3601), .A4(n3602), .ZN(n3598)
         );
  AOI221_X1 U3425 ( .B1(n13328), .B2(n14057), .C1(n13325), .C2(n14041), .A(
        n3606), .ZN(n3599) );
  AOI221_X1 U3426 ( .B1(n13355), .B2(n14229), .C1(n13352), .C2(n16044), .A(
        n3604), .ZN(n3601) );
  AOI221_X1 U3427 ( .B1(n13343), .B2(n14089), .C1(n13340), .C2(n15903), .A(
        n3605), .ZN(n3600) );
  NAND4_X1 U3428 ( .A1(n3562), .A2(n3563), .A3(n3564), .A4(n3565), .ZN(n3561)
         );
  AOI221_X1 U3429 ( .B1(n13328), .B2(n14056), .C1(n13325), .C2(n14040), .A(
        n3569), .ZN(n3562) );
  AOI221_X1 U3430 ( .B1(n13355), .B2(n14228), .C1(n13352), .C2(n16043), .A(
        n3567), .ZN(n3564) );
  AOI221_X1 U3431 ( .B1(n13343), .B2(n14088), .C1(n13340), .C2(n15902), .A(
        n3568), .ZN(n3563) );
  NAND4_X1 U3432 ( .A1(n3525), .A2(n3526), .A3(n3527), .A4(n3528), .ZN(n3524)
         );
  AOI221_X1 U3433 ( .B1(n13328), .B2(n14055), .C1(n13325), .C2(n14039), .A(
        n3532), .ZN(n3525) );
  AOI221_X1 U3434 ( .B1(n13355), .B2(n14227), .C1(n13352), .C2(n14215), .A(
        n3530), .ZN(n3527) );
  AOI221_X1 U3435 ( .B1(n13343), .B2(n14087), .C1(n13340), .C2(n15901), .A(
        n3531), .ZN(n3526) );
  NAND4_X1 U3436 ( .A1(n3488), .A2(n3489), .A3(n3490), .A4(n3491), .ZN(n3487)
         );
  AOI221_X1 U3437 ( .B1(n13328), .B2(n14054), .C1(n13325), .C2(n14038), .A(
        n3495), .ZN(n3488) );
  AOI221_X1 U3438 ( .B1(n13355), .B2(n14226), .C1(n13352), .C2(n14214), .A(
        n3493), .ZN(n3490) );
  AOI221_X1 U3439 ( .B1(n13343), .B2(n14086), .C1(n13340), .C2(n15900), .A(
        n3494), .ZN(n3489) );
  NAND4_X1 U3440 ( .A1(n3451), .A2(n3452), .A3(n3453), .A4(n3454), .ZN(n3450)
         );
  AOI221_X1 U3441 ( .B1(n13328), .B2(n14053), .C1(n13325), .C2(n14037), .A(
        n3458), .ZN(n3451) );
  AOI221_X1 U3442 ( .B1(n13355), .B2(n14225), .C1(n13352), .C2(n14213), .A(
        n3456), .ZN(n3453) );
  AOI221_X1 U3443 ( .B1(n13343), .B2(n14085), .C1(n13340), .C2(n15899), .A(
        n3457), .ZN(n3452) );
  NAND4_X1 U3444 ( .A1(n3414), .A2(n3415), .A3(n3416), .A4(n3417), .ZN(n3413)
         );
  AOI221_X1 U3445 ( .B1(n13328), .B2(n14052), .C1(n13325), .C2(n14036), .A(
        n3421), .ZN(n3414) );
  AOI221_X1 U3446 ( .B1(n13355), .B2(n14224), .C1(n13352), .C2(n14212), .A(
        n3419), .ZN(n3416) );
  AOI221_X1 U3447 ( .B1(n13343), .B2(n14084), .C1(n13340), .C2(n15898), .A(
        n3420), .ZN(n3415) );
  NAND4_X1 U3448 ( .A1(n3377), .A2(n3378), .A3(n3379), .A4(n3380), .ZN(n3376)
         );
  AOI221_X1 U3449 ( .B1(n13329), .B2(n14051), .C1(n13326), .C2(n14035), .A(
        n3384), .ZN(n3377) );
  AOI221_X1 U3450 ( .B1(n13356), .B2(n14223), .C1(n13353), .C2(n14211), .A(
        n3382), .ZN(n3379) );
  AOI221_X1 U3451 ( .B1(n13344), .B2(n14083), .C1(n13341), .C2(n15605), .A(
        n3383), .ZN(n3378) );
  NAND4_X1 U3452 ( .A1(n3340), .A2(n3341), .A3(n3342), .A4(n3343), .ZN(n3339)
         );
  AOI221_X1 U3453 ( .B1(n13329), .B2(n14050), .C1(n13326), .C2(n14034), .A(
        n3347), .ZN(n3340) );
  AOI221_X1 U3454 ( .B1(n13356), .B2(n14222), .C1(n13353), .C2(n14210), .A(
        n3345), .ZN(n3342) );
  AOI221_X1 U3455 ( .B1(n13344), .B2(n14082), .C1(n13341), .C2(n15604), .A(
        n3346), .ZN(n3341) );
  NAND4_X1 U3456 ( .A1(n3303), .A2(n3304), .A3(n3305), .A4(n3306), .ZN(n3302)
         );
  AOI221_X1 U3457 ( .B1(n13329), .B2(n14049), .C1(n13326), .C2(n14033), .A(
        n3310), .ZN(n3303) );
  AOI221_X1 U3458 ( .B1(n13356), .B2(n14221), .C1(n13353), .C2(n14209), .A(
        n3308), .ZN(n3305) );
  AOI221_X1 U3459 ( .B1(n13344), .B2(n14081), .C1(n13341), .C2(n15603), .A(
        n3309), .ZN(n3304) );
  NAND4_X1 U3460 ( .A1(n3266), .A2(n3267), .A3(n3268), .A4(n3269), .ZN(n3265)
         );
  AOI221_X1 U3461 ( .B1(n13329), .B2(n14048), .C1(n13326), .C2(n14032), .A(
        n3273), .ZN(n3266) );
  AOI221_X1 U3462 ( .B1(n13356), .B2(n14220), .C1(n13353), .C2(n14208), .A(
        n3271), .ZN(n3268) );
  AOI221_X1 U3463 ( .B1(n13344), .B2(n14080), .C1(n13341), .C2(n15602), .A(
        n3272), .ZN(n3267) );
  NAND4_X1 U3464 ( .A1(n3237), .A2(n3238), .A3(n3239), .A4(n3240), .ZN(n3227)
         );
  AOI221_X1 U3465 ( .B1(n13275), .B2(n15865), .C1(n13272), .C2(n15628), .A(
        n3244), .ZN(n3237) );
  AOI221_X1 U3466 ( .B1(n13302), .B2(n15577), .C1(n13299), .C2(n15793), .A(
        n3242), .ZN(n3239) );
  AOI221_X1 U3467 ( .B1(n13290), .B2(n14464), .C1(n13287), .C2(n15585), .A(
        n3243), .ZN(n3238) );
  NAND4_X1 U3468 ( .A1(n3200), .A2(n3201), .A3(n3202), .A4(n3203), .ZN(n3190)
         );
  AOI221_X1 U3469 ( .B1(n13275), .B2(n15864), .C1(n13272), .C2(n15627), .A(
        n3207), .ZN(n3200) );
  AOI221_X1 U3470 ( .B1(n13302), .B2(n15576), .C1(n13299), .C2(n15792), .A(
        n3205), .ZN(n3202) );
  AOI221_X1 U3471 ( .B1(n13290), .B2(n14463), .C1(n13287), .C2(n15584), .A(
        n3206), .ZN(n3201) );
  NAND4_X1 U3472 ( .A1(n4632), .A2(n4633), .A3(n4634), .A4(n4635), .ZN(n4622)
         );
  AOI221_X1 U3473 ( .B1(n13047), .B2(n15868), .C1(n13044), .C2(n15631), .A(
        n4639), .ZN(n4632) );
  AOI221_X1 U3474 ( .B1(n13074), .B2(n15796), .C1(n13071), .C2(n15580), .A(
        n4637), .ZN(n4634) );
  AOI221_X1 U3475 ( .B1(n13062), .B2(n14467), .C1(n13059), .C2(n15588), .A(
        n4638), .ZN(n4633) );
  NAND4_X1 U3476 ( .A1(n4595), .A2(n4596), .A3(n4597), .A4(n4598), .ZN(n4585)
         );
  AOI221_X1 U3477 ( .B1(n13047), .B2(n15867), .C1(n13044), .C2(n15630), .A(
        n4602), .ZN(n4595) );
  AOI221_X1 U3478 ( .B1(n13074), .B2(n15795), .C1(n13071), .C2(n15579), .A(
        n4600), .ZN(n4597) );
  AOI221_X1 U3479 ( .B1(n13062), .B2(n14466), .C1(n13059), .C2(n15587), .A(
        n4601), .ZN(n4596) );
  NAND4_X1 U3480 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n4548)
         );
  AOI221_X1 U3481 ( .B1(n13047), .B2(n15866), .C1(n13044), .C2(n15629), .A(
        n4565), .ZN(n4558) );
  AOI221_X1 U3482 ( .B1(n13074), .B2(n15794), .C1(n13071), .C2(n15578), .A(
        n4563), .ZN(n4560) );
  AOI221_X1 U3483 ( .B1(n13062), .B2(n14465), .C1(n13059), .C2(n15586), .A(
        n4564), .ZN(n4559) );
  NAND4_X1 U3484 ( .A1(n4521), .A2(n4522), .A3(n4523), .A4(n4524), .ZN(n4511)
         );
  AOI221_X1 U3485 ( .B1(n13047), .B2(n15865), .C1(n13044), .C2(n15628), .A(
        n4528), .ZN(n4521) );
  AOI221_X1 U3486 ( .B1(n13074), .B2(n15793), .C1(n13071), .C2(n15577), .A(
        n4526), .ZN(n4523) );
  AOI221_X1 U3487 ( .B1(n13062), .B2(n14464), .C1(n13059), .C2(n15585), .A(
        n4527), .ZN(n4522) );
  NAND4_X1 U3488 ( .A1(n4484), .A2(n4485), .A3(n4486), .A4(n4487), .ZN(n4474)
         );
  AOI221_X1 U3489 ( .B1(n13047), .B2(n15864), .C1(n13044), .C2(n15627), .A(
        n4491), .ZN(n4484) );
  AOI221_X1 U3490 ( .B1(n13074), .B2(n15792), .C1(n13071), .C2(n15576), .A(
        n4489), .ZN(n4486) );
  AOI221_X1 U3491 ( .B1(n13062), .B2(n14463), .C1(n13059), .C2(n15584), .A(
        n4490), .ZN(n4485) );
  NAND4_X1 U3492 ( .A1(n5681), .A2(n5684), .A3(n5686), .A4(n5688), .ZN(n5648)
         );
  AOI221_X1 U3493 ( .B1(n13045), .B2(n14458), .C1(n13042), .C2(n15861), .A(
        n5698), .ZN(n5681) );
  AOI221_X1 U3494 ( .B1(n13072), .B2(n14659), .C1(n13069), .C2(n15789), .A(
        n5694), .ZN(n5686) );
  AOI221_X1 U3495 ( .B1(n13060), .B2(n14492), .C1(n13057), .C2(n15837), .A(
        n5696), .ZN(n5684) );
  NAND4_X1 U3496 ( .A1(n5601), .A2(n5604), .A3(n5606), .A4(n5608), .ZN(n5586)
         );
  AOI221_X1 U3497 ( .B1(n13045), .B2(n14457), .C1(n13042), .C2(n15860), .A(
        n5614), .ZN(n5601) );
  AOI221_X1 U3498 ( .B1(n13072), .B2(n14658), .C1(n13069), .C2(n15788), .A(
        n5610), .ZN(n5606) );
  AOI221_X1 U3499 ( .B1(n13060), .B2(n14491), .C1(n13057), .C2(n15836), .A(
        n5611), .ZN(n5604) );
  NAND4_X1 U3500 ( .A1(n5540), .A2(n5541), .A3(n5544), .A4(n5546), .ZN(n5524)
         );
  AOI221_X1 U3501 ( .B1(n13045), .B2(n14456), .C1(n13042), .C2(n15859), .A(
        n5551), .ZN(n5540) );
  AOI221_X1 U3502 ( .B1(n13072), .B2(n14657), .C1(n13069), .C2(n15787), .A(
        n5549), .ZN(n5544) );
  AOI221_X1 U3503 ( .B1(n13060), .B2(n14490), .C1(n13057), .C2(n15835), .A(
        n5550), .ZN(n5541) );
  NAND4_X1 U3504 ( .A1(n5479), .A2(n5480), .A3(n5481), .A4(n5484), .ZN(n5461)
         );
  AOI221_X1 U3505 ( .B1(n13045), .B2(n14455), .C1(n13042), .C2(n15858), .A(
        n5490), .ZN(n5479) );
  AOI221_X1 U3506 ( .B1(n13072), .B2(n14656), .C1(n13069), .C2(n15786), .A(
        n5488), .ZN(n5481) );
  AOI221_X1 U3507 ( .B1(n13060), .B2(n14489), .C1(n13057), .C2(n15834), .A(
        n5489), .ZN(n5480) );
  NAND4_X1 U3508 ( .A1(n5421), .A2(n5422), .A3(n5424), .A4(n5426), .ZN(n5408)
         );
  AOI221_X1 U3509 ( .B1(n13045), .B2(n14454), .C1(n13042), .C2(n15857), .A(
        n5431), .ZN(n5421) );
  AOI221_X1 U3510 ( .B1(n13072), .B2(n14655), .C1(n13069), .C2(n15785), .A(
        n5429), .ZN(n5424) );
  AOI221_X1 U3511 ( .B1(n13060), .B2(n14488), .C1(n13057), .C2(n15833), .A(
        n5430), .ZN(n5422) );
  NAND4_X1 U3512 ( .A1(n5372), .A2(n5373), .A3(n5374), .A4(n5375), .ZN(n5362)
         );
  AOI221_X1 U3513 ( .B1(n13045), .B2(n14453), .C1(n13042), .C2(n15856), .A(
        n5379), .ZN(n5372) );
  AOI221_X1 U3514 ( .B1(n13072), .B2(n14654), .C1(n13069), .C2(n15784), .A(
        n5377), .ZN(n5374) );
  AOI221_X1 U3515 ( .B1(n13060), .B2(n14487), .C1(n13057), .C2(n15832), .A(
        n5378), .ZN(n5373) );
  NAND4_X1 U3516 ( .A1(n5335), .A2(n5336), .A3(n5337), .A4(n5338), .ZN(n5325)
         );
  AOI221_X1 U3517 ( .B1(n13045), .B2(n14452), .C1(n13042), .C2(n15855), .A(
        n5342), .ZN(n5335) );
  AOI221_X1 U3518 ( .B1(n13072), .B2(n14653), .C1(n13069), .C2(n15783), .A(
        n5340), .ZN(n5337) );
  AOI221_X1 U3519 ( .B1(n13060), .B2(n14486), .C1(n13057), .C2(n15831), .A(
        n5341), .ZN(n5336) );
  NAND4_X1 U3520 ( .A1(n5298), .A2(n5299), .A3(n5300), .A4(n5301), .ZN(n5288)
         );
  AOI221_X1 U3521 ( .B1(n13045), .B2(n14451), .C1(n13042), .C2(n15854), .A(
        n5305), .ZN(n5298) );
  AOI221_X1 U3522 ( .B1(n13072), .B2(n15633), .C1(n13069), .C2(n15782), .A(
        n5303), .ZN(n5300) );
  AOI221_X1 U3523 ( .B1(n13060), .B2(n14485), .C1(n13057), .C2(n15830), .A(
        n5304), .ZN(n5299) );
  NAND4_X1 U3524 ( .A1(n5261), .A2(n5262), .A3(n5263), .A4(n5264), .ZN(n5251)
         );
  AOI221_X1 U3525 ( .B1(n13045), .B2(n14450), .C1(n13042), .C2(n15853), .A(
        n5268), .ZN(n5261) );
  AOI221_X1 U3526 ( .B1(n13072), .B2(n15813), .C1(n13069), .C2(n15781), .A(
        n5266), .ZN(n5263) );
  AOI221_X1 U3527 ( .B1(n13060), .B2(n14484), .C1(n13057), .C2(n15829), .A(
        n5267), .ZN(n5262) );
  NAND4_X1 U3528 ( .A1(n5224), .A2(n5225), .A3(n5226), .A4(n5227), .ZN(n5214)
         );
  AOI221_X1 U3529 ( .B1(n13045), .B2(n14449), .C1(n13042), .C2(n15852), .A(
        n5231), .ZN(n5224) );
  AOI221_X1 U3530 ( .B1(n13072), .B2(n15812), .C1(n13069), .C2(n15780), .A(
        n5229), .ZN(n5226) );
  AOI221_X1 U3531 ( .B1(n13060), .B2(n14483), .C1(n13057), .C2(n15828), .A(
        n5230), .ZN(n5225) );
  NAND4_X1 U3532 ( .A1(n5187), .A2(n5188), .A3(n5189), .A4(n5190), .ZN(n5177)
         );
  AOI221_X1 U3533 ( .B1(n13045), .B2(n14448), .C1(n13042), .C2(n15851), .A(
        n5194), .ZN(n5187) );
  AOI221_X1 U3534 ( .B1(n13072), .B2(n15811), .C1(n13069), .C2(n15779), .A(
        n5192), .ZN(n5189) );
  AOI221_X1 U3535 ( .B1(n13060), .B2(n14482), .C1(n13057), .C2(n15827), .A(
        n5193), .ZN(n5188) );
  NAND4_X1 U3536 ( .A1(n5150), .A2(n5151), .A3(n5152), .A4(n5153), .ZN(n5140)
         );
  AOI221_X1 U3537 ( .B1(n13045), .B2(n14447), .C1(n13042), .C2(n15850), .A(
        n5157), .ZN(n5150) );
  AOI221_X1 U3538 ( .B1(n13072), .B2(n15810), .C1(n13069), .C2(n15778), .A(
        n5155), .ZN(n5152) );
  AOI221_X1 U3539 ( .B1(n13060), .B2(n14481), .C1(n13057), .C2(n15826), .A(
        n5156), .ZN(n5151) );
  NAND4_X1 U3540 ( .A1(n5113), .A2(n5114), .A3(n5115), .A4(n5116), .ZN(n5103)
         );
  AOI221_X1 U3541 ( .B1(n13046), .B2(n14446), .C1(n13043), .C2(n15849), .A(
        n5120), .ZN(n5113) );
  AOI221_X1 U3542 ( .B1(n13073), .B2(n15809), .C1(n13070), .C2(n15777), .A(
        n5118), .ZN(n5115) );
  AOI221_X1 U3543 ( .B1(n13061), .B2(n14480), .C1(n13058), .C2(n15825), .A(
        n5119), .ZN(n5114) );
  NAND4_X1 U3544 ( .A1(n5076), .A2(n5077), .A3(n5078), .A4(n5079), .ZN(n5066)
         );
  AOI221_X1 U3545 ( .B1(n13046), .B2(n14445), .C1(n13043), .C2(n15848), .A(
        n5083), .ZN(n5076) );
  AOI221_X1 U3546 ( .B1(n13073), .B2(n15808), .C1(n13070), .C2(n15776), .A(
        n5081), .ZN(n5078) );
  AOI221_X1 U3547 ( .B1(n13061), .B2(n14479), .C1(n13058), .C2(n15824), .A(
        n5082), .ZN(n5077) );
  NAND4_X1 U3548 ( .A1(n5039), .A2(n5040), .A3(n5041), .A4(n5042), .ZN(n5029)
         );
  AOI221_X1 U3549 ( .B1(n13046), .B2(n14444), .C1(n13043), .C2(n15847), .A(
        n5046), .ZN(n5039) );
  AOI221_X1 U3550 ( .B1(n13073), .B2(n15807), .C1(n13070), .C2(n15775), .A(
        n5044), .ZN(n5041) );
  AOI221_X1 U3551 ( .B1(n13061), .B2(n14478), .C1(n13058), .C2(n15823), .A(
        n5045), .ZN(n5040) );
  NAND4_X1 U3552 ( .A1(n5002), .A2(n5003), .A3(n5004), .A4(n5005), .ZN(n4992)
         );
  AOI221_X1 U3553 ( .B1(n13046), .B2(n14443), .C1(n13043), .C2(n15846), .A(
        n5009), .ZN(n5002) );
  AOI221_X1 U3554 ( .B1(n13073), .B2(n15806), .C1(n13070), .C2(n15774), .A(
        n5007), .ZN(n5004) );
  AOI221_X1 U3555 ( .B1(n13061), .B2(n14477), .C1(n13058), .C2(n15822), .A(
        n5008), .ZN(n5003) );
  NAND4_X1 U3556 ( .A1(n4965), .A2(n4966), .A3(n4967), .A4(n4968), .ZN(n4955)
         );
  AOI221_X1 U3557 ( .B1(n13046), .B2(n14442), .C1(n13043), .C2(n15845), .A(
        n4972), .ZN(n4965) );
  AOI221_X1 U3558 ( .B1(n13073), .B2(n15805), .C1(n13070), .C2(n15773), .A(
        n4970), .ZN(n4967) );
  AOI221_X1 U3559 ( .B1(n13061), .B2(n14476), .C1(n13058), .C2(n15821), .A(
        n4971), .ZN(n4966) );
  NAND4_X1 U3560 ( .A1(n4928), .A2(n4929), .A3(n4930), .A4(n4931), .ZN(n4918)
         );
  AOI221_X1 U3561 ( .B1(n13046), .B2(n14441), .C1(n13043), .C2(n15844), .A(
        n4935), .ZN(n4928) );
  AOI221_X1 U3562 ( .B1(n13073), .B2(n15804), .C1(n13070), .C2(n15772), .A(
        n4933), .ZN(n4930) );
  AOI221_X1 U3563 ( .B1(n13061), .B2(n14475), .C1(n13058), .C2(n15820), .A(
        n4934), .ZN(n4929) );
  NAND4_X1 U3564 ( .A1(n4891), .A2(n4892), .A3(n4893), .A4(n4894), .ZN(n4881)
         );
  AOI221_X1 U3565 ( .B1(n13046), .B2(n14440), .C1(n13043), .C2(n15843), .A(
        n4898), .ZN(n4891) );
  AOI221_X1 U3566 ( .B1(n13073), .B2(n15803), .C1(n13070), .C2(n15771), .A(
        n4896), .ZN(n4893) );
  AOI221_X1 U3567 ( .B1(n13061), .B2(n14474), .C1(n13058), .C2(n15819), .A(
        n4897), .ZN(n4892) );
  NAND4_X1 U3568 ( .A1(n4854), .A2(n4855), .A3(n4856), .A4(n4857), .ZN(n4844)
         );
  AOI221_X1 U3569 ( .B1(n13046), .B2(n15922), .C1(n13043), .C2(n15842), .A(
        n4861), .ZN(n4854) );
  AOI221_X1 U3570 ( .B1(n13073), .B2(n15802), .C1(n13070), .C2(n15770), .A(
        n4859), .ZN(n4856) );
  AOI221_X1 U3571 ( .B1(n13061), .B2(n14473), .C1(n13058), .C2(n15818), .A(
        n4860), .ZN(n4855) );
  NAND4_X1 U3572 ( .A1(n4817), .A2(n4818), .A3(n4819), .A4(n4820), .ZN(n4807)
         );
  AOI221_X1 U3573 ( .B1(n13046), .B2(n15873), .C1(n13043), .C2(n15841), .A(
        n4824), .ZN(n4817) );
  AOI221_X1 U3574 ( .B1(n13073), .B2(n15801), .C1(n13070), .C2(n15769), .A(
        n4822), .ZN(n4819) );
  AOI221_X1 U3575 ( .B1(n13061), .B2(n14472), .C1(n13058), .C2(n15817), .A(
        n4823), .ZN(n4818) );
  NAND4_X1 U3576 ( .A1(n4780), .A2(n4781), .A3(n4782), .A4(n4783), .ZN(n4770)
         );
  AOI221_X1 U3577 ( .B1(n13046), .B2(n15872), .C1(n13043), .C2(n15840), .A(
        n4787), .ZN(n4780) );
  AOI221_X1 U3578 ( .B1(n13073), .B2(n15800), .C1(n13070), .C2(n15768), .A(
        n4785), .ZN(n4782) );
  AOI221_X1 U3579 ( .B1(n13061), .B2(n14471), .C1(n13058), .C2(n15816), .A(
        n4786), .ZN(n4781) );
  NAND4_X1 U3580 ( .A1(n4743), .A2(n4744), .A3(n4745), .A4(n4746), .ZN(n4733)
         );
  AOI221_X1 U3581 ( .B1(n13046), .B2(n15871), .C1(n13043), .C2(n15839), .A(
        n4750), .ZN(n4743) );
  AOI221_X1 U3582 ( .B1(n13073), .B2(n15799), .C1(n13070), .C2(n15767), .A(
        n4748), .ZN(n4745) );
  AOI221_X1 U3583 ( .B1(n13061), .B2(n14470), .C1(n13058), .C2(n15815), .A(
        n4749), .ZN(n4744) );
  NAND4_X1 U3584 ( .A1(n4706), .A2(n4707), .A3(n4708), .A4(n4709), .ZN(n4696)
         );
  AOI221_X1 U3585 ( .B1(n13046), .B2(n15870), .C1(n13043), .C2(n15838), .A(
        n4713), .ZN(n4706) );
  AOI221_X1 U3586 ( .B1(n13073), .B2(n15798), .C1(n13070), .C2(n15766), .A(
        n4711), .ZN(n4708) );
  AOI221_X1 U3587 ( .B1(n13061), .B2(n14469), .C1(n13058), .C2(n15814), .A(
        n4712), .ZN(n4707) );
  NAND4_X1 U3588 ( .A1(n4669), .A2(n4670), .A3(n4671), .A4(n4672), .ZN(n4659)
         );
  AOI221_X1 U3589 ( .B1(n13047), .B2(n15869), .C1(n13044), .C2(n15632), .A(
        n4676), .ZN(n4669) );
  AOI221_X1 U3590 ( .B1(n13074), .B2(n15797), .C1(n13071), .C2(n15581), .A(
        n4674), .ZN(n4671) );
  AOI221_X1 U3591 ( .B1(n13062), .B2(n14468), .C1(n13059), .C2(n15589), .A(
        n4675), .ZN(n4670) );
  NAND4_X1 U3592 ( .A1(n4284), .A2(n4285), .A3(n4286), .A4(n4287), .ZN(n4263)
         );
  AOI221_X1 U3593 ( .B1(n13273), .B2(n14458), .C1(n13270), .C2(n15861), .A(
        n4293), .ZN(n4284) );
  AOI221_X1 U3594 ( .B1(n13300), .B2(n15789), .C1(n13297), .C2(n14659), .A(
        n4291), .ZN(n4286) );
  AOI221_X1 U3595 ( .B1(n13288), .B2(n14492), .C1(n13285), .C2(n15837), .A(
        n4292), .ZN(n4285) );
  NAND4_X1 U3596 ( .A1(n4236), .A2(n4237), .A3(n4238), .A4(n4239), .ZN(n4226)
         );
  AOI221_X1 U3597 ( .B1(n13273), .B2(n14457), .C1(n13270), .C2(n15860), .A(
        n4243), .ZN(n4236) );
  AOI221_X1 U3598 ( .B1(n13300), .B2(n15788), .C1(n13297), .C2(n14658), .A(
        n4241), .ZN(n4238) );
  AOI221_X1 U3599 ( .B1(n13288), .B2(n14491), .C1(n13285), .C2(n15836), .A(
        n4242), .ZN(n4237) );
  NAND4_X1 U3600 ( .A1(n4199), .A2(n4200), .A3(n4201), .A4(n4202), .ZN(n4189)
         );
  AOI221_X1 U3601 ( .B1(n13273), .B2(n14456), .C1(n13270), .C2(n15859), .A(
        n4206), .ZN(n4199) );
  AOI221_X1 U3602 ( .B1(n13300), .B2(n15787), .C1(n13297), .C2(n14657), .A(
        n4204), .ZN(n4201) );
  AOI221_X1 U3603 ( .B1(n13288), .B2(n14490), .C1(n13285), .C2(n15835), .A(
        n4205), .ZN(n4200) );
  NAND4_X1 U3604 ( .A1(n4162), .A2(n4163), .A3(n4164), .A4(n4165), .ZN(n4152)
         );
  AOI221_X1 U3605 ( .B1(n13273), .B2(n14455), .C1(n13270), .C2(n15858), .A(
        n4169), .ZN(n4162) );
  AOI221_X1 U3606 ( .B1(n13300), .B2(n15786), .C1(n13297), .C2(n14656), .A(
        n4167), .ZN(n4164) );
  AOI221_X1 U3607 ( .B1(n13288), .B2(n14489), .C1(n13285), .C2(n15834), .A(
        n4168), .ZN(n4163) );
  NAND4_X1 U3608 ( .A1(n4125), .A2(n4126), .A3(n4127), .A4(n4128), .ZN(n4115)
         );
  AOI221_X1 U3609 ( .B1(n13273), .B2(n14454), .C1(n13270), .C2(n15857), .A(
        n4132), .ZN(n4125) );
  AOI221_X1 U3610 ( .B1(n13300), .B2(n15785), .C1(n13297), .C2(n14655), .A(
        n4130), .ZN(n4127) );
  AOI221_X1 U3611 ( .B1(n13288), .B2(n14488), .C1(n13285), .C2(n15833), .A(
        n4131), .ZN(n4126) );
  NAND4_X1 U3612 ( .A1(n4088), .A2(n4089), .A3(n4090), .A4(n4091), .ZN(n4078)
         );
  AOI221_X1 U3613 ( .B1(n13273), .B2(n14453), .C1(n13270), .C2(n15856), .A(
        n4095), .ZN(n4088) );
  AOI221_X1 U3614 ( .B1(n13300), .B2(n15784), .C1(n13297), .C2(n14654), .A(
        n4093), .ZN(n4090) );
  AOI221_X1 U3615 ( .B1(n13288), .B2(n14487), .C1(n13285), .C2(n15832), .A(
        n4094), .ZN(n4089) );
  NAND4_X1 U3616 ( .A1(n4051), .A2(n4052), .A3(n4053), .A4(n4054), .ZN(n4041)
         );
  AOI221_X1 U3617 ( .B1(n13273), .B2(n14452), .C1(n13270), .C2(n15855), .A(
        n4058), .ZN(n4051) );
  AOI221_X1 U3618 ( .B1(n13300), .B2(n15783), .C1(n13297), .C2(n14653), .A(
        n4056), .ZN(n4053) );
  AOI221_X1 U3619 ( .B1(n13288), .B2(n14486), .C1(n13285), .C2(n15831), .A(
        n4057), .ZN(n4052) );
  NAND4_X1 U3620 ( .A1(n4014), .A2(n4015), .A3(n4016), .A4(n4017), .ZN(n4004)
         );
  AOI221_X1 U3621 ( .B1(n13273), .B2(n14451), .C1(n13270), .C2(n15854), .A(
        n4021), .ZN(n4014) );
  AOI221_X1 U3622 ( .B1(n13300), .B2(n15782), .C1(n13297), .C2(n15633), .A(
        n4019), .ZN(n4016) );
  AOI221_X1 U3623 ( .B1(n13288), .B2(n14485), .C1(n13285), .C2(n15830), .A(
        n4020), .ZN(n4015) );
  NAND4_X1 U3624 ( .A1(n3977), .A2(n3978), .A3(n3979), .A4(n3980), .ZN(n3967)
         );
  AOI221_X1 U3625 ( .B1(n13273), .B2(n14450), .C1(n13270), .C2(n15853), .A(
        n3984), .ZN(n3977) );
  AOI221_X1 U3626 ( .B1(n13300), .B2(n15781), .C1(n13297), .C2(n15813), .A(
        n3982), .ZN(n3979) );
  AOI221_X1 U3627 ( .B1(n13288), .B2(n14484), .C1(n13285), .C2(n15829), .A(
        n3983), .ZN(n3978) );
  NAND4_X1 U3628 ( .A1(n3940), .A2(n3941), .A3(n3942), .A4(n3943), .ZN(n3930)
         );
  AOI221_X1 U3629 ( .B1(n13273), .B2(n14449), .C1(n13270), .C2(n15852), .A(
        n3947), .ZN(n3940) );
  AOI221_X1 U3630 ( .B1(n13300), .B2(n15780), .C1(n13297), .C2(n15812), .A(
        n3945), .ZN(n3942) );
  AOI221_X1 U3631 ( .B1(n13288), .B2(n14483), .C1(n13285), .C2(n15828), .A(
        n3946), .ZN(n3941) );
  NAND4_X1 U3632 ( .A1(n3903), .A2(n3904), .A3(n3905), .A4(n3906), .ZN(n3893)
         );
  AOI221_X1 U3633 ( .B1(n13273), .B2(n14448), .C1(n13270), .C2(n15851), .A(
        n3910), .ZN(n3903) );
  AOI221_X1 U3634 ( .B1(n13300), .B2(n15779), .C1(n13297), .C2(n15811), .A(
        n3908), .ZN(n3905) );
  AOI221_X1 U3635 ( .B1(n13288), .B2(n14482), .C1(n13285), .C2(n15827), .A(
        n3909), .ZN(n3904) );
  NAND4_X1 U3636 ( .A1(n3866), .A2(n3867), .A3(n3868), .A4(n3869), .ZN(n3856)
         );
  AOI221_X1 U3637 ( .B1(n13273), .B2(n14447), .C1(n13270), .C2(n15850), .A(
        n3873), .ZN(n3866) );
  AOI221_X1 U3638 ( .B1(n13300), .B2(n15778), .C1(n13297), .C2(n15810), .A(
        n3871), .ZN(n3868) );
  AOI221_X1 U3639 ( .B1(n13288), .B2(n14481), .C1(n13285), .C2(n15826), .A(
        n3872), .ZN(n3867) );
  NAND4_X1 U3640 ( .A1(n3829), .A2(n3830), .A3(n3831), .A4(n3832), .ZN(n3819)
         );
  AOI221_X1 U3641 ( .B1(n13274), .B2(n14446), .C1(n13271), .C2(n15849), .A(
        n3836), .ZN(n3829) );
  AOI221_X1 U3642 ( .B1(n13301), .B2(n15777), .C1(n13298), .C2(n15809), .A(
        n3834), .ZN(n3831) );
  AOI221_X1 U3643 ( .B1(n13289), .B2(n14480), .C1(n13286), .C2(n15825), .A(
        n3835), .ZN(n3830) );
  NAND4_X1 U3644 ( .A1(n3792), .A2(n3793), .A3(n3794), .A4(n3795), .ZN(n3782)
         );
  AOI221_X1 U3645 ( .B1(n13274), .B2(n14445), .C1(n13271), .C2(n15848), .A(
        n3799), .ZN(n3792) );
  AOI221_X1 U3646 ( .B1(n13301), .B2(n15776), .C1(n13298), .C2(n15808), .A(
        n3797), .ZN(n3794) );
  AOI221_X1 U3647 ( .B1(n13289), .B2(n14479), .C1(n13286), .C2(n15824), .A(
        n3798), .ZN(n3793) );
  NAND4_X1 U3648 ( .A1(n3755), .A2(n3756), .A3(n3757), .A4(n3758), .ZN(n3745)
         );
  AOI221_X1 U3649 ( .B1(n13274), .B2(n14444), .C1(n13271), .C2(n15847), .A(
        n3762), .ZN(n3755) );
  AOI221_X1 U3650 ( .B1(n13301), .B2(n15775), .C1(n13298), .C2(n15807), .A(
        n3760), .ZN(n3757) );
  AOI221_X1 U3651 ( .B1(n13289), .B2(n14478), .C1(n13286), .C2(n15823), .A(
        n3761), .ZN(n3756) );
  NAND4_X1 U3652 ( .A1(n3718), .A2(n3719), .A3(n3720), .A4(n3721), .ZN(n3708)
         );
  AOI221_X1 U3653 ( .B1(n13274), .B2(n14443), .C1(n13271), .C2(n15846), .A(
        n3725), .ZN(n3718) );
  AOI221_X1 U3654 ( .B1(n13301), .B2(n15774), .C1(n13298), .C2(n15806), .A(
        n3723), .ZN(n3720) );
  AOI221_X1 U3655 ( .B1(n13289), .B2(n14477), .C1(n13286), .C2(n15822), .A(
        n3724), .ZN(n3719) );
  NAND4_X1 U3656 ( .A1(n3681), .A2(n3682), .A3(n3683), .A4(n3684), .ZN(n3671)
         );
  AOI221_X1 U3657 ( .B1(n13274), .B2(n14442), .C1(n13271), .C2(n15845), .A(
        n3688), .ZN(n3681) );
  AOI221_X1 U3658 ( .B1(n13301), .B2(n15773), .C1(n13298), .C2(n15805), .A(
        n3686), .ZN(n3683) );
  AOI221_X1 U3659 ( .B1(n13289), .B2(n14476), .C1(n13286), .C2(n15821), .A(
        n3687), .ZN(n3682) );
  NAND4_X1 U3660 ( .A1(n3644), .A2(n3645), .A3(n3646), .A4(n3647), .ZN(n3634)
         );
  AOI221_X1 U3661 ( .B1(n13274), .B2(n14441), .C1(n13271), .C2(n15844), .A(
        n3651), .ZN(n3644) );
  AOI221_X1 U3662 ( .B1(n13301), .B2(n15772), .C1(n13298), .C2(n15804), .A(
        n3649), .ZN(n3646) );
  AOI221_X1 U3663 ( .B1(n13289), .B2(n14475), .C1(n13286), .C2(n15820), .A(
        n3650), .ZN(n3645) );
  NAND4_X1 U3664 ( .A1(n3607), .A2(n3608), .A3(n3609), .A4(n3610), .ZN(n3597)
         );
  AOI221_X1 U3665 ( .B1(n13274), .B2(n14440), .C1(n13271), .C2(n15843), .A(
        n3614), .ZN(n3607) );
  AOI221_X1 U3666 ( .B1(n13301), .B2(n15771), .C1(n13298), .C2(n15803), .A(
        n3612), .ZN(n3609) );
  AOI221_X1 U3667 ( .B1(n13289), .B2(n14474), .C1(n13286), .C2(n15819), .A(
        n3613), .ZN(n3608) );
  NAND4_X1 U3668 ( .A1(n3570), .A2(n3571), .A3(n3572), .A4(n3573), .ZN(n3560)
         );
  AOI221_X1 U3669 ( .B1(n13274), .B2(n15922), .C1(n13271), .C2(n15842), .A(
        n3577), .ZN(n3570) );
  AOI221_X1 U3670 ( .B1(n13301), .B2(n15770), .C1(n13298), .C2(n15802), .A(
        n3575), .ZN(n3572) );
  AOI221_X1 U3671 ( .B1(n13289), .B2(n14473), .C1(n13286), .C2(n15818), .A(
        n3576), .ZN(n3571) );
  NAND4_X1 U3672 ( .A1(n3533), .A2(n3534), .A3(n3535), .A4(n3536), .ZN(n3523)
         );
  AOI221_X1 U3673 ( .B1(n13274), .B2(n15873), .C1(n13271), .C2(n15841), .A(
        n3540), .ZN(n3533) );
  AOI221_X1 U3674 ( .B1(n13301), .B2(n15769), .C1(n13298), .C2(n15801), .A(
        n3538), .ZN(n3535) );
  AOI221_X1 U3675 ( .B1(n13289), .B2(n14472), .C1(n13286), .C2(n15817), .A(
        n3539), .ZN(n3534) );
  NAND4_X1 U3676 ( .A1(n3496), .A2(n3497), .A3(n3498), .A4(n3499), .ZN(n3486)
         );
  AOI221_X1 U3677 ( .B1(n13274), .B2(n15872), .C1(n13271), .C2(n15840), .A(
        n3503), .ZN(n3496) );
  AOI221_X1 U3678 ( .B1(n13301), .B2(n15768), .C1(n13298), .C2(n15800), .A(
        n3501), .ZN(n3498) );
  AOI221_X1 U3679 ( .B1(n13289), .B2(n14471), .C1(n13286), .C2(n15816), .A(
        n3502), .ZN(n3497) );
  NAND4_X1 U3680 ( .A1(n3459), .A2(n3460), .A3(n3461), .A4(n3462), .ZN(n3449)
         );
  AOI221_X1 U3681 ( .B1(n13274), .B2(n15871), .C1(n13271), .C2(n15839), .A(
        n3466), .ZN(n3459) );
  AOI221_X1 U3682 ( .B1(n13301), .B2(n15767), .C1(n13298), .C2(n15799), .A(
        n3464), .ZN(n3461) );
  AOI221_X1 U3683 ( .B1(n13289), .B2(n14470), .C1(n13286), .C2(n15815), .A(
        n3465), .ZN(n3460) );
  NAND4_X1 U3684 ( .A1(n3422), .A2(n3423), .A3(n3424), .A4(n3425), .ZN(n3412)
         );
  AOI221_X1 U3685 ( .B1(n13274), .B2(n15870), .C1(n13271), .C2(n15838), .A(
        n3429), .ZN(n3422) );
  AOI221_X1 U3686 ( .B1(n13301), .B2(n15766), .C1(n13298), .C2(n15798), .A(
        n3427), .ZN(n3424) );
  AOI221_X1 U3687 ( .B1(n13289), .B2(n14469), .C1(n13286), .C2(n15814), .A(
        n3428), .ZN(n3423) );
  NAND4_X1 U3688 ( .A1(n3385), .A2(n3386), .A3(n3387), .A4(n3388), .ZN(n3375)
         );
  AOI221_X1 U3689 ( .B1(n13275), .B2(n15869), .C1(n13272), .C2(n15632), .A(
        n3392), .ZN(n3385) );
  AOI221_X1 U3690 ( .B1(n13302), .B2(n15581), .C1(n13299), .C2(n15797), .A(
        n3390), .ZN(n3387) );
  AOI221_X1 U3691 ( .B1(n13290), .B2(n14468), .C1(n13287), .C2(n15589), .A(
        n3391), .ZN(n3386) );
  NAND4_X1 U3692 ( .A1(n3348), .A2(n3349), .A3(n3350), .A4(n3351), .ZN(n3338)
         );
  AOI221_X1 U3693 ( .B1(n13275), .B2(n15868), .C1(n13272), .C2(n15631), .A(
        n3355), .ZN(n3348) );
  AOI221_X1 U3694 ( .B1(n13302), .B2(n15580), .C1(n13299), .C2(n15796), .A(
        n3353), .ZN(n3350) );
  AOI221_X1 U3695 ( .B1(n13290), .B2(n14467), .C1(n13287), .C2(n15588), .A(
        n3354), .ZN(n3349) );
  NAND4_X1 U3696 ( .A1(n3311), .A2(n3312), .A3(n3313), .A4(n3314), .ZN(n3301)
         );
  AOI221_X1 U3697 ( .B1(n13275), .B2(n15867), .C1(n13272), .C2(n15630), .A(
        n3318), .ZN(n3311) );
  AOI221_X1 U3698 ( .B1(n13302), .B2(n15579), .C1(n13299), .C2(n15795), .A(
        n3316), .ZN(n3313) );
  AOI221_X1 U3699 ( .B1(n13290), .B2(n14466), .C1(n13287), .C2(n15587), .A(
        n3317), .ZN(n3312) );
  NAND4_X1 U3700 ( .A1(n3274), .A2(n3275), .A3(n3276), .A4(n3277), .ZN(n3264)
         );
  AOI221_X1 U3701 ( .B1(n13275), .B2(n15866), .C1(n13272), .C2(n15629), .A(
        n3281), .ZN(n3274) );
  AOI221_X1 U3702 ( .B1(n13302), .B2(n15578), .C1(n13299), .C2(n15794), .A(
        n3279), .ZN(n3276) );
  AOI221_X1 U3703 ( .B1(n13290), .B2(n14465), .C1(n13287), .C2(n15586), .A(
        n3280), .ZN(n3275) );
  NOR3_X2 U3704 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[1]), .A3(n16066), .ZN(n4278) );
  NOR3_X2 U3705 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[2]), .A3(n16068), .ZN(n5671) );
  NOR3_X2 U3706 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n16067), .ZN(n5666) );
  NOR3_X2 U3707 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[2]), .A3(n16065), .ZN(n4280) );
  NOR3_X2 U3708 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[1]), .A3(n16069), .ZN(n5674) );
  NOR3_X2 U3709 ( .A1(n16067), .A2(ADD_RD2[2]), .A3(n16068), .ZN(n5676) );
  BUF_X1 U3710 ( .A(n16063), .Z(n12922) );
  BUF_X1 U3711 ( .A(n16063), .Z(n12923) );
  BUF_X1 U3712 ( .A(n16063), .Z(n12924) );
  BUF_X1 U3713 ( .A(n16063), .Z(n12925) );
  BUF_X1 U3714 ( .A(n16063), .Z(n12926) );
  BUF_X1 U3715 ( .A(n16063), .Z(n12927) );
  INV_X1 U3716 ( .A(ADD_RD2[0]), .ZN(n16067) );
  INV_X1 U3717 ( .A(ADD_RD1[0]), .ZN(n16064) );
  BUF_X1 U3718 ( .A(n2864), .Z(n13830) );
  BUF_X1 U3719 ( .A(n2863), .Z(n13836) );
  BUF_X1 U3720 ( .A(n2862), .Z(n13842) );
  BUF_X1 U3721 ( .A(n2861), .Z(n13848) );
  BUF_X1 U3722 ( .A(n2860), .Z(n13854) );
  BUF_X1 U3723 ( .A(n2859), .Z(n13860) );
  BUF_X1 U3724 ( .A(n2858), .Z(n13866) );
  BUF_X1 U3725 ( .A(n2857), .Z(n13872) );
  BUF_X1 U3726 ( .A(n2856), .Z(n13878) );
  BUF_X1 U3727 ( .A(n2855), .Z(n13884) );
  BUF_X1 U3728 ( .A(n2854), .Z(n13890) );
  BUF_X1 U3729 ( .A(n2853), .Z(n13896) );
  BUF_X1 U3730 ( .A(n2852), .Z(n13902) );
  BUF_X1 U3731 ( .A(n2851), .Z(n13908) );
  BUF_X1 U3732 ( .A(n2850), .Z(n13914) );
  BUF_X1 U3733 ( .A(n2849), .Z(n13920) );
  BUF_X1 U3734 ( .A(n2848), .Z(n13926) );
  BUF_X1 U3735 ( .A(n2847), .Z(n13932) );
  BUF_X1 U3736 ( .A(n2846), .Z(n13938) );
  BUF_X1 U3737 ( .A(n2845), .Z(n13944) );
  BUF_X1 U3738 ( .A(n2844), .Z(n13950) );
  BUF_X1 U3739 ( .A(n2843), .Z(n13956) );
  BUF_X1 U3740 ( .A(n2842), .Z(n13962) );
  BUF_X1 U3741 ( .A(n2841), .Z(n13968) );
  BUF_X1 U3742 ( .A(n2840), .Z(n13974) );
  BUF_X1 U3743 ( .A(n2839), .Z(n13980) );
  BUF_X1 U3744 ( .A(n2838), .Z(n13986) );
  BUF_X1 U3745 ( .A(n2837), .Z(n13992) );
  BUF_X1 U3746 ( .A(n2836), .Z(n13998) );
  BUF_X1 U3747 ( .A(n2835), .Z(n14004) );
  BUF_X1 U3748 ( .A(n2833), .Z(n14013) );
  BUF_X1 U3749 ( .A(n2865), .Z(n13824) );
  BUF_X1 U3750 ( .A(n2865), .Z(n13828) );
  BUF_X1 U3751 ( .A(n2864), .Z(n13834) );
  BUF_X1 U3752 ( .A(n2863), .Z(n13840) );
  BUF_X1 U3753 ( .A(n2862), .Z(n13846) );
  BUF_X1 U3754 ( .A(n2861), .Z(n13852) );
  BUF_X1 U3755 ( .A(n2860), .Z(n13858) );
  BUF_X1 U3756 ( .A(n2859), .Z(n13864) );
  BUF_X1 U3757 ( .A(n2858), .Z(n13870) );
  BUF_X1 U3758 ( .A(n2857), .Z(n13876) );
  BUF_X1 U3759 ( .A(n2856), .Z(n13882) );
  BUF_X1 U3760 ( .A(n2855), .Z(n13888) );
  BUF_X1 U3761 ( .A(n2854), .Z(n13894) );
  BUF_X1 U3762 ( .A(n2853), .Z(n13900) );
  BUF_X1 U3763 ( .A(n2852), .Z(n13906) );
  BUF_X1 U3764 ( .A(n2851), .Z(n13912) );
  BUF_X1 U3765 ( .A(n2850), .Z(n13918) );
  BUF_X1 U3766 ( .A(n2849), .Z(n13924) );
  BUF_X1 U3767 ( .A(n2848), .Z(n13930) );
  BUF_X1 U3768 ( .A(n2847), .Z(n13936) );
  BUF_X1 U3769 ( .A(n2846), .Z(n13942) );
  BUF_X1 U3770 ( .A(n2845), .Z(n13948) );
  BUF_X1 U3771 ( .A(n2844), .Z(n13954) );
  BUF_X1 U3772 ( .A(n2843), .Z(n13960) );
  BUF_X1 U3773 ( .A(n2842), .Z(n13966) );
  BUF_X1 U3774 ( .A(n2841), .Z(n13972) );
  BUF_X1 U3775 ( .A(n2840), .Z(n13978) );
  BUF_X1 U3776 ( .A(n2839), .Z(n13984) );
  BUF_X1 U3777 ( .A(n2838), .Z(n13990) );
  BUF_X1 U3778 ( .A(n2837), .Z(n13996) );
  BUF_X1 U3779 ( .A(n2836), .Z(n14002) );
  BUF_X1 U3780 ( .A(n2835), .Z(n14008) );
  BUF_X1 U3781 ( .A(n2833), .Z(n14017) );
  BUF_X1 U3782 ( .A(n2865), .Z(n13827) );
  BUF_X1 U3783 ( .A(n2864), .Z(n13833) );
  BUF_X1 U3784 ( .A(n2863), .Z(n13839) );
  BUF_X1 U3785 ( .A(n2862), .Z(n13845) );
  BUF_X1 U3786 ( .A(n2861), .Z(n13851) );
  BUF_X1 U3787 ( .A(n2860), .Z(n13857) );
  BUF_X1 U3788 ( .A(n2859), .Z(n13863) );
  BUF_X1 U3789 ( .A(n2858), .Z(n13869) );
  BUF_X1 U3790 ( .A(n2857), .Z(n13875) );
  BUF_X1 U3791 ( .A(n2856), .Z(n13881) );
  BUF_X1 U3792 ( .A(n2855), .Z(n13887) );
  BUF_X1 U3793 ( .A(n2854), .Z(n13893) );
  BUF_X1 U3794 ( .A(n2853), .Z(n13899) );
  BUF_X1 U3795 ( .A(n2852), .Z(n13905) );
  BUF_X1 U3796 ( .A(n2851), .Z(n13911) );
  BUF_X1 U3797 ( .A(n2850), .Z(n13917) );
  BUF_X1 U3798 ( .A(n2849), .Z(n13923) );
  BUF_X1 U3799 ( .A(n2848), .Z(n13929) );
  BUF_X1 U3800 ( .A(n2847), .Z(n13935) );
  BUF_X1 U3801 ( .A(n2846), .Z(n13941) );
  BUF_X1 U3802 ( .A(n2845), .Z(n13947) );
  BUF_X1 U3803 ( .A(n2844), .Z(n13953) );
  BUF_X1 U3804 ( .A(n2843), .Z(n13959) );
  BUF_X1 U3805 ( .A(n2842), .Z(n13965) );
  BUF_X1 U3806 ( .A(n2841), .Z(n13971) );
  BUF_X1 U3807 ( .A(n2840), .Z(n13977) );
  BUF_X1 U3808 ( .A(n2839), .Z(n13983) );
  BUF_X1 U3809 ( .A(n2838), .Z(n13989) );
  BUF_X1 U3810 ( .A(n2837), .Z(n13995) );
  BUF_X1 U3811 ( .A(n2836), .Z(n14001) );
  BUF_X1 U3812 ( .A(n2835), .Z(n14007) );
  BUF_X1 U3813 ( .A(n2833), .Z(n14016) );
  BUF_X1 U3814 ( .A(n2865), .Z(n13826) );
  BUF_X1 U3815 ( .A(n2864), .Z(n13832) );
  BUF_X1 U3816 ( .A(n2863), .Z(n13838) );
  BUF_X1 U3818 ( .A(n2862), .Z(n13844) );
  BUF_X1 U3819 ( .A(n2861), .Z(n13850) );
  BUF_X1 U3820 ( .A(n2860), .Z(n13856) );
  BUF_X1 U3821 ( .A(n2859), .Z(n13862) );
  BUF_X1 U3822 ( .A(n2858), .Z(n13868) );
  BUF_X1 U3823 ( .A(n2857), .Z(n13874) );
  BUF_X1 U3824 ( .A(n2856), .Z(n13880) );
  BUF_X1 U3825 ( .A(n2855), .Z(n13886) );
  BUF_X1 U3826 ( .A(n2854), .Z(n13892) );
  BUF_X1 U3827 ( .A(n2853), .Z(n13898) );
  BUF_X1 U3828 ( .A(n2852), .Z(n13904) );
  BUF_X1 U3829 ( .A(n2851), .Z(n13910) );
  BUF_X1 U3830 ( .A(n2850), .Z(n13916) );
  BUF_X1 U3831 ( .A(n2849), .Z(n13922) );
  BUF_X1 U3832 ( .A(n2848), .Z(n13928) );
  BUF_X1 U3833 ( .A(n2847), .Z(n13934) );
  BUF_X1 U3834 ( .A(n2846), .Z(n13940) );
  BUF_X1 U3835 ( .A(n2845), .Z(n13946) );
  BUF_X1 U3836 ( .A(n2844), .Z(n13952) );
  BUF_X1 U3837 ( .A(n2843), .Z(n13958) );
  BUF_X1 U3838 ( .A(n2842), .Z(n13964) );
  BUF_X1 U3839 ( .A(n2841), .Z(n13970) );
  BUF_X1 U3840 ( .A(n2840), .Z(n13976) );
  BUF_X1 U3841 ( .A(n2839), .Z(n13982) );
  BUF_X1 U3842 ( .A(n2838), .Z(n13988) );
  BUF_X1 U3843 ( .A(n2837), .Z(n13994) );
  BUF_X1 U3844 ( .A(n2836), .Z(n14000) );
  BUF_X1 U3845 ( .A(n2835), .Z(n14006) );
  BUF_X1 U3846 ( .A(n2833), .Z(n14015) );
  BUF_X1 U3847 ( .A(n2865), .Z(n13825) );
  BUF_X1 U3848 ( .A(n2864), .Z(n13831) );
  BUF_X1 U3849 ( .A(n2863), .Z(n13837) );
  BUF_X1 U3850 ( .A(n2862), .Z(n13843) );
  BUF_X1 U3851 ( .A(n2861), .Z(n13849) );
  BUF_X1 U3852 ( .A(n2860), .Z(n13855) );
  BUF_X1 U3853 ( .A(n2859), .Z(n13861) );
  BUF_X1 U3854 ( .A(n2858), .Z(n13867) );
  BUF_X1 U3855 ( .A(n2857), .Z(n13873) );
  BUF_X1 U3856 ( .A(n2856), .Z(n13879) );
  BUF_X1 U3857 ( .A(n2855), .Z(n13885) );
  BUF_X1 U3858 ( .A(n2854), .Z(n13891) );
  BUF_X1 U3859 ( .A(n2853), .Z(n13897) );
  BUF_X1 U3860 ( .A(n2852), .Z(n13903) );
  BUF_X1 U3861 ( .A(n2851), .Z(n13909) );
  BUF_X1 U3862 ( .A(n2850), .Z(n13915) );
  BUF_X1 U3863 ( .A(n2849), .Z(n13921) );
  BUF_X1 U3864 ( .A(n2848), .Z(n13927) );
  BUF_X1 U3865 ( .A(n2847), .Z(n13933) );
  BUF_X1 U3866 ( .A(n2846), .Z(n13939) );
  BUF_X1 U3867 ( .A(n2845), .Z(n13945) );
  BUF_X1 U3868 ( .A(n2844), .Z(n13951) );
  BUF_X1 U3869 ( .A(n2843), .Z(n13957) );
  BUF_X1 U3870 ( .A(n2842), .Z(n13963) );
  BUF_X1 U3871 ( .A(n2841), .Z(n13969) );
  BUF_X1 U3872 ( .A(n2840), .Z(n13975) );
  BUF_X1 U3873 ( .A(n2839), .Z(n13981) );
  BUF_X1 U3874 ( .A(n2838), .Z(n13987) );
  BUF_X1 U3875 ( .A(n2837), .Z(n13993) );
  BUF_X1 U3876 ( .A(n2836), .Z(n13999) );
  BUF_X1 U3877 ( .A(n2835), .Z(n14005) );
  BUF_X1 U3878 ( .A(n2833), .Z(n14014) );
  INV_X1 U3879 ( .A(ADD_RD2[1]), .ZN(n16068) );
  INV_X1 U3880 ( .A(ADD_RD1[1]), .ZN(n16065) );
  INV_X1 U3881 ( .A(ADD_RD2[2]), .ZN(n16069) );
  INV_X1 U3882 ( .A(ADD_RD1[2]), .ZN(n16066) );
  NAND2_X1 U3883 ( .A1(n14027), .A2(n16074), .ZN(n4325) );
  NAND2_X1 U3884 ( .A1(n14027), .A2(n16073), .ZN(n3041) );
  NAND4_X1 U3885 ( .A1(n5738), .A2(n5740), .A3(n5742), .A4(n5744), .ZN(n4322)
         );
  NOR3_X1 U3886 ( .A1(n5754), .A2(n16075), .A3(n16074), .ZN(n5742) );
  NAND4_X1 U3887 ( .A1(n4313), .A2(n4314), .A3(n4315), .A4(n4316), .ZN(n3038)
         );
  NOR3_X1 U3888 ( .A1(n4321), .A2(n16075), .A3(n16073), .ZN(n4315) );
  NOR2_X1 U3889 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .ZN(n3000) );
  NOR2_X1 U3890 ( .A1(n16070), .A2(ADD_WR[1]), .ZN(n3003) );
  NOR2_X1 U3891 ( .A1(n16071), .A2(ADD_WR[0]), .ZN(n3006) );
  NOR2_X1 U3892 ( .A1(ADD_WR[2]), .A2(ADD_WR[3]), .ZN(n3022) );
  INV_X1 U3893 ( .A(ADD_WR[1]), .ZN(n16071) );
  INV_X1 U3894 ( .A(ADD_WR[2]), .ZN(n16072) );
  AND2_X1 U3895 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .ZN(n3012) );
  INV_X1 U3896 ( .A(ADD_WR[0]), .ZN(n16070) );
  INV_X1 U3897 ( .A(n13810), .ZN(n13823) );
  AOI221_X1 U3898 ( .B1(n13182), .B2(n5982), .C1(n13179), .C2(n15177), .A(
        n3259), .ZN(n3254) );
  OAI222_X1 U3899 ( .A1(n15273), .A2(n13176), .B1(n15209), .B2(n13173), .C1(
        n15241), .C2(n13170), .ZN(n3259) );
  AOI221_X1 U3900 ( .B1(n13182), .B2(n5983), .C1(n13179), .C2(n15176), .A(
        n3222), .ZN(n3217) );
  OAI222_X1 U3901 ( .A1(n15272), .A2(n13176), .B1(n15208), .B2(n13173), .C1(
        n15240), .C2(n13170), .ZN(n3222) );
  AOI221_X1 U3902 ( .B1(n13182), .B2(n5984), .C1(n13179), .C2(n15175), .A(
        n3185), .ZN(n3180) );
  OAI222_X1 U3903 ( .A1(n15271), .A2(n13176), .B1(n15207), .B2(n13173), .C1(
        n15239), .C2(n13170), .ZN(n3185) );
  AOI221_X1 U3904 ( .B1(n13182), .B2(n5985), .C1(n13179), .C2(n15174), .A(
        n3141), .ZN(n3125) );
  OAI222_X1 U3905 ( .A1(n15270), .A2(n13176), .B1(n15206), .B2(n13173), .C1(
        n15238), .C2(n13170), .ZN(n3141) );
  AOI221_X1 U3906 ( .B1(n12954), .B2(n5979), .C1(n12951), .C2(n15180), .A(
        n4654), .ZN(n4649) );
  OAI222_X1 U3907 ( .A1(n15276), .A2(n12948), .B1(n15212), .B2(n12945), .C1(
        n15244), .C2(n12942), .ZN(n4654) );
  AOI221_X1 U3908 ( .B1(n12954), .B2(n5980), .C1(n12951), .C2(n15179), .A(
        n4617), .ZN(n4612) );
  OAI222_X1 U3909 ( .A1(n15275), .A2(n12948), .B1(n15211), .B2(n12945), .C1(
        n15243), .C2(n12942), .ZN(n4617) );
  AOI221_X1 U3910 ( .B1(n12954), .B2(n5981), .C1(n12951), .C2(n15178), .A(
        n4580), .ZN(n4575) );
  OAI222_X1 U3911 ( .A1(n15274), .A2(n12948), .B1(n15210), .B2(n12945), .C1(
        n15242), .C2(n12942), .ZN(n4580) );
  AOI221_X1 U3912 ( .B1(n12954), .B2(n5982), .C1(n12951), .C2(n15177), .A(
        n4543), .ZN(n4538) );
  OAI222_X1 U3913 ( .A1(n15273), .A2(n12948), .B1(n15209), .B2(n12945), .C1(
        n15241), .C2(n12942), .ZN(n4543) );
  AOI221_X1 U3914 ( .B1(n12954), .B2(n5983), .C1(n12951), .C2(n15176), .A(
        n4506), .ZN(n4501) );
  OAI222_X1 U3915 ( .A1(n15272), .A2(n12948), .B1(n15208), .B2(n12945), .C1(
        n15240), .C2(n12942), .ZN(n4506) );
  AOI221_X1 U3916 ( .B1(n12954), .B2(n5984), .C1(n12951), .C2(n15175), .A(
        n4469), .ZN(n4464) );
  OAI222_X1 U3917 ( .A1(n15271), .A2(n12948), .B1(n15207), .B2(n12945), .C1(
        n15239), .C2(n12942), .ZN(n4469) );
  AOI221_X1 U3918 ( .B1(n12954), .B2(n5985), .C1(n12951), .C2(n15174), .A(
        n4425), .ZN(n4409) );
  OAI222_X1 U3919 ( .A1(n15270), .A2(n12948), .B1(n15206), .B2(n12945), .C1(
        n15238), .C2(n12942), .ZN(n4425) );
  AOI221_X1 U3920 ( .B1(n13008), .B2(n6234), .C1(n13005), .C2(n15565), .A(
        n4683), .ZN(n4678) );
  OAI222_X1 U3921 ( .A1(n14923), .A2(n13002), .B1(n14859), .B2(n12999), .C1(
        n14891), .C2(n12996), .ZN(n4683) );
  AOI221_X1 U3922 ( .B1(n13236), .B2(n6234), .C1(n13233), .C2(n15565), .A(
        n3399), .ZN(n3394) );
  OAI222_X1 U3923 ( .A1(n14923), .A2(n13230), .B1(n14859), .B2(n13227), .C1(
        n14891), .C2(n13224), .ZN(n3399) );
  AOI221_X1 U3924 ( .B1(n13182), .B2(n5979), .C1(n13179), .C2(n15180), .A(
        n3370), .ZN(n3365) );
  OAI222_X1 U3925 ( .A1(n15276), .A2(n13176), .B1(n15212), .B2(n13173), .C1(
        n15244), .C2(n13170), .ZN(n3370) );
  AOI221_X1 U3926 ( .B1(n13182), .B2(n5980), .C1(n13179), .C2(n15179), .A(
        n3333), .ZN(n3328) );
  OAI222_X1 U3927 ( .A1(n15275), .A2(n13176), .B1(n15211), .B2(n13173), .C1(
        n15243), .C2(n13170), .ZN(n3333) );
  AOI221_X1 U3928 ( .B1(n13182), .B2(n5981), .C1(n13179), .C2(n15178), .A(
        n3296), .ZN(n3291) );
  OAI222_X1 U3929 ( .A1(n15274), .A2(n13176), .B1(n15210), .B2(n13173), .C1(
        n15242), .C2(n13170), .ZN(n3296) );
  OAI222_X1 U3930 ( .A1(n16082), .A2(n13155), .B1(n4619), .B2(n13152), .C1(
        n13144), .C2(n1487), .ZN(n7597) );
  NOR4_X1 U3931 ( .A1(n4620), .A2(n4621), .A3(n4622), .A4(n4623), .ZN(n4619)
         );
  NAND4_X1 U3932 ( .A1(n4648), .A2(n4649), .A3(n4650), .A4(n4651), .ZN(n4620)
         );
  NAND4_X1 U3933 ( .A1(n4640), .A2(n4641), .A3(n4642), .A4(n4643), .ZN(n4621)
         );
  OAI222_X1 U3934 ( .A1(n16081), .A2(n13155), .B1(n4582), .B2(n13152), .C1(
        n13144), .C2(n1486), .ZN(n7599) );
  NOR4_X1 U3935 ( .A1(n4583), .A2(n4584), .A3(n4585), .A4(n4586), .ZN(n4582)
         );
  NAND4_X1 U3936 ( .A1(n4611), .A2(n4612), .A3(n4613), .A4(n4614), .ZN(n4583)
         );
  NAND4_X1 U3937 ( .A1(n4603), .A2(n4604), .A3(n4605), .A4(n4606), .ZN(n4584)
         );
  OAI222_X1 U3938 ( .A1(n16080), .A2(n13155), .B1(n4545), .B2(n13152), .C1(
        n13144), .C2(n1485), .ZN(n7601) );
  NOR4_X1 U3939 ( .A1(n4546), .A2(n4547), .A3(n4548), .A4(n4549), .ZN(n4545)
         );
  NAND4_X1 U3940 ( .A1(n4574), .A2(n4575), .A3(n4576), .A4(n4577), .ZN(n4546)
         );
  NAND4_X1 U3941 ( .A1(n4566), .A2(n4567), .A3(n4568), .A4(n4569), .ZN(n4547)
         );
  OAI222_X1 U3942 ( .A1(n16079), .A2(n13155), .B1(n4508), .B2(n13152), .C1(
        n13144), .C2(n1484), .ZN(n7603) );
  NOR4_X1 U3943 ( .A1(n4509), .A2(n4510), .A3(n4511), .A4(n4512), .ZN(n4508)
         );
  NAND4_X1 U3944 ( .A1(n4537), .A2(n4538), .A3(n4539), .A4(n4540), .ZN(n4509)
         );
  NAND4_X1 U3945 ( .A1(n4529), .A2(n4530), .A3(n4531), .A4(n4532), .ZN(n4510)
         );
  OAI222_X1 U3946 ( .A1(n16078), .A2(n13155), .B1(n4471), .B2(n13152), .C1(
        n13144), .C2(n1483), .ZN(n7605) );
  NOR4_X1 U3947 ( .A1(n4472), .A2(n4473), .A3(n4474), .A4(n4475), .ZN(n4471)
         );
  NAND4_X1 U3948 ( .A1(n4500), .A2(n4501), .A3(n4502), .A4(n4503), .ZN(n4472)
         );
  NAND4_X1 U3949 ( .A1(n4492), .A2(n4493), .A3(n4494), .A4(n4495), .ZN(n4473)
         );
  OAI222_X1 U3950 ( .A1(n16077), .A2(n13155), .B1(n4434), .B2(n13152), .C1(
        n13144), .C2(n1482), .ZN(n7607) );
  NOR4_X1 U3951 ( .A1(n4435), .A2(n4436), .A3(n4437), .A4(n4438), .ZN(n4434)
         );
  NAND4_X1 U3952 ( .A1(n4463), .A2(n4464), .A3(n4465), .A4(n4466), .ZN(n4435)
         );
  NAND4_X1 U3953 ( .A1(n4455), .A2(n4456), .A3(n4457), .A4(n4458), .ZN(n4436)
         );
  OAI222_X1 U3954 ( .A1(n16076), .A2(n13155), .B1(n4323), .B2(n13152), .C1(
        n13145), .C2(n1481), .ZN(n7609) );
  NOR4_X1 U3955 ( .A1(n4326), .A2(n4327), .A3(n4328), .A4(n4329), .ZN(n4323)
         );
  NAND4_X1 U3956 ( .A1(n4408), .A2(n4409), .A3(n4410), .A4(n4411), .ZN(n4326)
         );
  NAND4_X1 U3957 ( .A1(n4382), .A2(n4383), .A3(n4384), .A4(n4385), .ZN(n4327)
         );
  AOI221_X1 U3958 ( .B1(n13248), .B2(n6174), .C1(n13245), .C2(n15615), .A(
        n3250), .ZN(n3247) );
  OAI22_X1 U3959 ( .A1(n14952), .A2(n13242), .B1(n15926), .B2(n13239), .ZN(
        n3250) );
  AOI221_X1 U3960 ( .B1(n13194), .B2(n5918), .C1(n13191), .C2(n15305), .A(
        n3258), .ZN(n3255) );
  OAI22_X1 U3961 ( .A1(n15337), .A2(n13188), .B1(n15369), .B2(n13185), .ZN(
        n3258) );
  AOI221_X1 U3962 ( .B1(n13248), .B2(n6175), .C1(n13245), .C2(n15614), .A(
        n3213), .ZN(n3210) );
  OAI22_X1 U3963 ( .A1(n14951), .A2(n13242), .B1(n15925), .B2(n13239), .ZN(
        n3213) );
  AOI221_X1 U3964 ( .B1(n13194), .B2(n5919), .C1(n13191), .C2(n15304), .A(
        n3221), .ZN(n3218) );
  OAI22_X1 U3965 ( .A1(n15336), .A2(n13188), .B1(n15368), .B2(n13185), .ZN(
        n3221) );
  AOI221_X1 U3966 ( .B1(n13248), .B2(n6176), .C1(n13245), .C2(n15613), .A(
        n3176), .ZN(n3173) );
  OAI22_X1 U3967 ( .A1(n14950), .A2(n13242), .B1(n15924), .B2(n13239), .ZN(
        n3176) );
  AOI221_X1 U3968 ( .B1(n13194), .B2(n5920), .C1(n13191), .C2(n15303), .A(
        n3184), .ZN(n3181) );
  OAI22_X1 U3969 ( .A1(n15335), .A2(n13188), .B1(n15367), .B2(n13185), .ZN(
        n3184) );
  AOI221_X1 U3970 ( .B1(n13248), .B2(n6177), .C1(n13245), .C2(n14948), .A(
        n3110), .ZN(n3100) );
  OAI22_X1 U3971 ( .A1(n14949), .A2(n13242), .B1(n15923), .B2(n13239), .ZN(
        n3110) );
  AOI221_X1 U3972 ( .B1(n13194), .B2(n5921), .C1(n13191), .C2(n15302), .A(
        n3136), .ZN(n3126) );
  OAI22_X1 U3973 ( .A1(n15334), .A2(n13188), .B1(n15366), .B2(n13185), .ZN(
        n3136) );
  AOI221_X1 U3974 ( .B1(n13020), .B2(n6171), .C1(n13017), .C2(n15618), .A(
        n4645), .ZN(n4642) );
  OAI22_X1 U3975 ( .A1(n14955), .A2(n13014), .B1(n15929), .B2(n13011), .ZN(
        n4645) );
  AOI221_X1 U3976 ( .B1(n12966), .B2(n5915), .C1(n12963), .C2(n15308), .A(
        n4653), .ZN(n4650) );
  OAI22_X1 U3977 ( .A1(n15340), .A2(n12960), .B1(n15372), .B2(n12957), .ZN(
        n4653) );
  AOI221_X1 U3978 ( .B1(n13020), .B2(n6172), .C1(n13017), .C2(n15617), .A(
        n4608), .ZN(n4605) );
  OAI22_X1 U3979 ( .A1(n14954), .A2(n13014), .B1(n15928), .B2(n13011), .ZN(
        n4608) );
  AOI221_X1 U3980 ( .B1(n12966), .B2(n5916), .C1(n12963), .C2(n15307), .A(
        n4616), .ZN(n4613) );
  OAI22_X1 U3981 ( .A1(n15339), .A2(n12960), .B1(n15371), .B2(n12957), .ZN(
        n4616) );
  AOI221_X1 U3982 ( .B1(n13020), .B2(n6173), .C1(n13017), .C2(n15616), .A(
        n4571), .ZN(n4568) );
  OAI22_X1 U3983 ( .A1(n14953), .A2(n13014), .B1(n15927), .B2(n13011), .ZN(
        n4571) );
  AOI221_X1 U3984 ( .B1(n12966), .B2(n5917), .C1(n12963), .C2(n15306), .A(
        n4579), .ZN(n4576) );
  OAI22_X1 U3985 ( .A1(n15338), .A2(n12960), .B1(n15370), .B2(n12957), .ZN(
        n4579) );
  AOI221_X1 U3986 ( .B1(n13020), .B2(n6174), .C1(n13017), .C2(n15615), .A(
        n4534), .ZN(n4531) );
  OAI22_X1 U3987 ( .A1(n14952), .A2(n13014), .B1(n15926), .B2(n13011), .ZN(
        n4534) );
  AOI221_X1 U3988 ( .B1(n12966), .B2(n5918), .C1(n12963), .C2(n15305), .A(
        n4542), .ZN(n4539) );
  OAI22_X1 U3989 ( .A1(n15337), .A2(n12960), .B1(n15369), .B2(n12957), .ZN(
        n4542) );
  AOI221_X1 U3990 ( .B1(n13020), .B2(n6175), .C1(n13017), .C2(n15614), .A(
        n4497), .ZN(n4494) );
  OAI22_X1 U3991 ( .A1(n14951), .A2(n13014), .B1(n15925), .B2(n13011), .ZN(
        n4497) );
  AOI221_X1 U3992 ( .B1(n12966), .B2(n5919), .C1(n12963), .C2(n15304), .A(
        n4505), .ZN(n4502) );
  OAI22_X1 U3993 ( .A1(n15336), .A2(n12960), .B1(n15368), .B2(n12957), .ZN(
        n4505) );
  AOI221_X1 U3994 ( .B1(n13020), .B2(n6176), .C1(n13017), .C2(n15613), .A(
        n4460), .ZN(n4457) );
  OAI22_X1 U3995 ( .A1(n14950), .A2(n13014), .B1(n15924), .B2(n13011), .ZN(
        n4460) );
  AOI221_X1 U3996 ( .B1(n12966), .B2(n5920), .C1(n12963), .C2(n15303), .A(
        n4468), .ZN(n4465) );
  OAI22_X1 U3997 ( .A1(n15335), .A2(n12960), .B1(n15367), .B2(n12957), .ZN(
        n4468) );
  AOI221_X1 U3998 ( .B1(n13020), .B2(n6177), .C1(n13017), .C2(n14948), .A(
        n4394), .ZN(n4384) );
  OAI22_X1 U3999 ( .A1(n14949), .A2(n13014), .B1(n15923), .B2(n13011), .ZN(
        n4394) );
  AOI221_X1 U4000 ( .B1(n12966), .B2(n5921), .C1(n12963), .C2(n15302), .A(
        n4420), .ZN(n4410) );
  OAI22_X1 U4001 ( .A1(n15334), .A2(n12960), .B1(n15366), .B2(n12957), .ZN(
        n4420) );
  AOI221_X1 U4002 ( .B1(n13018), .B2(n6146), .C1(n13015), .C2(n15681), .A(
        n5712), .ZN(n5704) );
  OAI22_X1 U4003 ( .A1(n14980), .A2(n13012), .B1(n15970), .B2(n13009), .ZN(
        n5712) );
  AOI221_X1 U4004 ( .B1(n12964), .B2(n5890), .C1(n12961), .C2(n15333), .A(
        n5730), .ZN(n5724) );
  OAI22_X1 U4005 ( .A1(n15365), .A2(n12958), .B1(n15397), .B2(n12955), .ZN(
        n5730) );
  AOI221_X1 U4006 ( .B1(n13018), .B2(n6147), .C1(n13015), .C2(n15680), .A(
        n5624), .ZN(n5619) );
  OAI22_X1 U4007 ( .A1(n14979), .A2(n13012), .B1(n15969), .B2(n13009), .ZN(
        n5624) );
  AOI221_X1 U4008 ( .B1(n12964), .B2(n5891), .C1(n12961), .C2(n15332), .A(
        n5638), .ZN(n5631) );
  OAI22_X1 U4009 ( .A1(n15364), .A2(n12958), .B1(n15396), .B2(n12955), .ZN(
        n5638) );
  AOI221_X1 U4010 ( .B1(n13018), .B2(n6148), .C1(n13015), .C2(n15679), .A(
        n5561), .ZN(n5558) );
  OAI22_X1 U4011 ( .A1(n14978), .A2(n13012), .B1(n15968), .B2(n13009), .ZN(
        n5561) );
  AOI221_X1 U4012 ( .B1(n12964), .B2(n5892), .C1(n12961), .C2(n15331), .A(
        n5576), .ZN(n5570) );
  OAI22_X1 U4013 ( .A1(n15363), .A2(n12958), .B1(n15395), .B2(n12955), .ZN(
        n5576) );
  AOI221_X1 U4014 ( .B1(n13018), .B2(n6149), .C1(n13015), .C2(n15678), .A(
        n5500), .ZN(n5496) );
  OAI22_X1 U4015 ( .A1(n14977), .A2(n13012), .B1(n15967), .B2(n13009), .ZN(
        n5500) );
  AOI221_X1 U4016 ( .B1(n12964), .B2(n5893), .C1(n12961), .C2(n15330), .A(
        n5514), .ZN(n5509) );
  OAI22_X1 U4017 ( .A1(n15362), .A2(n12958), .B1(n15394), .B2(n12955), .ZN(
        n5514) );
  AOI221_X1 U4018 ( .B1(n13018), .B2(n6150), .C1(n13015), .C2(n15677), .A(
        n5440), .ZN(n5436) );
  OAI22_X1 U4019 ( .A1(n14976), .A2(n13012), .B1(n15966), .B2(n13009), .ZN(
        n5440) );
  AOI221_X1 U4020 ( .B1(n12964), .B2(n5894), .C1(n12961), .C2(n15329), .A(
        n5451), .ZN(n5448) );
  OAI22_X1 U4021 ( .A1(n15361), .A2(n12958), .B1(n15393), .B2(n12955), .ZN(
        n5451) );
  AOI221_X1 U4022 ( .B1(n13018), .B2(n6151), .C1(n13015), .C2(n15676), .A(
        n5388), .ZN(n5382) );
  OAI22_X1 U4023 ( .A1(n14975), .A2(n13012), .B1(n15965), .B2(n13009), .ZN(
        n5388) );
  AOI221_X1 U4024 ( .B1(n12964), .B2(n5895), .C1(n12961), .C2(n15328), .A(
        n5399), .ZN(n5394) );
  OAI22_X1 U4025 ( .A1(n15360), .A2(n12958), .B1(n15392), .B2(n12955), .ZN(
        n5399) );
  AOI221_X1 U4026 ( .B1(n13018), .B2(n6152), .C1(n13015), .C2(n15675), .A(
        n5348), .ZN(n5345) );
  OAI22_X1 U4027 ( .A1(n14974), .A2(n13012), .B1(n15964), .B2(n13009), .ZN(
        n5348) );
  AOI221_X1 U4028 ( .B1(n12964), .B2(n5896), .C1(n12961), .C2(n15327), .A(
        n5356), .ZN(n5353) );
  OAI22_X1 U4029 ( .A1(n15359), .A2(n12958), .B1(n15391), .B2(n12955), .ZN(
        n5356) );
  AOI221_X1 U4030 ( .B1(n13018), .B2(n6153), .C1(n13015), .C2(n15674), .A(
        n5311), .ZN(n5308) );
  OAI22_X1 U4031 ( .A1(n14973), .A2(n13012), .B1(n15963), .B2(n13009), .ZN(
        n5311) );
  AOI221_X1 U4032 ( .B1(n12964), .B2(n5897), .C1(n12961), .C2(n15326), .A(
        n5319), .ZN(n5316) );
  OAI22_X1 U4033 ( .A1(n15358), .A2(n12958), .B1(n15390), .B2(n12955), .ZN(
        n5319) );
  AOI221_X1 U4034 ( .B1(n13018), .B2(n6154), .C1(n13015), .C2(n15673), .A(
        n5274), .ZN(n5271) );
  OAI22_X1 U4035 ( .A1(n14972), .A2(n13012), .B1(n15962), .B2(n13009), .ZN(
        n5274) );
  AOI221_X1 U4036 ( .B1(n12964), .B2(n5898), .C1(n12961), .C2(n15325), .A(
        n5282), .ZN(n5279) );
  OAI22_X1 U4037 ( .A1(n15357), .A2(n12958), .B1(n15389), .B2(n12955), .ZN(
        n5282) );
  AOI221_X1 U4038 ( .B1(n13018), .B2(n6155), .C1(n13015), .C2(n15672), .A(
        n5237), .ZN(n5234) );
  OAI22_X1 U4039 ( .A1(n14971), .A2(n13012), .B1(n15961), .B2(n13009), .ZN(
        n5237) );
  AOI221_X1 U4040 ( .B1(n12964), .B2(n5899), .C1(n12961), .C2(n15324), .A(
        n5245), .ZN(n5242) );
  OAI22_X1 U4041 ( .A1(n15356), .A2(n12958), .B1(n15388), .B2(n12955), .ZN(
        n5245) );
  AOI221_X1 U4042 ( .B1(n13018), .B2(n6156), .C1(n13015), .C2(n15671), .A(
        n5200), .ZN(n5197) );
  OAI22_X1 U4043 ( .A1(n14970), .A2(n13012), .B1(n15960), .B2(n13009), .ZN(
        n5200) );
  AOI221_X1 U4044 ( .B1(n12964), .B2(n5900), .C1(n12961), .C2(n15323), .A(
        n5208), .ZN(n5205) );
  OAI22_X1 U4045 ( .A1(n15355), .A2(n12958), .B1(n15387), .B2(n12955), .ZN(
        n5208) );
  AOI221_X1 U4046 ( .B1(n13018), .B2(n6157), .C1(n13015), .C2(n15670), .A(
        n5163), .ZN(n5160) );
  OAI22_X1 U4047 ( .A1(n14969), .A2(n13012), .B1(n15959), .B2(n13009), .ZN(
        n5163) );
  AOI221_X1 U4048 ( .B1(n12964), .B2(n5901), .C1(n12961), .C2(n15322), .A(
        n5171), .ZN(n5168) );
  OAI22_X1 U4049 ( .A1(n15354), .A2(n12958), .B1(n15386), .B2(n12955), .ZN(
        n5171) );
  AOI221_X1 U4050 ( .B1(n13019), .B2(n6158), .C1(n13016), .C2(n15669), .A(
        n5126), .ZN(n5123) );
  OAI22_X1 U4051 ( .A1(n14968), .A2(n13013), .B1(n15958), .B2(n13010), .ZN(
        n5126) );
  AOI221_X1 U4052 ( .B1(n12965), .B2(n5902), .C1(n12962), .C2(n15321), .A(
        n5134), .ZN(n5131) );
  OAI22_X1 U4053 ( .A1(n15353), .A2(n12959), .B1(n15385), .B2(n12956), .ZN(
        n5134) );
  AOI221_X1 U4054 ( .B1(n13019), .B2(n6159), .C1(n13016), .C2(n15668), .A(
        n5089), .ZN(n5086) );
  OAI22_X1 U4055 ( .A1(n14967), .A2(n13013), .B1(n15957), .B2(n13010), .ZN(
        n5089) );
  AOI221_X1 U4056 ( .B1(n12965), .B2(n5903), .C1(n12962), .C2(n15320), .A(
        n5097), .ZN(n5094) );
  OAI22_X1 U4057 ( .A1(n15352), .A2(n12959), .B1(n15384), .B2(n12956), .ZN(
        n5097) );
  AOI221_X1 U4058 ( .B1(n13019), .B2(n6160), .C1(n13016), .C2(n15667), .A(
        n5052), .ZN(n5049) );
  OAI22_X1 U4059 ( .A1(n14966), .A2(n13013), .B1(n15956), .B2(n13010), .ZN(
        n5052) );
  AOI221_X1 U4060 ( .B1(n12965), .B2(n5904), .C1(n12962), .C2(n15319), .A(
        n5060), .ZN(n5057) );
  OAI22_X1 U4061 ( .A1(n15351), .A2(n12959), .B1(n15383), .B2(n12956), .ZN(
        n5060) );
  AOI221_X1 U4062 ( .B1(n13019), .B2(n6161), .C1(n13016), .C2(n15666), .A(
        n5015), .ZN(n5012) );
  OAI22_X1 U4063 ( .A1(n14965), .A2(n13013), .B1(n15955), .B2(n13010), .ZN(
        n5015) );
  AOI221_X1 U4064 ( .B1(n12965), .B2(n5905), .C1(n12962), .C2(n15318), .A(
        n5023), .ZN(n5020) );
  OAI22_X1 U4065 ( .A1(n15350), .A2(n12959), .B1(n15382), .B2(n12956), .ZN(
        n5023) );
  AOI221_X1 U4066 ( .B1(n13019), .B2(n6162), .C1(n13016), .C2(n15665), .A(
        n4978), .ZN(n4975) );
  OAI22_X1 U4067 ( .A1(n14964), .A2(n13013), .B1(n15954), .B2(n13010), .ZN(
        n4978) );
  AOI221_X1 U4068 ( .B1(n12965), .B2(n5906), .C1(n12962), .C2(n15317), .A(
        n4986), .ZN(n4983) );
  OAI22_X1 U4069 ( .A1(n15349), .A2(n12959), .B1(n15381), .B2(n12956), .ZN(
        n4986) );
  AOI221_X1 U4070 ( .B1(n13019), .B2(n6163), .C1(n13016), .C2(n15664), .A(
        n4941), .ZN(n4938) );
  OAI22_X1 U4071 ( .A1(n14963), .A2(n13013), .B1(n15953), .B2(n13010), .ZN(
        n4941) );
  AOI221_X1 U4072 ( .B1(n12965), .B2(n5907), .C1(n12962), .C2(n15316), .A(
        n4949), .ZN(n4946) );
  OAI22_X1 U4073 ( .A1(n15348), .A2(n12959), .B1(n15380), .B2(n12956), .ZN(
        n4949) );
  AOI221_X1 U4074 ( .B1(n13019), .B2(n6164), .C1(n13016), .C2(n15663), .A(
        n4904), .ZN(n4901) );
  OAI22_X1 U4075 ( .A1(n14962), .A2(n13013), .B1(n15952), .B2(n13010), .ZN(
        n4904) );
  AOI221_X1 U4076 ( .B1(n12965), .B2(n5908), .C1(n12962), .C2(n15315), .A(
        n4912), .ZN(n4909) );
  OAI22_X1 U4077 ( .A1(n15347), .A2(n12959), .B1(n15379), .B2(n12956), .ZN(
        n4912) );
  AOI221_X1 U4078 ( .B1(n13019), .B2(n6165), .C1(n13016), .C2(n15662), .A(
        n4867), .ZN(n4864) );
  OAI22_X1 U4079 ( .A1(n14961), .A2(n13013), .B1(n15951), .B2(n13010), .ZN(
        n4867) );
  AOI221_X1 U4080 ( .B1(n12965), .B2(n5909), .C1(n12962), .C2(n15314), .A(
        n4875), .ZN(n4872) );
  OAI22_X1 U4081 ( .A1(n15346), .A2(n12959), .B1(n15378), .B2(n12956), .ZN(
        n4875) );
  AOI221_X1 U4082 ( .B1(n13019), .B2(n6166), .C1(n13016), .C2(n15661), .A(
        n4830), .ZN(n4827) );
  OAI22_X1 U4083 ( .A1(n14960), .A2(n13013), .B1(n15950), .B2(n13010), .ZN(
        n4830) );
  AOI221_X1 U4084 ( .B1(n12965), .B2(n5910), .C1(n12962), .C2(n15313), .A(
        n4838), .ZN(n4835) );
  OAI22_X1 U4085 ( .A1(n15345), .A2(n12959), .B1(n15377), .B2(n12956), .ZN(
        n4838) );
  AOI221_X1 U4086 ( .B1(n13019), .B2(n6167), .C1(n13016), .C2(n15660), .A(
        n4793), .ZN(n4790) );
  OAI22_X1 U4087 ( .A1(n14959), .A2(n13013), .B1(n15949), .B2(n13010), .ZN(
        n4793) );
  AOI221_X1 U4088 ( .B1(n12965), .B2(n5911), .C1(n12962), .C2(n15312), .A(
        n4801), .ZN(n4798) );
  OAI22_X1 U4089 ( .A1(n15344), .A2(n12959), .B1(n15376), .B2(n12956), .ZN(
        n4801) );
  AOI221_X1 U4090 ( .B1(n13019), .B2(n6168), .C1(n13016), .C2(n15659), .A(
        n4756), .ZN(n4753) );
  OAI22_X1 U4091 ( .A1(n14958), .A2(n13013), .B1(n15948), .B2(n13010), .ZN(
        n4756) );
  AOI221_X1 U4092 ( .B1(n12965), .B2(n5912), .C1(n12962), .C2(n15311), .A(
        n4764), .ZN(n4761) );
  OAI22_X1 U4093 ( .A1(n15343), .A2(n12959), .B1(n15375), .B2(n12956), .ZN(
        n4764) );
  AOI221_X1 U4094 ( .B1(n13019), .B2(n6169), .C1(n13016), .C2(n15658), .A(
        n4719), .ZN(n4716) );
  OAI22_X1 U4095 ( .A1(n14957), .A2(n13013), .B1(n15947), .B2(n13010), .ZN(
        n4719) );
  AOI221_X1 U4096 ( .B1(n12965), .B2(n5913), .C1(n12962), .C2(n15310), .A(
        n4727), .ZN(n4724) );
  OAI22_X1 U4097 ( .A1(n15342), .A2(n12959), .B1(n15374), .B2(n12956), .ZN(
        n4727) );
  AOI221_X1 U4098 ( .B1(n12966), .B2(n5914), .C1(n12963), .C2(n15309), .A(
        n4690), .ZN(n4687) );
  OAI22_X1 U4099 ( .A1(n15341), .A2(n12960), .B1(n15373), .B2(n12957), .ZN(
        n4690) );
  AOI221_X1 U4100 ( .B1(n13246), .B2(n6146), .C1(n13243), .C2(n15681), .A(
        n4300), .ZN(n4296) );
  OAI22_X1 U4101 ( .A1(n14980), .A2(n13240), .B1(n15970), .B2(n13237), .ZN(
        n4300) );
  AOI221_X1 U4102 ( .B1(n13192), .B2(n5890), .C1(n13189), .C2(n15333), .A(
        n4309), .ZN(n4306) );
  OAI22_X1 U4103 ( .A1(n15365), .A2(n13186), .B1(n15397), .B2(n13183), .ZN(
        n4309) );
  AOI221_X1 U4104 ( .B1(n13246), .B2(n6147), .C1(n13243), .C2(n15680), .A(
        n4249), .ZN(n4246) );
  OAI22_X1 U4105 ( .A1(n14979), .A2(n13240), .B1(n15969), .B2(n13237), .ZN(
        n4249) );
  AOI221_X1 U4106 ( .B1(n13192), .B2(n5891), .C1(n13189), .C2(n15332), .A(
        n4257), .ZN(n4254) );
  OAI22_X1 U4107 ( .A1(n15364), .A2(n13186), .B1(n15396), .B2(n13183), .ZN(
        n4257) );
  AOI221_X1 U4108 ( .B1(n13246), .B2(n6148), .C1(n13243), .C2(n15679), .A(
        n4212), .ZN(n4209) );
  OAI22_X1 U4109 ( .A1(n14978), .A2(n13240), .B1(n15968), .B2(n13237), .ZN(
        n4212) );
  AOI221_X1 U4110 ( .B1(n13192), .B2(n5892), .C1(n13189), .C2(n15331), .A(
        n4220), .ZN(n4217) );
  OAI22_X1 U4111 ( .A1(n15363), .A2(n13186), .B1(n15395), .B2(n13183), .ZN(
        n4220) );
  AOI221_X1 U4112 ( .B1(n13246), .B2(n6149), .C1(n13243), .C2(n15678), .A(
        n4175), .ZN(n4172) );
  OAI22_X1 U4113 ( .A1(n14977), .A2(n13240), .B1(n15967), .B2(n13237), .ZN(
        n4175) );
  AOI221_X1 U4114 ( .B1(n13192), .B2(n5893), .C1(n13189), .C2(n15330), .A(
        n4183), .ZN(n4180) );
  OAI22_X1 U4115 ( .A1(n15362), .A2(n13186), .B1(n15394), .B2(n13183), .ZN(
        n4183) );
  AOI221_X1 U4116 ( .B1(n13246), .B2(n6150), .C1(n13243), .C2(n15677), .A(
        n4138), .ZN(n4135) );
  OAI22_X1 U4117 ( .A1(n14976), .A2(n13240), .B1(n15966), .B2(n13237), .ZN(
        n4138) );
  AOI221_X1 U4118 ( .B1(n13192), .B2(n5894), .C1(n13189), .C2(n15329), .A(
        n4146), .ZN(n4143) );
  OAI22_X1 U4119 ( .A1(n15361), .A2(n13186), .B1(n15393), .B2(n13183), .ZN(
        n4146) );
  AOI221_X1 U4120 ( .B1(n13246), .B2(n6151), .C1(n13243), .C2(n15676), .A(
        n4101), .ZN(n4098) );
  OAI22_X1 U4121 ( .A1(n14975), .A2(n13240), .B1(n15965), .B2(n13237), .ZN(
        n4101) );
  AOI221_X1 U4122 ( .B1(n13192), .B2(n5895), .C1(n13189), .C2(n15328), .A(
        n4109), .ZN(n4106) );
  OAI22_X1 U4123 ( .A1(n15360), .A2(n13186), .B1(n15392), .B2(n13183), .ZN(
        n4109) );
  AOI221_X1 U4124 ( .B1(n13246), .B2(n6152), .C1(n13243), .C2(n15675), .A(
        n4064), .ZN(n4061) );
  OAI22_X1 U4125 ( .A1(n14974), .A2(n13240), .B1(n15964), .B2(n13237), .ZN(
        n4064) );
  AOI221_X1 U4126 ( .B1(n13192), .B2(n5896), .C1(n13189), .C2(n15327), .A(
        n4072), .ZN(n4069) );
  OAI22_X1 U4127 ( .A1(n15359), .A2(n13186), .B1(n15391), .B2(n13183), .ZN(
        n4072) );
  AOI221_X1 U4128 ( .B1(n13246), .B2(n6153), .C1(n13243), .C2(n15674), .A(
        n4027), .ZN(n4024) );
  OAI22_X1 U4129 ( .A1(n14973), .A2(n13240), .B1(n15963), .B2(n13237), .ZN(
        n4027) );
  AOI221_X1 U4130 ( .B1(n13192), .B2(n5897), .C1(n13189), .C2(n15326), .A(
        n4035), .ZN(n4032) );
  OAI22_X1 U4131 ( .A1(n15358), .A2(n13186), .B1(n15390), .B2(n13183), .ZN(
        n4035) );
  AOI221_X1 U4132 ( .B1(n13246), .B2(n6154), .C1(n13243), .C2(n15673), .A(
        n3990), .ZN(n3987) );
  OAI22_X1 U4133 ( .A1(n14972), .A2(n13240), .B1(n15962), .B2(n13237), .ZN(
        n3990) );
  AOI221_X1 U4134 ( .B1(n13192), .B2(n5898), .C1(n13189), .C2(n15325), .A(
        n3998), .ZN(n3995) );
  OAI22_X1 U4135 ( .A1(n15357), .A2(n13186), .B1(n15389), .B2(n13183), .ZN(
        n3998) );
  AOI221_X1 U4136 ( .B1(n13246), .B2(n6155), .C1(n13243), .C2(n15672), .A(
        n3953), .ZN(n3950) );
  OAI22_X1 U4137 ( .A1(n14971), .A2(n13240), .B1(n15961), .B2(n13237), .ZN(
        n3953) );
  AOI221_X1 U4138 ( .B1(n13192), .B2(n5899), .C1(n13189), .C2(n15324), .A(
        n3961), .ZN(n3958) );
  OAI22_X1 U4139 ( .A1(n15356), .A2(n13186), .B1(n15388), .B2(n13183), .ZN(
        n3961) );
  AOI221_X1 U4140 ( .B1(n13246), .B2(n6156), .C1(n13243), .C2(n15671), .A(
        n3916), .ZN(n3913) );
  OAI22_X1 U4141 ( .A1(n14970), .A2(n13240), .B1(n15960), .B2(n13237), .ZN(
        n3916) );
  AOI221_X1 U4142 ( .B1(n13192), .B2(n5900), .C1(n13189), .C2(n15323), .A(
        n3924), .ZN(n3921) );
  OAI22_X1 U4143 ( .A1(n15355), .A2(n13186), .B1(n15387), .B2(n13183), .ZN(
        n3924) );
  AOI221_X1 U4144 ( .B1(n13246), .B2(n6157), .C1(n13243), .C2(n15670), .A(
        n3879), .ZN(n3876) );
  OAI22_X1 U4145 ( .A1(n14969), .A2(n13240), .B1(n15959), .B2(n13237), .ZN(
        n3879) );
  AOI221_X1 U4146 ( .B1(n13192), .B2(n5901), .C1(n13189), .C2(n15322), .A(
        n3887), .ZN(n3884) );
  OAI22_X1 U4147 ( .A1(n15354), .A2(n13186), .B1(n15386), .B2(n13183), .ZN(
        n3887) );
  AOI221_X1 U4148 ( .B1(n13247), .B2(n6158), .C1(n13244), .C2(n15669), .A(
        n3842), .ZN(n3839) );
  OAI22_X1 U4149 ( .A1(n14968), .A2(n13241), .B1(n15958), .B2(n13238), .ZN(
        n3842) );
  AOI221_X1 U4150 ( .B1(n13193), .B2(n5902), .C1(n13190), .C2(n15321), .A(
        n3850), .ZN(n3847) );
  OAI22_X1 U4151 ( .A1(n15353), .A2(n13187), .B1(n15385), .B2(n13184), .ZN(
        n3850) );
  AOI221_X1 U4152 ( .B1(n13247), .B2(n6159), .C1(n13244), .C2(n15668), .A(
        n3805), .ZN(n3802) );
  OAI22_X1 U4153 ( .A1(n14967), .A2(n13241), .B1(n15957), .B2(n13238), .ZN(
        n3805) );
  AOI221_X1 U4154 ( .B1(n13193), .B2(n5903), .C1(n13190), .C2(n15320), .A(
        n3813), .ZN(n3810) );
  OAI22_X1 U4155 ( .A1(n15352), .A2(n13187), .B1(n15384), .B2(n13184), .ZN(
        n3813) );
  AOI221_X1 U4156 ( .B1(n13247), .B2(n6160), .C1(n13244), .C2(n15667), .A(
        n3768), .ZN(n3765) );
  OAI22_X1 U4157 ( .A1(n14966), .A2(n13241), .B1(n15956), .B2(n13238), .ZN(
        n3768) );
  AOI221_X1 U4158 ( .B1(n13193), .B2(n5904), .C1(n13190), .C2(n15319), .A(
        n3776), .ZN(n3773) );
  OAI22_X1 U4159 ( .A1(n15351), .A2(n13187), .B1(n15383), .B2(n13184), .ZN(
        n3776) );
  AOI221_X1 U4160 ( .B1(n13247), .B2(n6161), .C1(n13244), .C2(n15666), .A(
        n3731), .ZN(n3728) );
  OAI22_X1 U4161 ( .A1(n14965), .A2(n13241), .B1(n15955), .B2(n13238), .ZN(
        n3731) );
  AOI221_X1 U4162 ( .B1(n13193), .B2(n5905), .C1(n13190), .C2(n15318), .A(
        n3739), .ZN(n3736) );
  OAI22_X1 U4163 ( .A1(n15350), .A2(n13187), .B1(n15382), .B2(n13184), .ZN(
        n3739) );
  AOI221_X1 U4164 ( .B1(n13247), .B2(n6162), .C1(n13244), .C2(n15665), .A(
        n3694), .ZN(n3691) );
  OAI22_X1 U4165 ( .A1(n14964), .A2(n13241), .B1(n15954), .B2(n13238), .ZN(
        n3694) );
  AOI221_X1 U4166 ( .B1(n13193), .B2(n5906), .C1(n13190), .C2(n15317), .A(
        n3702), .ZN(n3699) );
  OAI22_X1 U4167 ( .A1(n15349), .A2(n13187), .B1(n15381), .B2(n13184), .ZN(
        n3702) );
  AOI221_X1 U4168 ( .B1(n13247), .B2(n6163), .C1(n13244), .C2(n15664), .A(
        n3657), .ZN(n3654) );
  OAI22_X1 U4169 ( .A1(n14963), .A2(n13241), .B1(n15953), .B2(n13238), .ZN(
        n3657) );
  AOI221_X1 U4170 ( .B1(n13193), .B2(n5907), .C1(n13190), .C2(n15316), .A(
        n3665), .ZN(n3662) );
  OAI22_X1 U4171 ( .A1(n15348), .A2(n13187), .B1(n15380), .B2(n13184), .ZN(
        n3665) );
  AOI221_X1 U4172 ( .B1(n13247), .B2(n6164), .C1(n13244), .C2(n15663), .A(
        n3620), .ZN(n3617) );
  OAI22_X1 U4173 ( .A1(n14962), .A2(n13241), .B1(n15952), .B2(n13238), .ZN(
        n3620) );
  AOI221_X1 U4174 ( .B1(n13193), .B2(n5908), .C1(n13190), .C2(n15315), .A(
        n3628), .ZN(n3625) );
  OAI22_X1 U4175 ( .A1(n15347), .A2(n13187), .B1(n15379), .B2(n13184), .ZN(
        n3628) );
  AOI221_X1 U4176 ( .B1(n13247), .B2(n6165), .C1(n13244), .C2(n15662), .A(
        n3583), .ZN(n3580) );
  OAI22_X1 U4177 ( .A1(n14961), .A2(n13241), .B1(n15951), .B2(n13238), .ZN(
        n3583) );
  AOI221_X1 U4178 ( .B1(n13193), .B2(n5909), .C1(n13190), .C2(n15314), .A(
        n3591), .ZN(n3588) );
  OAI22_X1 U4179 ( .A1(n15346), .A2(n13187), .B1(n15378), .B2(n13184), .ZN(
        n3591) );
  AOI221_X1 U4180 ( .B1(n13247), .B2(n6166), .C1(n13244), .C2(n15661), .A(
        n3546), .ZN(n3543) );
  OAI22_X1 U4181 ( .A1(n14960), .A2(n13241), .B1(n15950), .B2(n13238), .ZN(
        n3546) );
  AOI221_X1 U4182 ( .B1(n13193), .B2(n5910), .C1(n13190), .C2(n15313), .A(
        n3554), .ZN(n3551) );
  OAI22_X1 U4183 ( .A1(n15345), .A2(n13187), .B1(n15377), .B2(n13184), .ZN(
        n3554) );
  AOI221_X1 U4184 ( .B1(n13247), .B2(n6167), .C1(n13244), .C2(n15660), .A(
        n3509), .ZN(n3506) );
  OAI22_X1 U4185 ( .A1(n14959), .A2(n13241), .B1(n15949), .B2(n13238), .ZN(
        n3509) );
  AOI221_X1 U4186 ( .B1(n13193), .B2(n5911), .C1(n13190), .C2(n15312), .A(
        n3517), .ZN(n3514) );
  OAI22_X1 U4187 ( .A1(n15344), .A2(n13187), .B1(n15376), .B2(n13184), .ZN(
        n3517) );
  AOI221_X1 U4188 ( .B1(n13247), .B2(n6168), .C1(n13244), .C2(n15659), .A(
        n3472), .ZN(n3469) );
  OAI22_X1 U4189 ( .A1(n14958), .A2(n13241), .B1(n15948), .B2(n13238), .ZN(
        n3472) );
  AOI221_X1 U4190 ( .B1(n13193), .B2(n5912), .C1(n13190), .C2(n15311), .A(
        n3480), .ZN(n3477) );
  OAI22_X1 U4191 ( .A1(n15343), .A2(n13187), .B1(n15375), .B2(n13184), .ZN(
        n3480) );
  AOI221_X1 U4192 ( .B1(n13247), .B2(n6169), .C1(n13244), .C2(n15658), .A(
        n3435), .ZN(n3432) );
  OAI22_X1 U4193 ( .A1(n14957), .A2(n13241), .B1(n15947), .B2(n13238), .ZN(
        n3435) );
  AOI221_X1 U4194 ( .B1(n13193), .B2(n5913), .C1(n13190), .C2(n15310), .A(
        n3443), .ZN(n3440) );
  OAI22_X1 U4195 ( .A1(n15342), .A2(n13187), .B1(n15374), .B2(n13184), .ZN(
        n3443) );
  AOI221_X1 U4196 ( .B1(n13194), .B2(n5914), .C1(n13191), .C2(n15309), .A(
        n3406), .ZN(n3403) );
  OAI22_X1 U4197 ( .A1(n15341), .A2(n13188), .B1(n15373), .B2(n13185), .ZN(
        n3406) );
  AOI221_X1 U4198 ( .B1(n13248), .B2(n6171), .C1(n13245), .C2(n15618), .A(
        n3361), .ZN(n3358) );
  OAI22_X1 U4199 ( .A1(n14955), .A2(n13242), .B1(n15929), .B2(n13239), .ZN(
        n3361) );
  AOI221_X1 U4200 ( .B1(n13194), .B2(n5915), .C1(n13191), .C2(n15308), .A(
        n3369), .ZN(n3366) );
  OAI22_X1 U4201 ( .A1(n15340), .A2(n13188), .B1(n15372), .B2(n13185), .ZN(
        n3369) );
  AOI221_X1 U4202 ( .B1(n13248), .B2(n6172), .C1(n13245), .C2(n15617), .A(
        n3324), .ZN(n3321) );
  OAI22_X1 U4203 ( .A1(n14954), .A2(n13242), .B1(n15928), .B2(n13239), .ZN(
        n3324) );
  AOI221_X1 U4204 ( .B1(n13194), .B2(n5916), .C1(n13191), .C2(n15307), .A(
        n3332), .ZN(n3329) );
  OAI22_X1 U4205 ( .A1(n15339), .A2(n13188), .B1(n15371), .B2(n13185), .ZN(
        n3332) );
  AOI221_X1 U4206 ( .B1(n13248), .B2(n6173), .C1(n13245), .C2(n15616), .A(
        n3287), .ZN(n3284) );
  OAI22_X1 U4207 ( .A1(n14953), .A2(n13242), .B1(n15927), .B2(n13239), .ZN(
        n3287) );
  AOI221_X1 U4208 ( .B1(n13194), .B2(n5917), .C1(n13191), .C2(n15306), .A(
        n3295), .ZN(n3292) );
  OAI22_X1 U4209 ( .A1(n15338), .A2(n13188), .B1(n15370), .B2(n13185), .ZN(
        n3295) );
  OAI222_X1 U4210 ( .A1(n16079), .A2(n13383), .B1(n3224), .B2(n13380), .C1(
        n13372), .C2(n1452), .ZN(n7667) );
  NOR4_X1 U4211 ( .A1(n3225), .A2(n3226), .A3(n3227), .A4(n3228), .ZN(n3224)
         );
  NAND4_X1 U4212 ( .A1(n3253), .A2(n3254), .A3(n3255), .A4(n3256), .ZN(n3225)
         );
  NAND4_X1 U4213 ( .A1(n3245), .A2(n3246), .A3(n3247), .A4(n3248), .ZN(n3226)
         );
  OAI222_X1 U4214 ( .A1(n16078), .A2(n13383), .B1(n3187), .B2(n13380), .C1(
        n13372), .C2(n1451), .ZN(n7669) );
  NOR4_X1 U4215 ( .A1(n3188), .A2(n3189), .A3(n3190), .A4(n3191), .ZN(n3187)
         );
  NAND4_X1 U4216 ( .A1(n3216), .A2(n3217), .A3(n3218), .A4(n3219), .ZN(n3188)
         );
  NAND4_X1 U4217 ( .A1(n3208), .A2(n3209), .A3(n3210), .A4(n3211), .ZN(n3189)
         );
  OAI222_X1 U4218 ( .A1(n16077), .A2(n13383), .B1(n3150), .B2(n13380), .C1(
        n13372), .C2(n1450), .ZN(n7671) );
  NOR4_X1 U4219 ( .A1(n3151), .A2(n3152), .A3(n3153), .A4(n3154), .ZN(n3150)
         );
  NAND4_X1 U4220 ( .A1(n3179), .A2(n3180), .A3(n3181), .A4(n3182), .ZN(n3151)
         );
  NAND4_X1 U4221 ( .A1(n3171), .A2(n3172), .A3(n3173), .A4(n3174), .ZN(n3152)
         );
  OAI222_X1 U4222 ( .A1(n16076), .A2(n13383), .B1(n3039), .B2(n13380), .C1(
        n13373), .C2(n1449), .ZN(n7673) );
  NOR4_X1 U4223 ( .A1(n3042), .A2(n3043), .A3(n3044), .A4(n3045), .ZN(n3039)
         );
  NAND4_X1 U4224 ( .A1(n3124), .A2(n3125), .A3(n3126), .A4(n3127), .ZN(n3042)
         );
  NAND4_X1 U4225 ( .A1(n3098), .A2(n3099), .A3(n3100), .A4(n3101), .ZN(n3043)
         );
  OAI222_X1 U4226 ( .A1(n16107), .A2(n13153), .B1(n5641), .B2(n13150), .C1(
        n13146), .C2(n1512), .ZN(n7547) );
  NOR4_X1 U4227 ( .A1(n5644), .A2(n5646), .A3(n5648), .A4(n5649), .ZN(n5641)
         );
  NAND4_X1 U4228 ( .A1(n5720), .A2(n5722), .A3(n5724), .A4(n5726), .ZN(n5644)
         );
  NAND4_X1 U4229 ( .A1(n5700), .A2(n5702), .A3(n5704), .A4(n5706), .ZN(n5646)
         );
  OAI222_X1 U4230 ( .A1(n16106), .A2(n13153), .B1(n5580), .B2(n13150), .C1(
        n13146), .C2(n1511), .ZN(n7549) );
  NOR4_X1 U4231 ( .A1(n5581), .A2(n5584), .A3(n5586), .A4(n5588), .ZN(n5580)
         );
  NAND4_X1 U4232 ( .A1(n5629), .A2(n5630), .A3(n5631), .A4(n5634), .ZN(n5581)
         );
  NAND4_X1 U4233 ( .A1(n5616), .A2(n5618), .A3(n5619), .A4(n5620), .ZN(n5584)
         );
  OAI222_X1 U4234 ( .A1(n16105), .A2(n13153), .B1(n5519), .B2(n13150), .C1(
        n13146), .C2(n1510), .ZN(n7551) );
  NOR4_X1 U4235 ( .A1(n5520), .A2(n5521), .A3(n5524), .A4(n5526), .ZN(n5519)
         );
  NAND4_X1 U4236 ( .A1(n5568), .A2(n5569), .A3(n5570), .A4(n5571), .ZN(n5520)
         );
  NAND4_X1 U4237 ( .A1(n5554), .A2(n5556), .A3(n5558), .A4(n5559), .ZN(n5521)
         );
  OAI222_X1 U4238 ( .A1(n16104), .A2(n13153), .B1(n5458), .B2(n13150), .C1(
        n13146), .C2(n1509), .ZN(n7553) );
  NOR4_X1 U4239 ( .A1(n5459), .A2(n5460), .A3(n5461), .A4(n5464), .ZN(n5458)
         );
  NAND4_X1 U4240 ( .A1(n5506), .A2(n5508), .A3(n5509), .A4(n5510), .ZN(n5459)
         );
  NAND4_X1 U4241 ( .A1(n5491), .A2(n5494), .A3(n5496), .A4(n5498), .ZN(n5460)
         );
  OAI222_X1 U4242 ( .A1(n16103), .A2(n13153), .B1(n5402), .B2(n13150), .C1(
        n13146), .C2(n1508), .ZN(n7555) );
  NOR4_X1 U4243 ( .A1(n5404), .A2(n5406), .A3(n5408), .A4(n5409), .ZN(n5402)
         );
  NAND4_X1 U4244 ( .A1(n5444), .A2(n5446), .A3(n5448), .A4(n5449), .ZN(n5404)
         );
  NAND4_X1 U4245 ( .A1(n5432), .A2(n5434), .A3(n5436), .A4(n5438), .ZN(n5406)
         );
  OAI222_X1 U4246 ( .A1(n16102), .A2(n13153), .B1(n5359), .B2(n13150), .C1(
        n13146), .C2(n1507), .ZN(n7557) );
  NOR4_X1 U4247 ( .A1(n5360), .A2(n5361), .A3(n5362), .A4(n5363), .ZN(n5359)
         );
  NAND4_X1 U4248 ( .A1(n5391), .A2(n5392), .A3(n5394), .A4(n5396), .ZN(n5360)
         );
  NAND4_X1 U4249 ( .A1(n5380), .A2(n5381), .A3(n5382), .A4(n5384), .ZN(n5361)
         );
  OAI222_X1 U4250 ( .A1(n16101), .A2(n13153), .B1(n5322), .B2(n13150), .C1(
        n13146), .C2(n1506), .ZN(n7559) );
  NOR4_X1 U4251 ( .A1(n5323), .A2(n5324), .A3(n5325), .A4(n5326), .ZN(n5322)
         );
  NAND4_X1 U4252 ( .A1(n5351), .A2(n5352), .A3(n5353), .A4(n5354), .ZN(n5323)
         );
  NAND4_X1 U4253 ( .A1(n5343), .A2(n5344), .A3(n5345), .A4(n5346), .ZN(n5324)
         );
  OAI222_X1 U4254 ( .A1(n16100), .A2(n13153), .B1(n5285), .B2(n13150), .C1(
        n13146), .C2(n1505), .ZN(n7561) );
  NOR4_X1 U4255 ( .A1(n5286), .A2(n5287), .A3(n5288), .A4(n5289), .ZN(n5285)
         );
  NAND4_X1 U4256 ( .A1(n5314), .A2(n5315), .A3(n5316), .A4(n5317), .ZN(n5286)
         );
  NAND4_X1 U4257 ( .A1(n5306), .A2(n5307), .A3(n5308), .A4(n5309), .ZN(n5287)
         );
  OAI222_X1 U4258 ( .A1(n16099), .A2(n13153), .B1(n5248), .B2(n13150), .C1(
        n13145), .C2(n1504), .ZN(n7563) );
  NOR4_X1 U4259 ( .A1(n5249), .A2(n5250), .A3(n5251), .A4(n5252), .ZN(n5248)
         );
  NAND4_X1 U4260 ( .A1(n5277), .A2(n5278), .A3(n5279), .A4(n5280), .ZN(n5249)
         );
  NAND4_X1 U4261 ( .A1(n5269), .A2(n5270), .A3(n5271), .A4(n5272), .ZN(n5250)
         );
  OAI222_X1 U4262 ( .A1(n16098), .A2(n13153), .B1(n5211), .B2(n13150), .C1(
        n13145), .C2(n1503), .ZN(n7565) );
  NOR4_X1 U4263 ( .A1(n5212), .A2(n5213), .A3(n5214), .A4(n5215), .ZN(n5211)
         );
  NAND4_X1 U4264 ( .A1(n5240), .A2(n5241), .A3(n5242), .A4(n5243), .ZN(n5212)
         );
  NAND4_X1 U4265 ( .A1(n5232), .A2(n5233), .A3(n5234), .A4(n5235), .ZN(n5213)
         );
  OAI222_X1 U4266 ( .A1(n16097), .A2(n13153), .B1(n5174), .B2(n13150), .C1(
        n13145), .C2(n1502), .ZN(n7567) );
  NOR4_X1 U4267 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .ZN(n5174)
         );
  NAND4_X1 U4268 ( .A1(n5203), .A2(n5204), .A3(n5205), .A4(n5206), .ZN(n5175)
         );
  NAND4_X1 U4269 ( .A1(n5195), .A2(n5196), .A3(n5197), .A4(n5198), .ZN(n5176)
         );
  OAI222_X1 U4270 ( .A1(n16096), .A2(n13153), .B1(n5137), .B2(n13150), .C1(
        n13145), .C2(n1501), .ZN(n7569) );
  NOR4_X1 U4271 ( .A1(n5138), .A2(n5139), .A3(n5140), .A4(n5141), .ZN(n5137)
         );
  NAND4_X1 U4272 ( .A1(n5166), .A2(n5167), .A3(n5168), .A4(n5169), .ZN(n5138)
         );
  NAND4_X1 U4273 ( .A1(n5158), .A2(n5159), .A3(n5160), .A4(n5161), .ZN(n5139)
         );
  OAI222_X1 U4274 ( .A1(n16095), .A2(n13154), .B1(n5100), .B2(n13151), .C1(
        n13145), .C2(n1500), .ZN(n7571) );
  NOR4_X1 U4275 ( .A1(n5101), .A2(n5102), .A3(n5103), .A4(n5104), .ZN(n5100)
         );
  NAND4_X1 U4276 ( .A1(n5129), .A2(n5130), .A3(n5131), .A4(n5132), .ZN(n5101)
         );
  NAND4_X1 U4277 ( .A1(n5121), .A2(n5122), .A3(n5123), .A4(n5124), .ZN(n5102)
         );
  OAI222_X1 U4278 ( .A1(n16094), .A2(n13154), .B1(n5063), .B2(n13151), .C1(
        n13145), .C2(n1499), .ZN(n7573) );
  NOR4_X1 U4279 ( .A1(n5064), .A2(n5065), .A3(n5066), .A4(n5067), .ZN(n5063)
         );
  NAND4_X1 U4280 ( .A1(n5092), .A2(n5093), .A3(n5094), .A4(n5095), .ZN(n5064)
         );
  NAND4_X1 U4281 ( .A1(n5084), .A2(n5085), .A3(n5086), .A4(n5087), .ZN(n5065)
         );
  OAI222_X1 U4282 ( .A1(n16093), .A2(n13154), .B1(n5026), .B2(n13151), .C1(
        n13145), .C2(n1498), .ZN(n7575) );
  NOR4_X1 U4283 ( .A1(n5027), .A2(n5028), .A3(n5029), .A4(n5030), .ZN(n5026)
         );
  NAND4_X1 U4284 ( .A1(n5055), .A2(n5056), .A3(n5057), .A4(n5058), .ZN(n5027)
         );
  NAND4_X1 U4285 ( .A1(n5047), .A2(n5048), .A3(n5049), .A4(n5050), .ZN(n5028)
         );
  OAI222_X1 U4286 ( .A1(n16092), .A2(n13154), .B1(n4989), .B2(n13151), .C1(
        n13145), .C2(n1497), .ZN(n7577) );
  NOR4_X1 U4287 ( .A1(n4990), .A2(n4991), .A3(n4992), .A4(n4993), .ZN(n4989)
         );
  NAND4_X1 U4288 ( .A1(n5018), .A2(n5019), .A3(n5020), .A4(n5021), .ZN(n4990)
         );
  NAND4_X1 U4289 ( .A1(n5010), .A2(n5011), .A3(n5012), .A4(n5013), .ZN(n4991)
         );
  OAI222_X1 U4290 ( .A1(n16091), .A2(n13154), .B1(n4952), .B2(n13151), .C1(
        n13145), .C2(n1496), .ZN(n7579) );
  NOR4_X1 U4291 ( .A1(n4953), .A2(n4954), .A3(n4955), .A4(n4956), .ZN(n4952)
         );
  NAND4_X1 U4292 ( .A1(n4981), .A2(n4982), .A3(n4983), .A4(n4984), .ZN(n4953)
         );
  NAND4_X1 U4293 ( .A1(n4973), .A2(n4974), .A3(n4975), .A4(n4976), .ZN(n4954)
         );
  OAI222_X1 U4294 ( .A1(n16090), .A2(n13154), .B1(n4915), .B2(n13151), .C1(
        n13145), .C2(n1495), .ZN(n7581) );
  NOR4_X1 U4295 ( .A1(n4916), .A2(n4917), .A3(n4918), .A4(n4919), .ZN(n4915)
         );
  NAND4_X1 U4296 ( .A1(n4944), .A2(n4945), .A3(n4946), .A4(n4947), .ZN(n4916)
         );
  NAND4_X1 U4297 ( .A1(n4936), .A2(n4937), .A3(n4938), .A4(n4939), .ZN(n4917)
         );
  OAI222_X1 U4298 ( .A1(n16089), .A2(n13154), .B1(n4878), .B2(n13151), .C1(
        n13145), .C2(n1494), .ZN(n7583) );
  NOR4_X1 U4299 ( .A1(n4879), .A2(n4880), .A3(n4881), .A4(n4882), .ZN(n4878)
         );
  NAND4_X1 U4300 ( .A1(n4907), .A2(n4908), .A3(n4909), .A4(n4910), .ZN(n4879)
         );
  NAND4_X1 U4301 ( .A1(n4899), .A2(n4900), .A3(n4901), .A4(n4902), .ZN(n4880)
         );
  OAI222_X1 U4302 ( .A1(n16088), .A2(n13154), .B1(n4841), .B2(n13151), .C1(
        n13144), .C2(n1493), .ZN(n7585) );
  NOR4_X1 U4303 ( .A1(n4842), .A2(n4843), .A3(n4844), .A4(n4845), .ZN(n4841)
         );
  NAND4_X1 U4304 ( .A1(n4870), .A2(n4871), .A3(n4872), .A4(n4873), .ZN(n4842)
         );
  NAND4_X1 U4305 ( .A1(n4862), .A2(n4863), .A3(n4864), .A4(n4865), .ZN(n4843)
         );
  OAI222_X1 U4306 ( .A1(n16087), .A2(n13154), .B1(n4804), .B2(n13151), .C1(
        n13144), .C2(n1492), .ZN(n7587) );
  NOR4_X1 U4307 ( .A1(n4805), .A2(n4806), .A3(n4807), .A4(n4808), .ZN(n4804)
         );
  NAND4_X1 U4308 ( .A1(n4833), .A2(n4834), .A3(n4835), .A4(n4836), .ZN(n4805)
         );
  NAND4_X1 U4309 ( .A1(n4825), .A2(n4826), .A3(n4827), .A4(n4828), .ZN(n4806)
         );
  OAI222_X1 U4310 ( .A1(n16086), .A2(n13154), .B1(n4767), .B2(n13151), .C1(
        n13144), .C2(n1491), .ZN(n7589) );
  NOR4_X1 U4311 ( .A1(n4768), .A2(n4769), .A3(n4770), .A4(n4771), .ZN(n4767)
         );
  NAND4_X1 U4312 ( .A1(n4796), .A2(n4797), .A3(n4798), .A4(n4799), .ZN(n4768)
         );
  NAND4_X1 U4313 ( .A1(n4788), .A2(n4789), .A3(n4790), .A4(n4791), .ZN(n4769)
         );
  OAI222_X1 U4314 ( .A1(n16085), .A2(n13154), .B1(n4730), .B2(n13151), .C1(
        n13144), .C2(n1490), .ZN(n7591) );
  NOR4_X1 U4315 ( .A1(n4731), .A2(n4732), .A3(n4733), .A4(n4734), .ZN(n4730)
         );
  NAND4_X1 U4316 ( .A1(n4759), .A2(n4760), .A3(n4761), .A4(n4762), .ZN(n4731)
         );
  NAND4_X1 U4317 ( .A1(n4751), .A2(n4752), .A3(n4753), .A4(n4754), .ZN(n4732)
         );
  OAI222_X1 U4318 ( .A1(n16084), .A2(n13154), .B1(n4693), .B2(n13151), .C1(
        n13144), .C2(n1489), .ZN(n7593) );
  NOR4_X1 U4319 ( .A1(n4694), .A2(n4695), .A3(n4696), .A4(n4697), .ZN(n4693)
         );
  NAND4_X1 U4320 ( .A1(n4722), .A2(n4723), .A3(n4724), .A4(n4725), .ZN(n4694)
         );
  NAND4_X1 U4321 ( .A1(n4714), .A2(n4715), .A3(n4716), .A4(n4717), .ZN(n4695)
         );
  OAI222_X1 U4322 ( .A1(n16083), .A2(n13154), .B1(n4656), .B2(n13152), .C1(
        n13144), .C2(n1488), .ZN(n7595) );
  NOR4_X1 U4323 ( .A1(n4657), .A2(n4658), .A3(n4659), .A4(n4660), .ZN(n4656)
         );
  NAND4_X1 U4324 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .ZN(n4657)
         );
  NAND4_X1 U4325 ( .A1(n4677), .A2(n4678), .A3(n4679), .A4(n4680), .ZN(n4658)
         );
  OAI222_X1 U4326 ( .A1(n16107), .A2(n13381), .B1(n4260), .B2(n13378), .C1(
        n13374), .C2(n1480), .ZN(n7611) );
  NOR4_X1 U4327 ( .A1(n4261), .A2(n4262), .A3(n4263), .A4(n4264), .ZN(n4260)
         );
  NAND4_X1 U4328 ( .A1(n4304), .A2(n4305), .A3(n4306), .A4(n4307), .ZN(n4261)
         );
  NAND4_X1 U4329 ( .A1(n4294), .A2(n4295), .A3(n4296), .A4(n4297), .ZN(n4262)
         );
  OAI222_X1 U4330 ( .A1(n16106), .A2(n13381), .B1(n4223), .B2(n13378), .C1(
        n13374), .C2(n1479), .ZN(n7613) );
  NOR4_X1 U4331 ( .A1(n4224), .A2(n4225), .A3(n4226), .A4(n4227), .ZN(n4223)
         );
  NAND4_X1 U4332 ( .A1(n4252), .A2(n4253), .A3(n4254), .A4(n4255), .ZN(n4224)
         );
  NAND4_X1 U4333 ( .A1(n4244), .A2(n4245), .A3(n4246), .A4(n4247), .ZN(n4225)
         );
  OAI222_X1 U4334 ( .A1(n16105), .A2(n13381), .B1(n4186), .B2(n13378), .C1(
        n13374), .C2(n1478), .ZN(n7615) );
  NOR4_X1 U4335 ( .A1(n4187), .A2(n4188), .A3(n4189), .A4(n4190), .ZN(n4186)
         );
  NAND4_X1 U4336 ( .A1(n4215), .A2(n4216), .A3(n4217), .A4(n4218), .ZN(n4187)
         );
  NAND4_X1 U4337 ( .A1(n4207), .A2(n4208), .A3(n4209), .A4(n4210), .ZN(n4188)
         );
  OAI222_X1 U4338 ( .A1(n16104), .A2(n13381), .B1(n4149), .B2(n13378), .C1(
        n13374), .C2(n1477), .ZN(n7617) );
  NOR4_X1 U4339 ( .A1(n4150), .A2(n4151), .A3(n4152), .A4(n4153), .ZN(n4149)
         );
  NAND4_X1 U4340 ( .A1(n4178), .A2(n4179), .A3(n4180), .A4(n4181), .ZN(n4150)
         );
  NAND4_X1 U4341 ( .A1(n4170), .A2(n4171), .A3(n4172), .A4(n4173), .ZN(n4151)
         );
  OAI222_X1 U4342 ( .A1(n16103), .A2(n13381), .B1(n4112), .B2(n13378), .C1(
        n13374), .C2(n1476), .ZN(n7619) );
  NOR4_X1 U4343 ( .A1(n4113), .A2(n4114), .A3(n4115), .A4(n4116), .ZN(n4112)
         );
  NAND4_X1 U4344 ( .A1(n4141), .A2(n4142), .A3(n4143), .A4(n4144), .ZN(n4113)
         );
  NAND4_X1 U4345 ( .A1(n4133), .A2(n4134), .A3(n4135), .A4(n4136), .ZN(n4114)
         );
  OAI222_X1 U4346 ( .A1(n16102), .A2(n13381), .B1(n4075), .B2(n13378), .C1(
        n13374), .C2(n1475), .ZN(n7621) );
  NOR4_X1 U4347 ( .A1(n4076), .A2(n4077), .A3(n4078), .A4(n4079), .ZN(n4075)
         );
  NAND4_X1 U4348 ( .A1(n4104), .A2(n4105), .A3(n4106), .A4(n4107), .ZN(n4076)
         );
  NAND4_X1 U4349 ( .A1(n4096), .A2(n4097), .A3(n4098), .A4(n4099), .ZN(n4077)
         );
  OAI222_X1 U4350 ( .A1(n16101), .A2(n13381), .B1(n4038), .B2(n13378), .C1(
        n13374), .C2(n1474), .ZN(n7623) );
  NOR4_X1 U4351 ( .A1(n4039), .A2(n4040), .A3(n4041), .A4(n4042), .ZN(n4038)
         );
  NAND4_X1 U4352 ( .A1(n4067), .A2(n4068), .A3(n4069), .A4(n4070), .ZN(n4039)
         );
  NAND4_X1 U4353 ( .A1(n4059), .A2(n4060), .A3(n4061), .A4(n4062), .ZN(n4040)
         );
  OAI222_X1 U4354 ( .A1(n16100), .A2(n13381), .B1(n4001), .B2(n13378), .C1(
        n13374), .C2(n1473), .ZN(n7625) );
  NOR4_X1 U4355 ( .A1(n4002), .A2(n4003), .A3(n4004), .A4(n4005), .ZN(n4001)
         );
  NAND4_X1 U4356 ( .A1(n4030), .A2(n4031), .A3(n4032), .A4(n4033), .ZN(n4002)
         );
  NAND4_X1 U4357 ( .A1(n4022), .A2(n4023), .A3(n4024), .A4(n4025), .ZN(n4003)
         );
  OAI222_X1 U4358 ( .A1(n16099), .A2(n13381), .B1(n3964), .B2(n13378), .C1(
        n13373), .C2(n1472), .ZN(n7627) );
  NOR4_X1 U4359 ( .A1(n3965), .A2(n3966), .A3(n3967), .A4(n3968), .ZN(n3964)
         );
  NAND4_X1 U4360 ( .A1(n3993), .A2(n3994), .A3(n3995), .A4(n3996), .ZN(n3965)
         );
  NAND4_X1 U4361 ( .A1(n3985), .A2(n3986), .A3(n3987), .A4(n3988), .ZN(n3966)
         );
  OAI222_X1 U4362 ( .A1(n16098), .A2(n13381), .B1(n3927), .B2(n13378), .C1(
        n13373), .C2(n1471), .ZN(n7629) );
  NOR4_X1 U4363 ( .A1(n3928), .A2(n3929), .A3(n3930), .A4(n3931), .ZN(n3927)
         );
  NAND4_X1 U4364 ( .A1(n3956), .A2(n3957), .A3(n3958), .A4(n3959), .ZN(n3928)
         );
  NAND4_X1 U4365 ( .A1(n3948), .A2(n3949), .A3(n3950), .A4(n3951), .ZN(n3929)
         );
  OAI222_X1 U4366 ( .A1(n16097), .A2(n13381), .B1(n3890), .B2(n13378), .C1(
        n13373), .C2(n1470), .ZN(n7631) );
  NOR4_X1 U4367 ( .A1(n3891), .A2(n3892), .A3(n3893), .A4(n3894), .ZN(n3890)
         );
  NAND4_X1 U4368 ( .A1(n3919), .A2(n3920), .A3(n3921), .A4(n3922), .ZN(n3891)
         );
  NAND4_X1 U4369 ( .A1(n3911), .A2(n3912), .A3(n3913), .A4(n3914), .ZN(n3892)
         );
  OAI222_X1 U4370 ( .A1(n16096), .A2(n13381), .B1(n3853), .B2(n13378), .C1(
        n13373), .C2(n1469), .ZN(n7633) );
  NOR4_X1 U4371 ( .A1(n3854), .A2(n3855), .A3(n3856), .A4(n3857), .ZN(n3853)
         );
  NAND4_X1 U4372 ( .A1(n3882), .A2(n3883), .A3(n3884), .A4(n3885), .ZN(n3854)
         );
  NAND4_X1 U4373 ( .A1(n3874), .A2(n3875), .A3(n3876), .A4(n3877), .ZN(n3855)
         );
  OAI222_X1 U4374 ( .A1(n16095), .A2(n13382), .B1(n3816), .B2(n13379), .C1(
        n13373), .C2(n1468), .ZN(n7635) );
  NOR4_X1 U4375 ( .A1(n3817), .A2(n3818), .A3(n3819), .A4(n3820), .ZN(n3816)
         );
  NAND4_X1 U4376 ( .A1(n3845), .A2(n3846), .A3(n3847), .A4(n3848), .ZN(n3817)
         );
  NAND4_X1 U4377 ( .A1(n3837), .A2(n3838), .A3(n3839), .A4(n3840), .ZN(n3818)
         );
  OAI222_X1 U4378 ( .A1(n16094), .A2(n13382), .B1(n3779), .B2(n13379), .C1(
        n13373), .C2(n1467), .ZN(n7637) );
  NOR4_X1 U4379 ( .A1(n3780), .A2(n3781), .A3(n3782), .A4(n3783), .ZN(n3779)
         );
  NAND4_X1 U4380 ( .A1(n3808), .A2(n3809), .A3(n3810), .A4(n3811), .ZN(n3780)
         );
  NAND4_X1 U4381 ( .A1(n3800), .A2(n3801), .A3(n3802), .A4(n3803), .ZN(n3781)
         );
  OAI222_X1 U4382 ( .A1(n16093), .A2(n13382), .B1(n3742), .B2(n13379), .C1(
        n13373), .C2(n1466), .ZN(n7639) );
  NOR4_X1 U4383 ( .A1(n3743), .A2(n3744), .A3(n3745), .A4(n3746), .ZN(n3742)
         );
  NAND4_X1 U4384 ( .A1(n3771), .A2(n3772), .A3(n3773), .A4(n3774), .ZN(n3743)
         );
  NAND4_X1 U4385 ( .A1(n3763), .A2(n3764), .A3(n3765), .A4(n3766), .ZN(n3744)
         );
  OAI222_X1 U4386 ( .A1(n16092), .A2(n13382), .B1(n3705), .B2(n13379), .C1(
        n13373), .C2(n1465), .ZN(n7641) );
  NOR4_X1 U4387 ( .A1(n3706), .A2(n3707), .A3(n3708), .A4(n3709), .ZN(n3705)
         );
  NAND4_X1 U4388 ( .A1(n3734), .A2(n3735), .A3(n3736), .A4(n3737), .ZN(n3706)
         );
  NAND4_X1 U4389 ( .A1(n3726), .A2(n3727), .A3(n3728), .A4(n3729), .ZN(n3707)
         );
  OAI222_X1 U4390 ( .A1(n16091), .A2(n13382), .B1(n3668), .B2(n13379), .C1(
        n13373), .C2(n1464), .ZN(n7643) );
  NOR4_X1 U4391 ( .A1(n3669), .A2(n3670), .A3(n3671), .A4(n3672), .ZN(n3668)
         );
  NAND4_X1 U4392 ( .A1(n3697), .A2(n3698), .A3(n3699), .A4(n3700), .ZN(n3669)
         );
  NAND4_X1 U4393 ( .A1(n3689), .A2(n3690), .A3(n3691), .A4(n3692), .ZN(n3670)
         );
  OAI222_X1 U4394 ( .A1(n16090), .A2(n13382), .B1(n3631), .B2(n13379), .C1(
        n13373), .C2(n1463), .ZN(n7645) );
  NOR4_X1 U4395 ( .A1(n3632), .A2(n3633), .A3(n3634), .A4(n3635), .ZN(n3631)
         );
  NAND4_X1 U4396 ( .A1(n3660), .A2(n3661), .A3(n3662), .A4(n3663), .ZN(n3632)
         );
  NAND4_X1 U4397 ( .A1(n3652), .A2(n3653), .A3(n3654), .A4(n3655), .ZN(n3633)
         );
  OAI222_X1 U4398 ( .A1(n16089), .A2(n13382), .B1(n3594), .B2(n13379), .C1(
        n13373), .C2(n1462), .ZN(n7647) );
  NOR4_X1 U4399 ( .A1(n3595), .A2(n3596), .A3(n3597), .A4(n3598), .ZN(n3594)
         );
  NAND4_X1 U4400 ( .A1(n3623), .A2(n3624), .A3(n3625), .A4(n3626), .ZN(n3595)
         );
  NAND4_X1 U4401 ( .A1(n3615), .A2(n3616), .A3(n3617), .A4(n3618), .ZN(n3596)
         );
  OAI222_X1 U4402 ( .A1(n16088), .A2(n13382), .B1(n3557), .B2(n13379), .C1(
        n13372), .C2(n1461), .ZN(n7649) );
  NOR4_X1 U4403 ( .A1(n3558), .A2(n3559), .A3(n3560), .A4(n3561), .ZN(n3557)
         );
  NAND4_X1 U4404 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3558)
         );
  NAND4_X1 U4405 ( .A1(n3578), .A2(n3579), .A3(n3580), .A4(n3581), .ZN(n3559)
         );
  OAI222_X1 U4406 ( .A1(n16087), .A2(n13382), .B1(n3520), .B2(n13379), .C1(
        n13372), .C2(n1460), .ZN(n7651) );
  NOR4_X1 U4407 ( .A1(n3521), .A2(n3522), .A3(n3523), .A4(n3524), .ZN(n3520)
         );
  NAND4_X1 U4408 ( .A1(n3549), .A2(n3550), .A3(n3551), .A4(n3552), .ZN(n3521)
         );
  NAND4_X1 U4409 ( .A1(n3541), .A2(n3542), .A3(n3543), .A4(n3544), .ZN(n3522)
         );
  OAI222_X1 U4410 ( .A1(n16086), .A2(n13382), .B1(n3483), .B2(n13379), .C1(
        n13372), .C2(n1459), .ZN(n7653) );
  NOR4_X1 U4411 ( .A1(n3484), .A2(n3485), .A3(n3486), .A4(n3487), .ZN(n3483)
         );
  NAND4_X1 U4412 ( .A1(n3512), .A2(n3513), .A3(n3514), .A4(n3515), .ZN(n3484)
         );
  NAND4_X1 U4413 ( .A1(n3504), .A2(n3505), .A3(n3506), .A4(n3507), .ZN(n3485)
         );
  OAI222_X1 U4414 ( .A1(n16085), .A2(n13382), .B1(n3446), .B2(n13379), .C1(
        n13372), .C2(n1458), .ZN(n7655) );
  NOR4_X1 U4415 ( .A1(n3447), .A2(n3448), .A3(n3449), .A4(n3450), .ZN(n3446)
         );
  NAND4_X1 U4416 ( .A1(n3475), .A2(n3476), .A3(n3477), .A4(n3478), .ZN(n3447)
         );
  NAND4_X1 U4417 ( .A1(n3467), .A2(n3468), .A3(n3469), .A4(n3470), .ZN(n3448)
         );
  OAI222_X1 U4418 ( .A1(n16084), .A2(n13382), .B1(n3409), .B2(n13379), .C1(
        n13372), .C2(n1457), .ZN(n7657) );
  NOR4_X1 U4419 ( .A1(n3410), .A2(n3411), .A3(n3412), .A4(n3413), .ZN(n3409)
         );
  NAND4_X1 U4420 ( .A1(n3438), .A2(n3439), .A3(n3440), .A4(n3441), .ZN(n3410)
         );
  NAND4_X1 U4421 ( .A1(n3430), .A2(n3431), .A3(n3432), .A4(n3433), .ZN(n3411)
         );
  OAI222_X1 U4422 ( .A1(n16083), .A2(n13382), .B1(n3372), .B2(n13380), .C1(
        n13372), .C2(n1456), .ZN(n7659) );
  NOR4_X1 U4423 ( .A1(n3373), .A2(n3374), .A3(n3375), .A4(n3376), .ZN(n3372)
         );
  NAND4_X1 U4424 ( .A1(n3401), .A2(n3402), .A3(n3403), .A4(n3404), .ZN(n3373)
         );
  NAND4_X1 U4425 ( .A1(n3393), .A2(n3394), .A3(n3395), .A4(n3396), .ZN(n3374)
         );
  OAI222_X1 U4426 ( .A1(n16082), .A2(n13383), .B1(n3335), .B2(n13380), .C1(
        n13372), .C2(n1455), .ZN(n7661) );
  NOR4_X1 U4427 ( .A1(n3336), .A2(n3337), .A3(n3338), .A4(n3339), .ZN(n3335)
         );
  NAND4_X1 U4428 ( .A1(n3364), .A2(n3365), .A3(n3366), .A4(n3367), .ZN(n3336)
         );
  NAND4_X1 U4429 ( .A1(n3356), .A2(n3357), .A3(n3358), .A4(n3359), .ZN(n3337)
         );
  OAI222_X1 U4430 ( .A1(n16081), .A2(n13383), .B1(n3298), .B2(n13380), .C1(
        n13372), .C2(n1454), .ZN(n7663) );
  NOR4_X1 U4431 ( .A1(n3299), .A2(n3300), .A3(n3301), .A4(n3302), .ZN(n3298)
         );
  NAND4_X1 U4432 ( .A1(n3327), .A2(n3328), .A3(n3329), .A4(n3330), .ZN(n3299)
         );
  NAND4_X1 U4433 ( .A1(n3319), .A2(n3320), .A3(n3321), .A4(n3322), .ZN(n3300)
         );
  OAI222_X1 U4434 ( .A1(n16080), .A2(n13383), .B1(n3261), .B2(n13380), .C1(
        n13372), .C2(n1453), .ZN(n7665) );
  NOR4_X1 U4435 ( .A1(n3262), .A2(n3263), .A3(n3264), .A4(n3265), .ZN(n3261)
         );
  NAND4_X1 U4436 ( .A1(n3290), .A2(n3291), .A3(n3292), .A4(n3293), .ZN(n3262)
         );
  NAND4_X1 U4437 ( .A1(n3282), .A2(n3283), .A3(n3284), .A4(n3285), .ZN(n3263)
         );
  AOI221_X1 U4438 ( .B1(n13236), .B2(n6238), .C1(n13233), .C2(n15561), .A(
        n3251), .ZN(n3246) );
  OAI222_X1 U4439 ( .A1(n14919), .A2(n13230), .B1(n14855), .B2(n13227), .C1(
        n14887), .C2(n13224), .ZN(n3251) );
  AOI221_X1 U4440 ( .B1(n13236), .B2(n6239), .C1(n13233), .C2(n15560), .A(
        n3214), .ZN(n3209) );
  OAI222_X1 U4441 ( .A1(n14918), .A2(n13230), .B1(n14854), .B2(n13227), .C1(
        n14886), .C2(n13224), .ZN(n3214) );
  AOI221_X1 U4442 ( .B1(n13236), .B2(n6240), .C1(n13233), .C2(n15559), .A(
        n3177), .ZN(n3172) );
  OAI222_X1 U4443 ( .A1(n14917), .A2(n13230), .B1(n14853), .B2(n13227), .C1(
        n14885), .C2(n13224), .ZN(n3177) );
  AOI221_X1 U4444 ( .B1(n13236), .B2(n6241), .C1(n13233), .C2(n15558), .A(
        n3115), .ZN(n3099) );
  OAI222_X1 U4445 ( .A1(n14916), .A2(n13230), .B1(n14852), .B2(n13227), .C1(
        n14884), .C2(n13224), .ZN(n3115) );
  AOI221_X1 U4446 ( .B1(n13008), .B2(n6235), .C1(n13005), .C2(n15564), .A(
        n4646), .ZN(n4641) );
  OAI222_X1 U4447 ( .A1(n14922), .A2(n13002), .B1(n14858), .B2(n12999), .C1(
        n14890), .C2(n12996), .ZN(n4646) );
  AOI221_X1 U4448 ( .B1(n13008), .B2(n6236), .C1(n13005), .C2(n15563), .A(
        n4609), .ZN(n4604) );
  OAI222_X1 U4449 ( .A1(n14921), .A2(n13002), .B1(n14857), .B2(n12999), .C1(
        n14889), .C2(n12996), .ZN(n4609) );
  AOI221_X1 U4450 ( .B1(n13008), .B2(n6237), .C1(n13005), .C2(n15562), .A(
        n4572), .ZN(n4567) );
  OAI222_X1 U4451 ( .A1(n14920), .A2(n13002), .B1(n14856), .B2(n12999), .C1(
        n14888), .C2(n12996), .ZN(n4572) );
  AOI221_X1 U4452 ( .B1(n13008), .B2(n6238), .C1(n13005), .C2(n15561), .A(
        n4535), .ZN(n4530) );
  OAI222_X1 U4453 ( .A1(n14919), .A2(n13002), .B1(n14855), .B2(n12999), .C1(
        n14887), .C2(n12996), .ZN(n4535) );
  AOI221_X1 U4454 ( .B1(n13008), .B2(n6239), .C1(n13005), .C2(n15560), .A(
        n4498), .ZN(n4493) );
  OAI222_X1 U4455 ( .A1(n14918), .A2(n13002), .B1(n14854), .B2(n12999), .C1(
        n14886), .C2(n12996), .ZN(n4498) );
  AOI221_X1 U4456 ( .B1(n13008), .B2(n6240), .C1(n13005), .C2(n15559), .A(
        n4461), .ZN(n4456) );
  OAI222_X1 U4457 ( .A1(n14917), .A2(n13002), .B1(n14853), .B2(n12999), .C1(
        n14885), .C2(n12996), .ZN(n4461) );
  AOI221_X1 U4458 ( .B1(n13008), .B2(n6241), .C1(n13005), .C2(n15558), .A(
        n4399), .ZN(n4383) );
  OAI222_X1 U4459 ( .A1(n14916), .A2(n13002), .B1(n14852), .B2(n12999), .C1(
        n14884), .C2(n12996), .ZN(n4399) );
  AOI221_X1 U4460 ( .B1(n13006), .B2(n6210), .C1(n13003), .C2(n15705), .A(
        n5716), .ZN(n5702) );
  OAI222_X1 U4461 ( .A1(n14947), .A2(n13000), .B1(n14883), .B2(n12997), .C1(
        n14915), .C2(n12994), .ZN(n5716) );
  AOI221_X1 U4462 ( .B1(n12952), .B2(n5954), .C1(n12949), .C2(n15205), .A(
        n5734), .ZN(n5722) );
  OAI222_X1 U4463 ( .A1(n15301), .A2(n12946), .B1(n15237), .B2(n12943), .C1(
        n15269), .C2(n12940), .ZN(n5734) );
  AOI221_X1 U4464 ( .B1(n13006), .B2(n6211), .C1(n13003), .C2(n15704), .A(
        n5626), .ZN(n5618) );
  OAI222_X1 U4465 ( .A1(n14946), .A2(n13000), .B1(n14882), .B2(n12997), .C1(
        n14914), .C2(n12994), .ZN(n5626) );
  AOI221_X1 U4466 ( .B1(n12952), .B2(n5955), .C1(n12949), .C2(n15204), .A(
        n5639), .ZN(n5630) );
  OAI222_X1 U4467 ( .A1(n15300), .A2(n12946), .B1(n15236), .B2(n12943), .C1(
        n15268), .C2(n12940), .ZN(n5639) );
  AOI221_X1 U4468 ( .B1(n13006), .B2(n6212), .C1(n13003), .C2(n15703), .A(
        n5564), .ZN(n5556) );
  OAI222_X1 U4469 ( .A1(n14945), .A2(n13000), .B1(n14881), .B2(n12997), .C1(
        n14913), .C2(n12994), .ZN(n5564) );
  AOI221_X1 U4470 ( .B1(n12952), .B2(n5956), .C1(n12949), .C2(n15203), .A(
        n5578), .ZN(n5569) );
  OAI222_X1 U4471 ( .A1(n15299), .A2(n12946), .B1(n15235), .B2(n12943), .C1(
        n15267), .C2(n12940), .ZN(n5578) );
  AOI221_X1 U4472 ( .B1(n13006), .B2(n6213), .C1(n13003), .C2(n15702), .A(
        n5501), .ZN(n5494) );
  OAI222_X1 U4473 ( .A1(n14944), .A2(n13000), .B1(n14880), .B2(n12997), .C1(
        n14912), .C2(n12994), .ZN(n5501) );
  AOI221_X1 U4474 ( .B1(n12952), .B2(n5957), .C1(n12949), .C2(n15202), .A(
        n5516), .ZN(n5508) );
  OAI222_X1 U4475 ( .A1(n15298), .A2(n12946), .B1(n15234), .B2(n12943), .C1(
        n15266), .C2(n12940), .ZN(n5516) );
  AOI221_X1 U4476 ( .B1(n13006), .B2(n6214), .C1(n13003), .C2(n15701), .A(
        n5441), .ZN(n5434) );
  OAI222_X1 U4477 ( .A1(n14943), .A2(n13000), .B1(n14879), .B2(n12997), .C1(
        n14911), .C2(n12994), .ZN(n5441) );
  AOI221_X1 U4478 ( .B1(n12952), .B2(n5958), .C1(n12949), .C2(n15201), .A(
        n5454), .ZN(n5446) );
  OAI222_X1 U4479 ( .A1(n15297), .A2(n12946), .B1(n15233), .B2(n12943), .C1(
        n15265), .C2(n12940), .ZN(n5454) );
  AOI221_X1 U4480 ( .B1(n13006), .B2(n6215), .C1(n13003), .C2(n15700), .A(
        n5389), .ZN(n5381) );
  OAI222_X1 U4481 ( .A1(n14942), .A2(n13000), .B1(n14878), .B2(n12997), .C1(
        n14910), .C2(n12994), .ZN(n5389) );
  AOI221_X1 U4482 ( .B1(n12952), .B2(n5959), .C1(n12949), .C2(n15200), .A(
        n5400), .ZN(n5392) );
  OAI222_X1 U4483 ( .A1(n15296), .A2(n12946), .B1(n15232), .B2(n12943), .C1(
        n15264), .C2(n12940), .ZN(n5400) );
  AOI221_X1 U4484 ( .B1(n13006), .B2(n6216), .C1(n13003), .C2(n15699), .A(
        n5349), .ZN(n5344) );
  OAI222_X1 U4485 ( .A1(n14941), .A2(n13000), .B1(n14877), .B2(n12997), .C1(
        n14909), .C2(n12994), .ZN(n5349) );
  AOI221_X1 U4486 ( .B1(n12952), .B2(n5960), .C1(n12949), .C2(n15199), .A(
        n5357), .ZN(n5352) );
  OAI222_X1 U4487 ( .A1(n15295), .A2(n12946), .B1(n15231), .B2(n12943), .C1(
        n15263), .C2(n12940), .ZN(n5357) );
  AOI221_X1 U4488 ( .B1(n13006), .B2(n6217), .C1(n13003), .C2(n15698), .A(
        n5312), .ZN(n5307) );
  OAI222_X1 U4489 ( .A1(n14940), .A2(n13000), .B1(n14876), .B2(n12997), .C1(
        n14908), .C2(n12994), .ZN(n5312) );
  AOI221_X1 U4490 ( .B1(n12952), .B2(n5961), .C1(n12949), .C2(n15198), .A(
        n5320), .ZN(n5315) );
  OAI222_X1 U4491 ( .A1(n15294), .A2(n12946), .B1(n15230), .B2(n12943), .C1(
        n15262), .C2(n12940), .ZN(n5320) );
  AOI221_X1 U4492 ( .B1(n13006), .B2(n6218), .C1(n13003), .C2(n15697), .A(
        n5275), .ZN(n5270) );
  OAI222_X1 U4493 ( .A1(n14939), .A2(n13000), .B1(n14875), .B2(n12997), .C1(
        n14907), .C2(n12994), .ZN(n5275) );
  AOI221_X1 U4494 ( .B1(n12952), .B2(n5962), .C1(n12949), .C2(n15197), .A(
        n5283), .ZN(n5278) );
  OAI222_X1 U4495 ( .A1(n15293), .A2(n12946), .B1(n15229), .B2(n12943), .C1(
        n15261), .C2(n12940), .ZN(n5283) );
  AOI221_X1 U4496 ( .B1(n13006), .B2(n6219), .C1(n13003), .C2(n15696), .A(
        n5238), .ZN(n5233) );
  OAI222_X1 U4497 ( .A1(n14938), .A2(n13000), .B1(n14874), .B2(n12997), .C1(
        n14906), .C2(n12994), .ZN(n5238) );
  AOI221_X1 U4498 ( .B1(n12952), .B2(n5963), .C1(n12949), .C2(n15196), .A(
        n5246), .ZN(n5241) );
  OAI222_X1 U4499 ( .A1(n15292), .A2(n12946), .B1(n15228), .B2(n12943), .C1(
        n15260), .C2(n12940), .ZN(n5246) );
  AOI221_X1 U4500 ( .B1(n13006), .B2(n6220), .C1(n13003), .C2(n15695), .A(
        n5201), .ZN(n5196) );
  OAI222_X1 U4501 ( .A1(n14937), .A2(n13000), .B1(n14873), .B2(n12997), .C1(
        n14905), .C2(n12994), .ZN(n5201) );
  AOI221_X1 U4502 ( .B1(n12952), .B2(n5964), .C1(n12949), .C2(n15195), .A(
        n5209), .ZN(n5204) );
  OAI222_X1 U4503 ( .A1(n15291), .A2(n12946), .B1(n15227), .B2(n12943), .C1(
        n15259), .C2(n12940), .ZN(n5209) );
  AOI221_X1 U4504 ( .B1(n13006), .B2(n6221), .C1(n13003), .C2(n15694), .A(
        n5164), .ZN(n5159) );
  OAI222_X1 U4505 ( .A1(n14936), .A2(n13000), .B1(n14872), .B2(n12997), .C1(
        n14904), .C2(n12994), .ZN(n5164) );
  AOI221_X1 U4506 ( .B1(n12952), .B2(n5965), .C1(n12949), .C2(n15194), .A(
        n5172), .ZN(n5167) );
  OAI222_X1 U4507 ( .A1(n15290), .A2(n12946), .B1(n15226), .B2(n12943), .C1(
        n15258), .C2(n12940), .ZN(n5172) );
  AOI221_X1 U4508 ( .B1(n13007), .B2(n6222), .C1(n13004), .C2(n15693), .A(
        n5127), .ZN(n5122) );
  OAI222_X1 U4509 ( .A1(n14935), .A2(n13001), .B1(n14871), .B2(n12998), .C1(
        n14903), .C2(n12995), .ZN(n5127) );
  AOI221_X1 U4510 ( .B1(n12953), .B2(n5966), .C1(n12950), .C2(n15193), .A(
        n5135), .ZN(n5130) );
  OAI222_X1 U4511 ( .A1(n15289), .A2(n12947), .B1(n15225), .B2(n12944), .C1(
        n15257), .C2(n12941), .ZN(n5135) );
  AOI221_X1 U4512 ( .B1(n13007), .B2(n6223), .C1(n13004), .C2(n15692), .A(
        n5090), .ZN(n5085) );
  OAI222_X1 U4513 ( .A1(n14934), .A2(n13001), .B1(n14870), .B2(n12998), .C1(
        n14902), .C2(n12995), .ZN(n5090) );
  AOI221_X1 U4514 ( .B1(n12953), .B2(n5967), .C1(n12950), .C2(n15192), .A(
        n5098), .ZN(n5093) );
  OAI222_X1 U4515 ( .A1(n15288), .A2(n12947), .B1(n15224), .B2(n12944), .C1(
        n15256), .C2(n12941), .ZN(n5098) );
  AOI221_X1 U4516 ( .B1(n13007), .B2(n6224), .C1(n13004), .C2(n15691), .A(
        n5053), .ZN(n5048) );
  OAI222_X1 U4517 ( .A1(n14933), .A2(n13001), .B1(n14869), .B2(n12998), .C1(
        n14901), .C2(n12995), .ZN(n5053) );
  AOI221_X1 U4518 ( .B1(n12953), .B2(n5968), .C1(n12950), .C2(n15191), .A(
        n5061), .ZN(n5056) );
  OAI222_X1 U4519 ( .A1(n15287), .A2(n12947), .B1(n15223), .B2(n12944), .C1(
        n15255), .C2(n12941), .ZN(n5061) );
  AOI221_X1 U4520 ( .B1(n13007), .B2(n6225), .C1(n13004), .C2(n15690), .A(
        n5016), .ZN(n5011) );
  OAI222_X1 U4521 ( .A1(n14932), .A2(n13001), .B1(n14868), .B2(n12998), .C1(
        n14900), .C2(n12995), .ZN(n5016) );
  AOI221_X1 U4522 ( .B1(n12953), .B2(n5969), .C1(n12950), .C2(n15190), .A(
        n5024), .ZN(n5019) );
  OAI222_X1 U4523 ( .A1(n15286), .A2(n12947), .B1(n15222), .B2(n12944), .C1(
        n15254), .C2(n12941), .ZN(n5024) );
  AOI221_X1 U4524 ( .B1(n13007), .B2(n6226), .C1(n13004), .C2(n15689), .A(
        n4979), .ZN(n4974) );
  OAI222_X1 U4525 ( .A1(n14931), .A2(n13001), .B1(n14867), .B2(n12998), .C1(
        n14899), .C2(n12995), .ZN(n4979) );
  AOI221_X1 U4526 ( .B1(n12953), .B2(n5970), .C1(n12950), .C2(n15189), .A(
        n4987), .ZN(n4982) );
  OAI222_X1 U4527 ( .A1(n15285), .A2(n12947), .B1(n15221), .B2(n12944), .C1(
        n15253), .C2(n12941), .ZN(n4987) );
  AOI221_X1 U4528 ( .B1(n13007), .B2(n6227), .C1(n13004), .C2(n15688), .A(
        n4942), .ZN(n4937) );
  OAI222_X1 U4529 ( .A1(n14930), .A2(n13001), .B1(n14866), .B2(n12998), .C1(
        n14898), .C2(n12995), .ZN(n4942) );
  AOI221_X1 U4530 ( .B1(n12953), .B2(n5971), .C1(n12950), .C2(n15188), .A(
        n4950), .ZN(n4945) );
  OAI222_X1 U4531 ( .A1(n15284), .A2(n12947), .B1(n15220), .B2(n12944), .C1(
        n15252), .C2(n12941), .ZN(n4950) );
  AOI221_X1 U4532 ( .B1(n13007), .B2(n6228), .C1(n13004), .C2(n15687), .A(
        n4905), .ZN(n4900) );
  OAI222_X1 U4533 ( .A1(n14929), .A2(n13001), .B1(n14865), .B2(n12998), .C1(
        n14897), .C2(n12995), .ZN(n4905) );
  AOI221_X1 U4534 ( .B1(n12953), .B2(n5972), .C1(n12950), .C2(n15187), .A(
        n4913), .ZN(n4908) );
  OAI222_X1 U4535 ( .A1(n15283), .A2(n12947), .B1(n15219), .B2(n12944), .C1(
        n15251), .C2(n12941), .ZN(n4913) );
  AOI221_X1 U4536 ( .B1(n13007), .B2(n6229), .C1(n13004), .C2(n15686), .A(
        n4868), .ZN(n4863) );
  OAI222_X1 U4537 ( .A1(n14928), .A2(n13001), .B1(n14864), .B2(n12998), .C1(
        n14896), .C2(n12995), .ZN(n4868) );
  AOI221_X1 U4538 ( .B1(n12953), .B2(n5973), .C1(n12950), .C2(n15186), .A(
        n4876), .ZN(n4871) );
  OAI222_X1 U4539 ( .A1(n15282), .A2(n12947), .B1(n15218), .B2(n12944), .C1(
        n15250), .C2(n12941), .ZN(n4876) );
  AOI221_X1 U4540 ( .B1(n13007), .B2(n6230), .C1(n13004), .C2(n15685), .A(
        n4831), .ZN(n4826) );
  OAI222_X1 U4541 ( .A1(n14927), .A2(n13001), .B1(n14863), .B2(n12998), .C1(
        n14895), .C2(n12995), .ZN(n4831) );
  AOI221_X1 U4542 ( .B1(n12953), .B2(n5974), .C1(n12950), .C2(n15185), .A(
        n4839), .ZN(n4834) );
  OAI222_X1 U4543 ( .A1(n15281), .A2(n12947), .B1(n15217), .B2(n12944), .C1(
        n15249), .C2(n12941), .ZN(n4839) );
  AOI221_X1 U4544 ( .B1(n13007), .B2(n6231), .C1(n13004), .C2(n15684), .A(
        n4794), .ZN(n4789) );
  OAI222_X1 U4545 ( .A1(n14926), .A2(n13001), .B1(n14862), .B2(n12998), .C1(
        n14894), .C2(n12995), .ZN(n4794) );
  AOI221_X1 U4546 ( .B1(n12953), .B2(n5975), .C1(n12950), .C2(n15184), .A(
        n4802), .ZN(n4797) );
  OAI222_X1 U4547 ( .A1(n15280), .A2(n12947), .B1(n15216), .B2(n12944), .C1(
        n15248), .C2(n12941), .ZN(n4802) );
  AOI221_X1 U4548 ( .B1(n13007), .B2(n6232), .C1(n13004), .C2(n15683), .A(
        n4757), .ZN(n4752) );
  OAI222_X1 U4549 ( .A1(n14925), .A2(n13001), .B1(n14861), .B2(n12998), .C1(
        n14893), .C2(n12995), .ZN(n4757) );
  AOI221_X1 U4550 ( .B1(n12953), .B2(n5976), .C1(n12950), .C2(n15183), .A(
        n4765), .ZN(n4760) );
  OAI222_X1 U4551 ( .A1(n15279), .A2(n12947), .B1(n15215), .B2(n12944), .C1(
        n15247), .C2(n12941), .ZN(n4765) );
  AOI221_X1 U4552 ( .B1(n13007), .B2(n6233), .C1(n13004), .C2(n15682), .A(
        n4720), .ZN(n4715) );
  OAI222_X1 U4553 ( .A1(n14924), .A2(n13001), .B1(n14860), .B2(n12998), .C1(
        n14892), .C2(n12995), .ZN(n4720) );
  AOI221_X1 U4554 ( .B1(n12953), .B2(n5977), .C1(n12950), .C2(n15182), .A(
        n4728), .ZN(n4723) );
  OAI222_X1 U4555 ( .A1(n15278), .A2(n12947), .B1(n15214), .B2(n12944), .C1(
        n15246), .C2(n12941), .ZN(n4728) );
  AOI221_X1 U4556 ( .B1(n12954), .B2(n5978), .C1(n12951), .C2(n15181), .A(
        n4691), .ZN(n4686) );
  OAI222_X1 U4557 ( .A1(n15277), .A2(n12948), .B1(n15213), .B2(n12945), .C1(
        n15245), .C2(n12942), .ZN(n4691) );
  AOI221_X1 U4558 ( .B1(n13234), .B2(n6210), .C1(n13231), .C2(n15705), .A(
        n4302), .ZN(n4295) );
  OAI222_X1 U4559 ( .A1(n14947), .A2(n13228), .B1(n14883), .B2(n13225), .C1(
        n14915), .C2(n13222), .ZN(n4302) );
  AOI221_X1 U4560 ( .B1(n13180), .B2(n5954), .C1(n13177), .C2(n15205), .A(
        n4311), .ZN(n4305) );
  OAI222_X1 U4561 ( .A1(n15301), .A2(n13174), .B1(n15237), .B2(n13171), .C1(
        n15269), .C2(n13168), .ZN(n4311) );
  AOI221_X1 U4562 ( .B1(n13234), .B2(n6211), .C1(n13231), .C2(n15704), .A(
        n4250), .ZN(n4245) );
  OAI222_X1 U4563 ( .A1(n14946), .A2(n13228), .B1(n14882), .B2(n13225), .C1(
        n14914), .C2(n13222), .ZN(n4250) );
  AOI221_X1 U4564 ( .B1(n13180), .B2(n5955), .C1(n13177), .C2(n15204), .A(
        n4258), .ZN(n4253) );
  OAI222_X1 U4565 ( .A1(n15300), .A2(n13174), .B1(n15236), .B2(n13171), .C1(
        n15268), .C2(n13168), .ZN(n4258) );
  AOI221_X1 U4566 ( .B1(n13234), .B2(n6212), .C1(n13231), .C2(n15703), .A(
        n4213), .ZN(n4208) );
  OAI222_X1 U4567 ( .A1(n14945), .A2(n13228), .B1(n14881), .B2(n13225), .C1(
        n14913), .C2(n13222), .ZN(n4213) );
  AOI221_X1 U4568 ( .B1(n13180), .B2(n5956), .C1(n13177), .C2(n15203), .A(
        n4221), .ZN(n4216) );
  OAI222_X1 U4569 ( .A1(n15299), .A2(n13174), .B1(n15235), .B2(n13171), .C1(
        n15267), .C2(n13168), .ZN(n4221) );
  AOI221_X1 U4570 ( .B1(n13234), .B2(n6213), .C1(n13231), .C2(n15702), .A(
        n4176), .ZN(n4171) );
  OAI222_X1 U4571 ( .A1(n14944), .A2(n13228), .B1(n14880), .B2(n13225), .C1(
        n14912), .C2(n13222), .ZN(n4176) );
  AOI221_X1 U4572 ( .B1(n13180), .B2(n5957), .C1(n13177), .C2(n15202), .A(
        n4184), .ZN(n4179) );
  OAI222_X1 U4573 ( .A1(n15298), .A2(n13174), .B1(n15234), .B2(n13171), .C1(
        n15266), .C2(n13168), .ZN(n4184) );
  AOI221_X1 U4574 ( .B1(n13234), .B2(n6214), .C1(n13231), .C2(n15701), .A(
        n4139), .ZN(n4134) );
  OAI222_X1 U4575 ( .A1(n14943), .A2(n13228), .B1(n14879), .B2(n13225), .C1(
        n14911), .C2(n13222), .ZN(n4139) );
  AOI221_X1 U4576 ( .B1(n13180), .B2(n5958), .C1(n13177), .C2(n15201), .A(
        n4147), .ZN(n4142) );
  OAI222_X1 U4577 ( .A1(n15297), .A2(n13174), .B1(n15233), .B2(n13171), .C1(
        n15265), .C2(n13168), .ZN(n4147) );
  AOI221_X1 U4578 ( .B1(n13234), .B2(n6215), .C1(n13231), .C2(n15700), .A(
        n4102), .ZN(n4097) );
  OAI222_X1 U4579 ( .A1(n14942), .A2(n13228), .B1(n14878), .B2(n13225), .C1(
        n14910), .C2(n13222), .ZN(n4102) );
  AOI221_X1 U4580 ( .B1(n13180), .B2(n5959), .C1(n13177), .C2(n15200), .A(
        n4110), .ZN(n4105) );
  OAI222_X1 U4581 ( .A1(n15296), .A2(n13174), .B1(n15232), .B2(n13171), .C1(
        n15264), .C2(n13168), .ZN(n4110) );
  AOI221_X1 U4582 ( .B1(n13234), .B2(n6216), .C1(n13231), .C2(n15699), .A(
        n4065), .ZN(n4060) );
  OAI222_X1 U4583 ( .A1(n14941), .A2(n13228), .B1(n14877), .B2(n13225), .C1(
        n14909), .C2(n13222), .ZN(n4065) );
  AOI221_X1 U4584 ( .B1(n13180), .B2(n5960), .C1(n13177), .C2(n15199), .A(
        n4073), .ZN(n4068) );
  OAI222_X1 U4585 ( .A1(n15295), .A2(n13174), .B1(n15231), .B2(n13171), .C1(
        n15263), .C2(n13168), .ZN(n4073) );
  AOI221_X1 U4586 ( .B1(n13234), .B2(n6217), .C1(n13231), .C2(n15698), .A(
        n4028), .ZN(n4023) );
  OAI222_X1 U4587 ( .A1(n14940), .A2(n13228), .B1(n14876), .B2(n13225), .C1(
        n14908), .C2(n13222), .ZN(n4028) );
  AOI221_X1 U4588 ( .B1(n13180), .B2(n5961), .C1(n13177), .C2(n15198), .A(
        n4036), .ZN(n4031) );
  OAI222_X1 U4589 ( .A1(n15294), .A2(n13174), .B1(n15230), .B2(n13171), .C1(
        n15262), .C2(n13168), .ZN(n4036) );
  AOI221_X1 U4590 ( .B1(n13234), .B2(n6218), .C1(n13231), .C2(n15697), .A(
        n3991), .ZN(n3986) );
  OAI222_X1 U4591 ( .A1(n14939), .A2(n13228), .B1(n14875), .B2(n13225), .C1(
        n14907), .C2(n13222), .ZN(n3991) );
  AOI221_X1 U4592 ( .B1(n13180), .B2(n5962), .C1(n13177), .C2(n15197), .A(
        n3999), .ZN(n3994) );
  OAI222_X1 U4593 ( .A1(n15293), .A2(n13174), .B1(n15229), .B2(n13171), .C1(
        n15261), .C2(n13168), .ZN(n3999) );
  AOI221_X1 U4594 ( .B1(n13234), .B2(n6219), .C1(n13231), .C2(n15696), .A(
        n3954), .ZN(n3949) );
  OAI222_X1 U4595 ( .A1(n14938), .A2(n13228), .B1(n14874), .B2(n13225), .C1(
        n14906), .C2(n13222), .ZN(n3954) );
  AOI221_X1 U4596 ( .B1(n13180), .B2(n5963), .C1(n13177), .C2(n15196), .A(
        n3962), .ZN(n3957) );
  OAI222_X1 U4597 ( .A1(n15292), .A2(n13174), .B1(n15228), .B2(n13171), .C1(
        n15260), .C2(n13168), .ZN(n3962) );
  AOI221_X1 U4598 ( .B1(n13234), .B2(n6220), .C1(n13231), .C2(n15695), .A(
        n3917), .ZN(n3912) );
  OAI222_X1 U4599 ( .A1(n14937), .A2(n13228), .B1(n14873), .B2(n13225), .C1(
        n14905), .C2(n13222), .ZN(n3917) );
  AOI221_X1 U4600 ( .B1(n13180), .B2(n5964), .C1(n13177), .C2(n15195), .A(
        n3925), .ZN(n3920) );
  OAI222_X1 U4601 ( .A1(n15291), .A2(n13174), .B1(n15227), .B2(n13171), .C1(
        n15259), .C2(n13168), .ZN(n3925) );
  AOI221_X1 U4602 ( .B1(n13234), .B2(n6221), .C1(n13231), .C2(n15694), .A(
        n3880), .ZN(n3875) );
  OAI222_X1 U4603 ( .A1(n14936), .A2(n13228), .B1(n14872), .B2(n13225), .C1(
        n14904), .C2(n13222), .ZN(n3880) );
  AOI221_X1 U4604 ( .B1(n13180), .B2(n5965), .C1(n13177), .C2(n15194), .A(
        n3888), .ZN(n3883) );
  OAI222_X1 U4605 ( .A1(n15290), .A2(n13174), .B1(n15226), .B2(n13171), .C1(
        n15258), .C2(n13168), .ZN(n3888) );
  AOI221_X1 U4606 ( .B1(n13235), .B2(n6222), .C1(n13232), .C2(n15693), .A(
        n3843), .ZN(n3838) );
  OAI222_X1 U4607 ( .A1(n14935), .A2(n13229), .B1(n14871), .B2(n13226), .C1(
        n14903), .C2(n13223), .ZN(n3843) );
  AOI221_X1 U4608 ( .B1(n13181), .B2(n5966), .C1(n13178), .C2(n15193), .A(
        n3851), .ZN(n3846) );
  OAI222_X1 U4609 ( .A1(n15289), .A2(n13175), .B1(n15225), .B2(n13172), .C1(
        n15257), .C2(n13169), .ZN(n3851) );
  AOI221_X1 U4610 ( .B1(n13235), .B2(n6223), .C1(n13232), .C2(n15692), .A(
        n3806), .ZN(n3801) );
  OAI222_X1 U4611 ( .A1(n14934), .A2(n13229), .B1(n14870), .B2(n13226), .C1(
        n14902), .C2(n13223), .ZN(n3806) );
  AOI221_X1 U4612 ( .B1(n13181), .B2(n5967), .C1(n13178), .C2(n15192), .A(
        n3814), .ZN(n3809) );
  OAI222_X1 U4613 ( .A1(n15288), .A2(n13175), .B1(n15224), .B2(n13172), .C1(
        n15256), .C2(n13169), .ZN(n3814) );
  AOI221_X1 U4614 ( .B1(n13235), .B2(n6224), .C1(n13232), .C2(n15691), .A(
        n3769), .ZN(n3764) );
  OAI222_X1 U4615 ( .A1(n14933), .A2(n13229), .B1(n14869), .B2(n13226), .C1(
        n14901), .C2(n13223), .ZN(n3769) );
  AOI221_X1 U4616 ( .B1(n13181), .B2(n5968), .C1(n13178), .C2(n15191), .A(
        n3777), .ZN(n3772) );
  OAI222_X1 U4617 ( .A1(n15287), .A2(n13175), .B1(n15223), .B2(n13172), .C1(
        n15255), .C2(n13169), .ZN(n3777) );
  AOI221_X1 U4618 ( .B1(n13235), .B2(n6225), .C1(n13232), .C2(n15690), .A(
        n3732), .ZN(n3727) );
  OAI222_X1 U4619 ( .A1(n14932), .A2(n13229), .B1(n14868), .B2(n13226), .C1(
        n14900), .C2(n13223), .ZN(n3732) );
  AOI221_X1 U4620 ( .B1(n13181), .B2(n5969), .C1(n13178), .C2(n15190), .A(
        n3740), .ZN(n3735) );
  OAI222_X1 U4621 ( .A1(n15286), .A2(n13175), .B1(n15222), .B2(n13172), .C1(
        n15254), .C2(n13169), .ZN(n3740) );
  AOI221_X1 U4622 ( .B1(n13235), .B2(n6226), .C1(n13232), .C2(n15689), .A(
        n3695), .ZN(n3690) );
  OAI222_X1 U4623 ( .A1(n14931), .A2(n13229), .B1(n14867), .B2(n13226), .C1(
        n14899), .C2(n13223), .ZN(n3695) );
  AOI221_X1 U4624 ( .B1(n13181), .B2(n5970), .C1(n13178), .C2(n15189), .A(
        n3703), .ZN(n3698) );
  OAI222_X1 U4625 ( .A1(n15285), .A2(n13175), .B1(n15221), .B2(n13172), .C1(
        n15253), .C2(n13169), .ZN(n3703) );
  AOI221_X1 U4626 ( .B1(n13235), .B2(n6227), .C1(n13232), .C2(n15688), .A(
        n3658), .ZN(n3653) );
  OAI222_X1 U4627 ( .A1(n14930), .A2(n13229), .B1(n14866), .B2(n13226), .C1(
        n14898), .C2(n13223), .ZN(n3658) );
  AOI221_X1 U4628 ( .B1(n13181), .B2(n5971), .C1(n13178), .C2(n15188), .A(
        n3666), .ZN(n3661) );
  OAI222_X1 U4629 ( .A1(n15284), .A2(n13175), .B1(n15220), .B2(n13172), .C1(
        n15252), .C2(n13169), .ZN(n3666) );
  AOI221_X1 U4630 ( .B1(n13235), .B2(n6228), .C1(n13232), .C2(n15687), .A(
        n3621), .ZN(n3616) );
  OAI222_X1 U4631 ( .A1(n14929), .A2(n13229), .B1(n14865), .B2(n13226), .C1(
        n14897), .C2(n13223), .ZN(n3621) );
  AOI221_X1 U4632 ( .B1(n13181), .B2(n5972), .C1(n13178), .C2(n15187), .A(
        n3629), .ZN(n3624) );
  OAI222_X1 U4633 ( .A1(n15283), .A2(n13175), .B1(n15219), .B2(n13172), .C1(
        n15251), .C2(n13169), .ZN(n3629) );
  AOI221_X1 U4634 ( .B1(n13235), .B2(n6229), .C1(n13232), .C2(n15686), .A(
        n3584), .ZN(n3579) );
  OAI222_X1 U4635 ( .A1(n14928), .A2(n13229), .B1(n14864), .B2(n13226), .C1(
        n14896), .C2(n13223), .ZN(n3584) );
  AOI221_X1 U4636 ( .B1(n13181), .B2(n5973), .C1(n13178), .C2(n15186), .A(
        n3592), .ZN(n3587) );
  OAI222_X1 U4637 ( .A1(n15282), .A2(n13175), .B1(n15218), .B2(n13172), .C1(
        n15250), .C2(n13169), .ZN(n3592) );
  AOI221_X1 U4638 ( .B1(n13235), .B2(n6230), .C1(n13232), .C2(n15685), .A(
        n3547), .ZN(n3542) );
  OAI222_X1 U4639 ( .A1(n14927), .A2(n13229), .B1(n14863), .B2(n13226), .C1(
        n14895), .C2(n13223), .ZN(n3547) );
  AOI221_X1 U4640 ( .B1(n13181), .B2(n5974), .C1(n13178), .C2(n15185), .A(
        n3555), .ZN(n3550) );
  OAI222_X1 U4641 ( .A1(n15281), .A2(n13175), .B1(n15217), .B2(n13172), .C1(
        n15249), .C2(n13169), .ZN(n3555) );
  AOI221_X1 U4642 ( .B1(n13235), .B2(n6231), .C1(n13232), .C2(n15684), .A(
        n3510), .ZN(n3505) );
  OAI222_X1 U4643 ( .A1(n14926), .A2(n13229), .B1(n14862), .B2(n13226), .C1(
        n14894), .C2(n13223), .ZN(n3510) );
  AOI221_X1 U4644 ( .B1(n13181), .B2(n5975), .C1(n13178), .C2(n15184), .A(
        n3518), .ZN(n3513) );
  OAI222_X1 U4645 ( .A1(n15280), .A2(n13175), .B1(n15216), .B2(n13172), .C1(
        n15248), .C2(n13169), .ZN(n3518) );
  AOI221_X1 U4646 ( .B1(n13235), .B2(n6232), .C1(n13232), .C2(n15683), .A(
        n3473), .ZN(n3468) );
  OAI222_X1 U4647 ( .A1(n14925), .A2(n13229), .B1(n14861), .B2(n13226), .C1(
        n14893), .C2(n13223), .ZN(n3473) );
  AOI221_X1 U4648 ( .B1(n13181), .B2(n5976), .C1(n13178), .C2(n15183), .A(
        n3481), .ZN(n3476) );
  OAI222_X1 U4649 ( .A1(n15279), .A2(n13175), .B1(n15215), .B2(n13172), .C1(
        n15247), .C2(n13169), .ZN(n3481) );
  AOI221_X1 U4650 ( .B1(n13235), .B2(n6233), .C1(n13232), .C2(n15682), .A(
        n3436), .ZN(n3431) );
  OAI222_X1 U4651 ( .A1(n14924), .A2(n13229), .B1(n14860), .B2(n13226), .C1(
        n14892), .C2(n13223), .ZN(n3436) );
  AOI221_X1 U4652 ( .B1(n13181), .B2(n5977), .C1(n13178), .C2(n15182), .A(
        n3444), .ZN(n3439) );
  OAI222_X1 U4653 ( .A1(n15278), .A2(n13175), .B1(n15214), .B2(n13172), .C1(
        n15246), .C2(n13169), .ZN(n3444) );
  AOI221_X1 U4654 ( .B1(n13182), .B2(n5978), .C1(n13179), .C2(n15181), .A(
        n3407), .ZN(n3402) );
  OAI222_X1 U4655 ( .A1(n15277), .A2(n13176), .B1(n15213), .B2(n13173), .C1(
        n15245), .C2(n13170), .ZN(n3407) );
  AOI221_X1 U4656 ( .B1(n13236), .B2(n6235), .C1(n13233), .C2(n15564), .A(
        n3362), .ZN(n3357) );
  OAI222_X1 U4657 ( .A1(n14922), .A2(n13230), .B1(n14858), .B2(n13227), .C1(
        n14890), .C2(n13224), .ZN(n3362) );
  AOI221_X1 U4658 ( .B1(n13236), .B2(n6236), .C1(n13233), .C2(n15563), .A(
        n3325), .ZN(n3320) );
  OAI222_X1 U4659 ( .A1(n14921), .A2(n13230), .B1(n14857), .B2(n13227), .C1(
        n14889), .C2(n13224), .ZN(n3325) );
  AOI221_X1 U4660 ( .B1(n13236), .B2(n6237), .C1(n13233), .C2(n15562), .A(
        n3288), .ZN(n3283) );
  OAI222_X1 U4661 ( .A1(n14920), .A2(n13230), .B1(n14856), .B2(n13227), .C1(
        n14888), .C2(n13224), .ZN(n3288) );
  AOI221_X1 U4662 ( .B1(n13167), .B2(n6046), .C1(n13164), .C2(n6078), .A(n3260), .ZN(n3253) );
  OAI22_X1 U4663 ( .A1(n15113), .A2(n13161), .B1(n15145), .B2(n13158), .ZN(
        n3260) );
  AOI221_X1 U4664 ( .B1(n13167), .B2(n6047), .C1(n13164), .C2(n6079), .A(n3223), .ZN(n3216) );
  OAI22_X1 U4665 ( .A1(n15112), .A2(n13161), .B1(n15144), .B2(n13158), .ZN(
        n3223) );
  AOI221_X1 U4666 ( .B1(n13167), .B2(n6048), .C1(n13164), .C2(n6080), .A(n3186), .ZN(n3179) );
  OAI22_X1 U4667 ( .A1(n15111), .A2(n13161), .B1(n15143), .B2(n13158), .ZN(
        n3186) );
  AOI221_X1 U4668 ( .B1(n13167), .B2(n6049), .C1(n13164), .C2(n6081), .A(n3147), .ZN(n3124) );
  OAI22_X1 U4669 ( .A1(n15110), .A2(n13161), .B1(n15142), .B2(n13158), .ZN(
        n3147) );
  AOI221_X1 U4670 ( .B1(n12939), .B2(n6075), .C1(n12936), .C2(n6043), .A(n4655), .ZN(n4648) );
  OAI22_X1 U4671 ( .A1(n15148), .A2(n12933), .B1(n15116), .B2(n12930), .ZN(
        n4655) );
  AOI221_X1 U4672 ( .B1(n12939), .B2(n6076), .C1(n12936), .C2(n6044), .A(n4618), .ZN(n4611) );
  OAI22_X1 U4673 ( .A1(n15147), .A2(n12933), .B1(n15115), .B2(n12930), .ZN(
        n4618) );
  AOI221_X1 U4674 ( .B1(n12939), .B2(n6077), .C1(n12936), .C2(n6045), .A(n4581), .ZN(n4574) );
  OAI22_X1 U4675 ( .A1(n15146), .A2(n12933), .B1(n15114), .B2(n12930), .ZN(
        n4581) );
  AOI221_X1 U4676 ( .B1(n12939), .B2(n6078), .C1(n12936), .C2(n6046), .A(n4544), .ZN(n4537) );
  OAI22_X1 U4677 ( .A1(n15145), .A2(n12933), .B1(n15113), .B2(n12930), .ZN(
        n4544) );
  AOI221_X1 U4678 ( .B1(n12939), .B2(n6079), .C1(n12936), .C2(n6047), .A(n4507), .ZN(n4500) );
  OAI22_X1 U4679 ( .A1(n15144), .A2(n12933), .B1(n15112), .B2(n12930), .ZN(
        n4507) );
  AOI221_X1 U4680 ( .B1(n12939), .B2(n6080), .C1(n12936), .C2(n6048), .A(n4470), .ZN(n4463) );
  OAI22_X1 U4681 ( .A1(n15143), .A2(n12933), .B1(n15111), .B2(n12930), .ZN(
        n4470) );
  AOI221_X1 U4682 ( .B1(n12939), .B2(n6081), .C1(n12936), .C2(n6049), .A(n4431), .ZN(n4408) );
  OAI22_X1 U4683 ( .A1(n15142), .A2(n12933), .B1(n15110), .B2(n12930), .ZN(
        n4431) );
  AOI221_X1 U4684 ( .B1(n12992), .B2(n592), .C1(n12989), .C2(n15717), .A(n5128), .ZN(n5121) );
  OAI22_X1 U4685 ( .A1(n14839), .A2(n12986), .B1(n14807), .B2(n12983), .ZN(
        n5128) );
  AOI221_X1 U4686 ( .B1(n12992), .B2(n590), .C1(n12989), .C2(n15716), .A(n5091), .ZN(n5084) );
  OAI22_X1 U4687 ( .A1(n14838), .A2(n12986), .B1(n14806), .B2(n12983), .ZN(
        n5091) );
  AOI221_X1 U4688 ( .B1(n12992), .B2(n588), .C1(n12989), .C2(n15715), .A(n5054), .ZN(n5047) );
  OAI22_X1 U4689 ( .A1(n14837), .A2(n12986), .B1(n14805), .B2(n12983), .ZN(
        n5054) );
  AOI221_X1 U4690 ( .B1(n12992), .B2(n586), .C1(n12989), .C2(n15714), .A(n5017), .ZN(n5010) );
  OAI22_X1 U4691 ( .A1(n14836), .A2(n12986), .B1(n14804), .B2(n12983), .ZN(
        n5017) );
  AOI221_X1 U4692 ( .B1(n12992), .B2(n584), .C1(n12989), .C2(n15713), .A(n4980), .ZN(n4973) );
  OAI22_X1 U4693 ( .A1(n14835), .A2(n12986), .B1(n14803), .B2(n12983), .ZN(
        n4980) );
  AOI221_X1 U4694 ( .B1(n12992), .B2(n582), .C1(n12989), .C2(n15712), .A(n4943), .ZN(n4936) );
  OAI22_X1 U4695 ( .A1(n14834), .A2(n12986), .B1(n14802), .B2(n12983), .ZN(
        n4943) );
  AOI221_X1 U4696 ( .B1(n12992), .B2(n580), .C1(n12989), .C2(n15711), .A(n4906), .ZN(n4899) );
  OAI22_X1 U4697 ( .A1(n14833), .A2(n12986), .B1(n14801), .B2(n12983), .ZN(
        n4906) );
  AOI221_X1 U4698 ( .B1(n12992), .B2(n578), .C1(n12989), .C2(n15710), .A(n4869), .ZN(n4862) );
  OAI22_X1 U4699 ( .A1(n14832), .A2(n12986), .B1(n14800), .B2(n12983), .ZN(
        n4869) );
  AOI221_X1 U4700 ( .B1(n12939), .B2(n6074), .C1(n12936), .C2(n6042), .A(n4692), .ZN(n4685) );
  OAI22_X1 U4701 ( .A1(n15149), .A2(n12933), .B1(n15117), .B2(n12930), .ZN(
        n4692) );
  AOI221_X1 U4702 ( .B1(n13220), .B2(n592), .C1(n13217), .C2(n15717), .A(n3844), .ZN(n3837) );
  OAI22_X1 U4703 ( .A1(n14839), .A2(n13214), .B1(n14807), .B2(n13211), .ZN(
        n3844) );
  AOI221_X1 U4704 ( .B1(n13166), .B2(n6030), .C1(n13163), .C2(n6062), .A(n3852), .ZN(n3845) );
  OAI22_X1 U4705 ( .A1(n15129), .A2(n13160), .B1(n15161), .B2(n13157), .ZN(
        n3852) );
  AOI221_X1 U4706 ( .B1(n13220), .B2(n590), .C1(n13217), .C2(n15716), .A(n3807), .ZN(n3800) );
  OAI22_X1 U4707 ( .A1(n14838), .A2(n13214), .B1(n14806), .B2(n13211), .ZN(
        n3807) );
  AOI221_X1 U4708 ( .B1(n13166), .B2(n6031), .C1(n13163), .C2(n6063), .A(n3815), .ZN(n3808) );
  OAI22_X1 U4709 ( .A1(n15128), .A2(n13160), .B1(n15160), .B2(n13157), .ZN(
        n3815) );
  AOI221_X1 U4710 ( .B1(n13220), .B2(n588), .C1(n13217), .C2(n15715), .A(n3770), .ZN(n3763) );
  OAI22_X1 U4711 ( .A1(n14837), .A2(n13214), .B1(n14805), .B2(n13211), .ZN(
        n3770) );
  AOI221_X1 U4712 ( .B1(n13166), .B2(n6032), .C1(n13163), .C2(n6064), .A(n3778), .ZN(n3771) );
  OAI22_X1 U4713 ( .A1(n15127), .A2(n13160), .B1(n15159), .B2(n13157), .ZN(
        n3778) );
  AOI221_X1 U4714 ( .B1(n13220), .B2(n586), .C1(n13217), .C2(n15714), .A(n3733), .ZN(n3726) );
  OAI22_X1 U4715 ( .A1(n14836), .A2(n13214), .B1(n14804), .B2(n13211), .ZN(
        n3733) );
  AOI221_X1 U4716 ( .B1(n13166), .B2(n6033), .C1(n13163), .C2(n6065), .A(n3741), .ZN(n3734) );
  OAI22_X1 U4717 ( .A1(n15126), .A2(n13160), .B1(n15158), .B2(n13157), .ZN(
        n3741) );
  AOI221_X1 U4718 ( .B1(n13220), .B2(n584), .C1(n13217), .C2(n15713), .A(n3696), .ZN(n3689) );
  OAI22_X1 U4719 ( .A1(n14835), .A2(n13214), .B1(n14803), .B2(n13211), .ZN(
        n3696) );
  AOI221_X1 U4720 ( .B1(n13166), .B2(n6034), .C1(n13163), .C2(n6066), .A(n3704), .ZN(n3697) );
  OAI22_X1 U4721 ( .A1(n15125), .A2(n13160), .B1(n15157), .B2(n13157), .ZN(
        n3704) );
  AOI221_X1 U4722 ( .B1(n13220), .B2(n582), .C1(n13217), .C2(n15712), .A(n3659), .ZN(n3652) );
  OAI22_X1 U4723 ( .A1(n14834), .A2(n13214), .B1(n14802), .B2(n13211), .ZN(
        n3659) );
  AOI221_X1 U4724 ( .B1(n13166), .B2(n6035), .C1(n13163), .C2(n6067), .A(n3667), .ZN(n3660) );
  OAI22_X1 U4725 ( .A1(n15124), .A2(n13160), .B1(n15156), .B2(n13157), .ZN(
        n3667) );
  AOI221_X1 U4726 ( .B1(n13220), .B2(n580), .C1(n13217), .C2(n15711), .A(n3622), .ZN(n3615) );
  OAI22_X1 U4727 ( .A1(n14833), .A2(n13214), .B1(n14801), .B2(n13211), .ZN(
        n3622) );
  AOI221_X1 U4728 ( .B1(n13166), .B2(n6036), .C1(n13163), .C2(n6068), .A(n3630), .ZN(n3623) );
  OAI22_X1 U4729 ( .A1(n15123), .A2(n13160), .B1(n15155), .B2(n13157), .ZN(
        n3630) );
  AOI221_X1 U4730 ( .B1(n13220), .B2(n578), .C1(n13217), .C2(n15710), .A(n3585), .ZN(n3578) );
  OAI22_X1 U4731 ( .A1(n14832), .A2(n13214), .B1(n14800), .B2(n13211), .ZN(
        n3585) );
  AOI221_X1 U4732 ( .B1(n13166), .B2(n6037), .C1(n13163), .C2(n6069), .A(n3593), .ZN(n3586) );
  OAI22_X1 U4733 ( .A1(n15122), .A2(n13160), .B1(n15154), .B2(n13157), .ZN(
        n3593) );
  AOI221_X1 U4734 ( .B1(n13166), .B2(n6038), .C1(n13163), .C2(n6070), .A(n3556), .ZN(n3549) );
  OAI22_X1 U4735 ( .A1(n15121), .A2(n13160), .B1(n15153), .B2(n13157), .ZN(
        n3556) );
  AOI221_X1 U4736 ( .B1(n13166), .B2(n6039), .C1(n13163), .C2(n6071), .A(n3519), .ZN(n3512) );
  OAI22_X1 U4737 ( .A1(n15120), .A2(n13160), .B1(n15152), .B2(n13157), .ZN(
        n3519) );
  AOI221_X1 U4738 ( .B1(n13166), .B2(n6040), .C1(n13163), .C2(n6072), .A(n3482), .ZN(n3475) );
  OAI22_X1 U4739 ( .A1(n15119), .A2(n13160), .B1(n15151), .B2(n13157), .ZN(
        n3482) );
  AOI221_X1 U4740 ( .B1(n13166), .B2(n6041), .C1(n13163), .C2(n6073), .A(n3445), .ZN(n3438) );
  OAI22_X1 U4741 ( .A1(n15118), .A2(n13160), .B1(n15150), .B2(n13157), .ZN(
        n3445) );
  AOI221_X1 U4742 ( .B1(n13167), .B2(n6043), .C1(n13164), .C2(n6075), .A(n3371), .ZN(n3364) );
  OAI22_X1 U4743 ( .A1(n15116), .A2(n13161), .B1(n15148), .B2(n13158), .ZN(
        n3371) );
  AOI221_X1 U4744 ( .B1(n13167), .B2(n6044), .C1(n13164), .C2(n6076), .A(n3334), .ZN(n3327) );
  OAI22_X1 U4745 ( .A1(n15115), .A2(n13161), .B1(n15147), .B2(n13158), .ZN(
        n3334) );
  AOI221_X1 U4746 ( .B1(n13167), .B2(n6045), .C1(n13164), .C2(n6077), .A(n3297), .ZN(n3290) );
  OAI22_X1 U4747 ( .A1(n15114), .A2(n13161), .B1(n15146), .B2(n13158), .ZN(
        n3297) );
  AOI221_X1 U4748 ( .B1(n13221), .B2(n15730), .C1(n13218), .C2(n98), .A(n3121), 
        .ZN(n3098) );
  OAI22_X1 U4749 ( .A1(n14820), .A2(n13215), .B1(n14788), .B2(n13212), .ZN(
        n3121) );
  AOI221_X1 U4750 ( .B1(n12993), .B2(n15730), .C1(n12990), .C2(n98), .A(n4405), 
        .ZN(n4382) );
  OAI22_X1 U4751 ( .A1(n14820), .A2(n12987), .B1(n14788), .B2(n12984), .ZN(
        n4405) );
  OAI22_X1 U4752 ( .A1(n12645), .A2(n13323), .B1(n5667), .B2(n13320), .ZN(
        n3236) );
  OAI22_X1 U4753 ( .A1(n12646), .A2(n13323), .B1(n5677), .B2(n13320), .ZN(
        n3199) );
  OAI22_X1 U4754 ( .A1(n12647), .A2(n13323), .B1(n5687), .B2(n13320), .ZN(
        n3162) );
  OAI22_X1 U4755 ( .A1(n12648), .A2(n13323), .B1(n5697), .B2(n13320), .ZN(
        n3069) );
  OAI22_X1 U4756 ( .A1(n6803), .A2(n13095), .B1(n6931), .B2(n13092), .ZN(n4631) );
  OAI22_X1 U4757 ( .A1(n6804), .A2(n13095), .B1(n6932), .B2(n13092), .ZN(n4594) );
  OAI22_X1 U4758 ( .A1(n6805), .A2(n13095), .B1(n6933), .B2(n13092), .ZN(n4557) );
  OAI22_X1 U4759 ( .A1(n6806), .A2(n13095), .B1(n6934), .B2(n13092), .ZN(n4520) );
  OAI22_X1 U4760 ( .A1(n6807), .A2(n13095), .B1(n6935), .B2(n13092), .ZN(n4483) );
  OAI22_X1 U4761 ( .A1(n6808), .A2(n13095), .B1(n6936), .B2(n13092), .ZN(n4446) );
  OAI22_X1 U4762 ( .A1(n6809), .A2(n13095), .B1(n6937), .B2(n13092), .ZN(n4353) );
  OAI22_X1 U4763 ( .A1(n6802), .A2(n13095), .B1(n6930), .B2(n13092), .ZN(n4668) );
  OAI22_X1 U4764 ( .A1(n12649), .A2(n13323), .B1(n5627), .B2(n13320), .ZN(
        n3384) );
  OAI22_X1 U4765 ( .A1(n12650), .A2(n13323), .B1(n5637), .B2(n13320), .ZN(
        n3347) );
  OAI22_X1 U4766 ( .A1(n12651), .A2(n13323), .B1(n5647), .B2(n13320), .ZN(
        n3310) );
  OAI22_X1 U4767 ( .A1(n12652), .A2(n13323), .B1(n5657), .B2(n13320), .ZN(
        n3273) );
  OAI22_X1 U4768 ( .A1(n12653), .A2(n13350), .B1(n5665), .B2(n13347), .ZN(
        n3234) );
  OAI22_X1 U4769 ( .A1(n12654), .A2(n13350), .B1(n5675), .B2(n13347), .ZN(
        n3197) );
  OAI22_X1 U4770 ( .A1(n12655), .A2(n13350), .B1(n5685), .B2(n13347), .ZN(
        n3160) );
  OAI22_X1 U4771 ( .A1(n12656), .A2(n13350), .B1(n5695), .B2(n13347), .ZN(
        n3058) );
  OAI22_X1 U4772 ( .A1(n6787), .A2(n13122), .B1(n6915), .B2(n13119), .ZN(n4629) );
  OAI22_X1 U4773 ( .A1(n6788), .A2(n13122), .B1(n6916), .B2(n13119), .ZN(n4592) );
  OAI22_X1 U4774 ( .A1(n6789), .A2(n13122), .B1(n6917), .B2(n13119), .ZN(n4555) );
  OAI22_X1 U4775 ( .A1(n6790), .A2(n13122), .B1(n6918), .B2(n13119), .ZN(n4518) );
  OAI22_X1 U4776 ( .A1(n6791), .A2(n13122), .B1(n6919), .B2(n13119), .ZN(n4481) );
  OAI22_X1 U4777 ( .A1(n6792), .A2(n13122), .B1(n6920), .B2(n13119), .ZN(n4444) );
  OAI22_X1 U4778 ( .A1(n6793), .A2(n13122), .B1(n6921), .B2(n13119), .ZN(n4342) );
  OAI22_X1 U4779 ( .A1(n6786), .A2(n13122), .B1(n6914), .B2(n13119), .ZN(n4666) );
  OAI22_X1 U4780 ( .A1(n12657), .A2(n13350), .B1(n5625), .B2(n13347), .ZN(
        n3382) );
  OAI22_X1 U4781 ( .A1(n12658), .A2(n13350), .B1(n5635), .B2(n13347), .ZN(
        n3345) );
  OAI22_X1 U4782 ( .A1(n12659), .A2(n13350), .B1(n5645), .B2(n13347), .ZN(
        n3308) );
  OAI22_X1 U4783 ( .A1(n12660), .A2(n13350), .B1(n5655), .B2(n13347), .ZN(
        n3271) );
  AOI221_X1 U4784 ( .B1(n13020), .B2(n6170), .C1(n13017), .C2(n15619), .A(
        n4682), .ZN(n4679) );
  OAI22_X1 U4785 ( .A1(n14956), .A2(n13014), .B1(n15930), .B2(n13011), .ZN(
        n4682) );
  AOI221_X1 U4786 ( .B1(n13248), .B2(n6170), .C1(n13245), .C2(n15619), .A(
        n3398), .ZN(n3395) );
  OAI22_X1 U4787 ( .A1(n14956), .A2(n13242), .B1(n15930), .B2(n13239), .ZN(
        n3398) );
  AOI221_X1 U4788 ( .B1(n13167), .B2(n6042), .C1(n13164), .C2(n6074), .A(n3408), .ZN(n3401) );
  OAI22_X1 U4789 ( .A1(n15117), .A2(n13161), .B1(n15149), .B2(n13158), .ZN(
        n3408) );
  OAI22_X1 U4790 ( .A1(n6870), .A2(n13120), .B1(n710), .B2(n13117), .ZN(n5670)
         );
  OAI22_X1 U4791 ( .A1(n6830), .A2(n13093), .B1(n711), .B2(n13090), .ZN(n5680)
         );
  OAI22_X1 U4792 ( .A1(n6871), .A2(n13120), .B1(n707), .B2(n13117), .ZN(n5598)
         );
  OAI22_X1 U4793 ( .A1(n6831), .A2(n13093), .B1(n708), .B2(n13090), .ZN(n5600)
         );
  OAI22_X1 U4794 ( .A1(n6872), .A2(n13120), .B1(n704), .B2(n13117), .ZN(n5536)
         );
  OAI22_X1 U4795 ( .A1(n6832), .A2(n13093), .B1(n705), .B2(n13090), .ZN(n5539)
         );
  OAI22_X1 U4796 ( .A1(n6873), .A2(n13120), .B1(n701), .B2(n13117), .ZN(n5474)
         );
  OAI22_X1 U4797 ( .A1(n6833), .A2(n13093), .B1(n702), .B2(n13090), .ZN(n5478)
         );
  OAI22_X1 U4798 ( .A1(n6874), .A2(n13120), .B1(n698), .B2(n13117), .ZN(n5418)
         );
  OAI22_X1 U4799 ( .A1(n6834), .A2(n13093), .B1(n699), .B2(n13090), .ZN(n5420)
         );
  OAI22_X1 U4800 ( .A1(n6875), .A2(n13120), .B1(n695), .B2(n13117), .ZN(n5369)
         );
  OAI22_X1 U4801 ( .A1(n6835), .A2(n13093), .B1(n696), .B2(n13090), .ZN(n5371)
         );
  OAI22_X1 U4802 ( .A1(n6876), .A2(n13120), .B1(n692), .B2(n13117), .ZN(n5332)
         );
  OAI22_X1 U4803 ( .A1(n6836), .A2(n13093), .B1(n693), .B2(n13090), .ZN(n5334)
         );
  OAI22_X1 U4804 ( .A1(n6877), .A2(n13120), .B1(n689), .B2(n13117), .ZN(n5295)
         );
  OAI22_X1 U4805 ( .A1(n6837), .A2(n13093), .B1(n690), .B2(n13090), .ZN(n5297)
         );
  OAI22_X1 U4806 ( .A1(n6878), .A2(n13120), .B1(n686), .B2(n13117), .ZN(n5258)
         );
  OAI22_X1 U4807 ( .A1(n6838), .A2(n13093), .B1(n687), .B2(n13090), .ZN(n5260)
         );
  OAI22_X1 U4808 ( .A1(n6879), .A2(n13120), .B1(n683), .B2(n13117), .ZN(n5221)
         );
  OAI22_X1 U4809 ( .A1(n6839), .A2(n13093), .B1(n684), .B2(n13090), .ZN(n5223)
         );
  OAI22_X1 U4810 ( .A1(n6880), .A2(n13120), .B1(n680), .B2(n13117), .ZN(n5184)
         );
  OAI22_X1 U4811 ( .A1(n6840), .A2(n13093), .B1(n681), .B2(n13090), .ZN(n5186)
         );
  OAI22_X1 U4812 ( .A1(n6881), .A2(n13120), .B1(n677), .B2(n13117), .ZN(n5147)
         );
  OAI22_X1 U4813 ( .A1(n6841), .A2(n13093), .B1(n678), .B2(n13090), .ZN(n5149)
         );
  OAI22_X1 U4814 ( .A1(n6882), .A2(n13121), .B1(n674), .B2(n13118), .ZN(n5110)
         );
  OAI22_X1 U4815 ( .A1(n6883), .A2(n13094), .B1(n675), .B2(n13091), .ZN(n5112)
         );
  OAI22_X1 U4816 ( .A1(n6884), .A2(n13121), .B1(n671), .B2(n13118), .ZN(n5073)
         );
  OAI22_X1 U4817 ( .A1(n6885), .A2(n13094), .B1(n672), .B2(n13091), .ZN(n5075)
         );
  OAI22_X1 U4818 ( .A1(n6886), .A2(n13121), .B1(n668), .B2(n13118), .ZN(n5036)
         );
  OAI22_X1 U4819 ( .A1(n6887), .A2(n13094), .B1(n669), .B2(n13091), .ZN(n5038)
         );
  OAI22_X1 U4820 ( .A1(n6888), .A2(n13121), .B1(n665), .B2(n13118), .ZN(n4999)
         );
  OAI22_X1 U4821 ( .A1(n6889), .A2(n13094), .B1(n666), .B2(n13091), .ZN(n5001)
         );
  OAI22_X1 U4822 ( .A1(n6890), .A2(n13121), .B1(n662), .B2(n13118), .ZN(n4962)
         );
  OAI22_X1 U4823 ( .A1(n6794), .A2(n13094), .B1(n6922), .B2(n13091), .ZN(n4964) );
  OAI22_X1 U4824 ( .A1(n6891), .A2(n13121), .B1(n659), .B2(n13118), .ZN(n4925)
         );
  OAI22_X1 U4825 ( .A1(n6795), .A2(n13094), .B1(n6923), .B2(n13091), .ZN(n4927) );
  OAI22_X1 U4826 ( .A1(n6892), .A2(n13121), .B1(n656), .B2(n13118), .ZN(n4888)
         );
  OAI22_X1 U4827 ( .A1(n6796), .A2(n13094), .B1(n6924), .B2(n13091), .ZN(n4890) );
  OAI22_X1 U4828 ( .A1(n6893), .A2(n13121), .B1(n653), .B2(n13118), .ZN(n4851)
         );
  OAI22_X1 U4829 ( .A1(n6797), .A2(n13094), .B1(n6925), .B2(n13091), .ZN(n4853) );
  OAI22_X1 U4830 ( .A1(n6810), .A2(n13121), .B1(n6938), .B2(n13118), .ZN(n4814) );
  OAI22_X1 U4831 ( .A1(n6798), .A2(n13094), .B1(n6926), .B2(n13091), .ZN(n4816) );
  OAI22_X1 U4832 ( .A1(n6811), .A2(n13121), .B1(n6939), .B2(n13118), .ZN(n4777) );
  OAI22_X1 U4833 ( .A1(n6799), .A2(n13094), .B1(n6927), .B2(n13091), .ZN(n4779) );
  OAI22_X1 U4834 ( .A1(n6812), .A2(n13121), .B1(n6940), .B2(n13118), .ZN(n4740) );
  OAI22_X1 U4835 ( .A1(n6800), .A2(n13094), .B1(n6928), .B2(n13091), .ZN(n4742) );
  OAI22_X1 U4836 ( .A1(n6813), .A2(n13121), .B1(n6941), .B2(n13118), .ZN(n4703) );
  OAI22_X1 U4837 ( .A1(n6801), .A2(n13094), .B1(n6929), .B2(n13091), .ZN(n4705) );
  OAI22_X1 U4838 ( .A1(n12661), .A2(n13348), .B1(n5385), .B2(n13345), .ZN(
        n4277) );
  OAI22_X1 U4839 ( .A1(n12662), .A2(n13321), .B1(n5387), .B2(n13318), .ZN(
        n4283) );
  OAI22_X1 U4840 ( .A1(n12663), .A2(n13348), .B1(n5395), .B2(n13345), .ZN(
        n4233) );
  OAI22_X1 U4841 ( .A1(n12664), .A2(n13321), .B1(n5397), .B2(n13318), .ZN(
        n4235) );
  OAI22_X1 U4842 ( .A1(n12665), .A2(n13348), .B1(n5405), .B2(n13345), .ZN(
        n4196) );
  OAI22_X1 U4843 ( .A1(n12666), .A2(n13321), .B1(n5407), .B2(n13318), .ZN(
        n4198) );
  OAI22_X1 U4844 ( .A1(n12667), .A2(n13348), .B1(n5415), .B2(n13345), .ZN(
        n4159) );
  OAI22_X1 U4845 ( .A1(n12668), .A2(n13321), .B1(n5417), .B2(n13318), .ZN(
        n4161) );
  OAI22_X1 U4846 ( .A1(n12669), .A2(n13348), .B1(n5425), .B2(n13345), .ZN(
        n4122) );
  OAI22_X1 U4847 ( .A1(n12670), .A2(n13321), .B1(n5427), .B2(n13318), .ZN(
        n4124) );
  OAI22_X1 U4848 ( .A1(n12671), .A2(n13348), .B1(n5435), .B2(n13345), .ZN(
        n4085) );
  OAI22_X1 U4849 ( .A1(n12672), .A2(n13321), .B1(n5437), .B2(n13318), .ZN(
        n4087) );
  OAI22_X1 U4850 ( .A1(n12673), .A2(n13348), .B1(n5445), .B2(n13345), .ZN(
        n4048) );
  OAI22_X1 U4851 ( .A1(n12674), .A2(n13321), .B1(n5447), .B2(n13318), .ZN(
        n4050) );
  OAI22_X1 U4852 ( .A1(n12675), .A2(n13348), .B1(n5455), .B2(n13345), .ZN(
        n4011) );
  OAI22_X1 U4853 ( .A1(n12676), .A2(n13321), .B1(n5457), .B2(n13318), .ZN(
        n4013) );
  OAI22_X1 U4854 ( .A1(n12677), .A2(n13348), .B1(n5465), .B2(n13345), .ZN(
        n3974) );
  OAI22_X1 U4855 ( .A1(n12678), .A2(n13321), .B1(n5467), .B2(n13318), .ZN(
        n3976) );
  OAI22_X1 U4856 ( .A1(n12679), .A2(n13348), .B1(n5475), .B2(n13345), .ZN(
        n3937) );
  OAI22_X1 U4857 ( .A1(n12680), .A2(n13321), .B1(n5477), .B2(n13318), .ZN(
        n3939) );
  OAI22_X1 U4858 ( .A1(n12681), .A2(n13348), .B1(n5485), .B2(n13345), .ZN(
        n3900) );
  OAI22_X1 U4859 ( .A1(n12682), .A2(n13321), .B1(n5487), .B2(n13318), .ZN(
        n3902) );
  OAI22_X1 U4860 ( .A1(n12683), .A2(n13348), .B1(n5495), .B2(n13345), .ZN(
        n3863) );
  OAI22_X1 U4861 ( .A1(n12684), .A2(n13321), .B1(n5497), .B2(n13318), .ZN(
        n3865) );
  OAI22_X1 U4862 ( .A1(n12685), .A2(n13349), .B1(n5505), .B2(n13346), .ZN(
        n3826) );
  OAI22_X1 U4863 ( .A1(n12686), .A2(n13322), .B1(n5507), .B2(n13319), .ZN(
        n3828) );
  OAI22_X1 U4864 ( .A1(n12687), .A2(n13349), .B1(n5515), .B2(n13346), .ZN(
        n3789) );
  OAI22_X1 U4865 ( .A1(n12688), .A2(n13322), .B1(n5517), .B2(n13319), .ZN(
        n3791) );
  OAI22_X1 U4866 ( .A1(n12689), .A2(n13349), .B1(n5525), .B2(n13346), .ZN(
        n3752) );
  OAI22_X1 U4867 ( .A1(n12690), .A2(n13322), .B1(n5527), .B2(n13319), .ZN(
        n3754) );
  OAI22_X1 U4868 ( .A1(n12691), .A2(n13349), .B1(n5535), .B2(n13346), .ZN(
        n3715) );
  OAI22_X1 U4869 ( .A1(n12692), .A2(n13322), .B1(n5537), .B2(n13319), .ZN(
        n3717) );
  OAI22_X1 U4870 ( .A1(n12693), .A2(n13349), .B1(n5545), .B2(n13346), .ZN(
        n3678) );
  OAI22_X1 U4871 ( .A1(n12694), .A2(n13322), .B1(n5547), .B2(n13319), .ZN(
        n3680) );
  OAI22_X1 U4872 ( .A1(n12695), .A2(n13349), .B1(n5555), .B2(n13346), .ZN(
        n3641) );
  OAI22_X1 U4873 ( .A1(n12696), .A2(n13322), .B1(n5557), .B2(n13319), .ZN(
        n3643) );
  OAI22_X1 U4874 ( .A1(n12697), .A2(n13349), .B1(n5565), .B2(n13346), .ZN(
        n3604) );
  OAI22_X1 U4875 ( .A1(n12698), .A2(n13322), .B1(n5567), .B2(n13319), .ZN(
        n3606) );
  OAI22_X1 U4876 ( .A1(n12699), .A2(n13349), .B1(n5575), .B2(n13346), .ZN(
        n3567) );
  OAI22_X1 U4877 ( .A1(n12700), .A2(n13322), .B1(n5577), .B2(n13319), .ZN(
        n3569) );
  OAI22_X1 U4878 ( .A1(n12701), .A2(n13349), .B1(n5585), .B2(n13346), .ZN(
        n3530) );
  OAI22_X1 U4879 ( .A1(n12702), .A2(n13322), .B1(n5587), .B2(n13319), .ZN(
        n3532) );
  OAI22_X1 U4880 ( .A1(n12703), .A2(n13349), .B1(n5595), .B2(n13346), .ZN(
        n3493) );
  OAI22_X1 U4881 ( .A1(n12704), .A2(n13322), .B1(n5597), .B2(n13319), .ZN(
        n3495) );
  OAI22_X1 U4882 ( .A1(n12705), .A2(n13349), .B1(n5605), .B2(n13346), .ZN(
        n3456) );
  OAI22_X1 U4883 ( .A1(n12706), .A2(n13322), .B1(n5607), .B2(n13319), .ZN(
        n3458) );
  OAI22_X1 U4884 ( .A1(n12707), .A2(n13349), .B1(n5615), .B2(n13346), .ZN(
        n3419) );
  OAI22_X1 U4885 ( .A1(n12708), .A2(n13322), .B1(n5617), .B2(n13319), .ZN(
        n3421) );
  AOI221_X1 U4886 ( .B1(n12991), .B2(n616), .C1(n12988), .C2(n15729), .A(n5718), .ZN(n5700) );
  OAI22_X1 U4887 ( .A1(n14851), .A2(n12985), .B1(n14819), .B2(n12982), .ZN(
        n5718) );
  AOI221_X1 U4888 ( .B1(n12937), .B2(n6050), .C1(n12934), .C2(n6018), .A(n5736), .ZN(n5720) );
  OAI22_X1 U4889 ( .A1(n15173), .A2(n12931), .B1(n15141), .B2(n12928), .ZN(
        n5736) );
  AOI221_X1 U4890 ( .B1(n12991), .B2(n614), .C1(n12988), .C2(n15728), .A(n5628), .ZN(n5616) );
  OAI22_X1 U4891 ( .A1(n14850), .A2(n12985), .B1(n14818), .B2(n12982), .ZN(
        n5628) );
  AOI221_X1 U4892 ( .B1(n12937), .B2(n6051), .C1(n12934), .C2(n6019), .A(n5640), .ZN(n5629) );
  OAI22_X1 U4893 ( .A1(n15172), .A2(n12931), .B1(n15140), .B2(n12928), .ZN(
        n5640) );
  AOI221_X1 U4894 ( .B1(n12991), .B2(n612), .C1(n12988), .C2(n15727), .A(n5566), .ZN(n5554) );
  OAI22_X1 U4895 ( .A1(n14849), .A2(n12985), .B1(n14817), .B2(n12982), .ZN(
        n5566) );
  AOI221_X1 U4896 ( .B1(n12937), .B2(n6052), .C1(n12934), .C2(n6020), .A(n5579), .ZN(n5568) );
  OAI22_X1 U4897 ( .A1(n15171), .A2(n12931), .B1(n15139), .B2(n12928), .ZN(
        n5579) );
  AOI221_X1 U4898 ( .B1(n12991), .B2(n610), .C1(n12988), .C2(n15726), .A(n5504), .ZN(n5491) );
  OAI22_X1 U4899 ( .A1(n14848), .A2(n12985), .B1(n14816), .B2(n12982), .ZN(
        n5504) );
  AOI221_X1 U4900 ( .B1(n12937), .B2(n6053), .C1(n12934), .C2(n6021), .A(n5518), .ZN(n5506) );
  OAI22_X1 U4901 ( .A1(n15170), .A2(n12931), .B1(n15138), .B2(n12928), .ZN(
        n5518) );
  AOI221_X1 U4902 ( .B1(n12991), .B2(n608), .C1(n12988), .C2(n15725), .A(n5442), .ZN(n5432) );
  OAI22_X1 U4903 ( .A1(n14847), .A2(n12985), .B1(n14815), .B2(n12982), .ZN(
        n5442) );
  AOI221_X1 U4904 ( .B1(n12937), .B2(n6054), .C1(n12934), .C2(n6022), .A(n5456), .ZN(n5444) );
  OAI22_X1 U4905 ( .A1(n15169), .A2(n12931), .B1(n15137), .B2(n12928), .ZN(
        n5456) );
  AOI221_X1 U4906 ( .B1(n12991), .B2(n606), .C1(n12988), .C2(n15724), .A(n5390), .ZN(n5380) );
  OAI22_X1 U4907 ( .A1(n14846), .A2(n12985), .B1(n14814), .B2(n12982), .ZN(
        n5390) );
  AOI221_X1 U4908 ( .B1(n12937), .B2(n6055), .C1(n12934), .C2(n6023), .A(n5401), .ZN(n5391) );
  OAI22_X1 U4909 ( .A1(n15168), .A2(n12931), .B1(n15136), .B2(n12928), .ZN(
        n5401) );
  AOI221_X1 U4910 ( .B1(n12991), .B2(n604), .C1(n12988), .C2(n15723), .A(n5350), .ZN(n5343) );
  OAI22_X1 U4911 ( .A1(n14845), .A2(n12985), .B1(n14813), .B2(n12982), .ZN(
        n5350) );
  AOI221_X1 U4912 ( .B1(n12937), .B2(n6056), .C1(n12934), .C2(n6024), .A(n5358), .ZN(n5351) );
  OAI22_X1 U4913 ( .A1(n15167), .A2(n12931), .B1(n15135), .B2(n12928), .ZN(
        n5358) );
  AOI221_X1 U4914 ( .B1(n12991), .B2(n602), .C1(n12988), .C2(n15722), .A(n5313), .ZN(n5306) );
  OAI22_X1 U4915 ( .A1(n14844), .A2(n12985), .B1(n14812), .B2(n12982), .ZN(
        n5313) );
  AOI221_X1 U4916 ( .B1(n12937), .B2(n6057), .C1(n12934), .C2(n6025), .A(n5321), .ZN(n5314) );
  OAI22_X1 U4917 ( .A1(n15166), .A2(n12931), .B1(n15134), .B2(n12928), .ZN(
        n5321) );
  AOI221_X1 U4918 ( .B1(n12991), .B2(n600), .C1(n12988), .C2(n15721), .A(n5276), .ZN(n5269) );
  OAI22_X1 U4919 ( .A1(n14843), .A2(n12985), .B1(n14811), .B2(n12982), .ZN(
        n5276) );
  AOI221_X1 U4920 ( .B1(n12937), .B2(n6058), .C1(n12934), .C2(n6026), .A(n5284), .ZN(n5277) );
  OAI22_X1 U4921 ( .A1(n15165), .A2(n12931), .B1(n15133), .B2(n12928), .ZN(
        n5284) );
  AOI221_X1 U4922 ( .B1(n12991), .B2(n598), .C1(n12988), .C2(n15720), .A(n5239), .ZN(n5232) );
  OAI22_X1 U4923 ( .A1(n14842), .A2(n12985), .B1(n14810), .B2(n12982), .ZN(
        n5239) );
  AOI221_X1 U4924 ( .B1(n12937), .B2(n6059), .C1(n12934), .C2(n6027), .A(n5247), .ZN(n5240) );
  OAI22_X1 U4925 ( .A1(n15164), .A2(n12931), .B1(n15132), .B2(n12928), .ZN(
        n5247) );
  AOI221_X1 U4926 ( .B1(n12991), .B2(n596), .C1(n12988), .C2(n15719), .A(n5202), .ZN(n5195) );
  OAI22_X1 U4927 ( .A1(n14841), .A2(n12985), .B1(n14809), .B2(n12982), .ZN(
        n5202) );
  AOI221_X1 U4928 ( .B1(n12937), .B2(n6060), .C1(n12934), .C2(n6028), .A(n5210), .ZN(n5203) );
  OAI22_X1 U4929 ( .A1(n15163), .A2(n12931), .B1(n15131), .B2(n12928), .ZN(
        n5210) );
  AOI221_X1 U4930 ( .B1(n12991), .B2(n594), .C1(n12988), .C2(n15718), .A(n5165), .ZN(n5158) );
  OAI22_X1 U4931 ( .A1(n14840), .A2(n12985), .B1(n14808), .B2(n12982), .ZN(
        n5165) );
  AOI221_X1 U4932 ( .B1(n12937), .B2(n6061), .C1(n12934), .C2(n6029), .A(n5173), .ZN(n5166) );
  OAI22_X1 U4933 ( .A1(n15162), .A2(n12931), .B1(n15130), .B2(n12928), .ZN(
        n5173) );
  AOI221_X1 U4934 ( .B1(n12938), .B2(n6062), .C1(n12935), .C2(n6030), .A(n5136), .ZN(n5129) );
  OAI22_X1 U4935 ( .A1(n15161), .A2(n12932), .B1(n15129), .B2(n12929), .ZN(
        n5136) );
  AOI221_X1 U4936 ( .B1(n12938), .B2(n6063), .C1(n12935), .C2(n6031), .A(n5099), .ZN(n5092) );
  OAI22_X1 U4937 ( .A1(n15160), .A2(n12932), .B1(n15128), .B2(n12929), .ZN(
        n5099) );
  AOI221_X1 U4938 ( .B1(n12938), .B2(n6064), .C1(n12935), .C2(n6032), .A(n5062), .ZN(n5055) );
  OAI22_X1 U4939 ( .A1(n15159), .A2(n12932), .B1(n15127), .B2(n12929), .ZN(
        n5062) );
  AOI221_X1 U4940 ( .B1(n12938), .B2(n6065), .C1(n12935), .C2(n6033), .A(n5025), .ZN(n5018) );
  OAI22_X1 U4941 ( .A1(n15158), .A2(n12932), .B1(n15126), .B2(n12929), .ZN(
        n5025) );
  AOI221_X1 U4942 ( .B1(n12938), .B2(n6066), .C1(n12935), .C2(n6034), .A(n4988), .ZN(n4981) );
  OAI22_X1 U4943 ( .A1(n15157), .A2(n12932), .B1(n15125), .B2(n12929), .ZN(
        n4988) );
  AOI221_X1 U4944 ( .B1(n12938), .B2(n6067), .C1(n12935), .C2(n6035), .A(n4951), .ZN(n4944) );
  OAI22_X1 U4945 ( .A1(n15156), .A2(n12932), .B1(n15124), .B2(n12929), .ZN(
        n4951) );
  AOI221_X1 U4946 ( .B1(n12938), .B2(n6068), .C1(n12935), .C2(n6036), .A(n4914), .ZN(n4907) );
  OAI22_X1 U4947 ( .A1(n15155), .A2(n12932), .B1(n15123), .B2(n12929), .ZN(
        n4914) );
  AOI221_X1 U4948 ( .B1(n12938), .B2(n6069), .C1(n12935), .C2(n6037), .A(n4877), .ZN(n4870) );
  OAI22_X1 U4949 ( .A1(n15154), .A2(n12932), .B1(n15122), .B2(n12929), .ZN(
        n4877) );
  AOI221_X1 U4950 ( .B1(n12938), .B2(n6070), .C1(n12935), .C2(n6038), .A(n4840), .ZN(n4833) );
  OAI22_X1 U4951 ( .A1(n15153), .A2(n12932), .B1(n15121), .B2(n12929), .ZN(
        n4840) );
  AOI221_X1 U4952 ( .B1(n12938), .B2(n6071), .C1(n12935), .C2(n6039), .A(n4803), .ZN(n4796) );
  OAI22_X1 U4953 ( .A1(n15152), .A2(n12932), .B1(n15120), .B2(n12929), .ZN(
        n4803) );
  AOI221_X1 U4954 ( .B1(n12938), .B2(n6072), .C1(n12935), .C2(n6040), .A(n4766), .ZN(n4759) );
  OAI22_X1 U4955 ( .A1(n15151), .A2(n12932), .B1(n15119), .B2(n12929), .ZN(
        n4766) );
  AOI221_X1 U4956 ( .B1(n12938), .B2(n6073), .C1(n12935), .C2(n6041), .A(n4729), .ZN(n4722) );
  OAI22_X1 U4957 ( .A1(n15150), .A2(n12932), .B1(n15118), .B2(n12929), .ZN(
        n4729) );
  AOI221_X1 U4958 ( .B1(n13219), .B2(n616), .C1(n13216), .C2(n15729), .A(n4303), .ZN(n4294) );
  OAI22_X1 U4959 ( .A1(n14851), .A2(n13213), .B1(n14819), .B2(n13210), .ZN(
        n4303) );
  AOI221_X1 U4960 ( .B1(n13165), .B2(n6018), .C1(n13162), .C2(n6050), .A(n4312), .ZN(n4304) );
  OAI22_X1 U4961 ( .A1(n15141), .A2(n13159), .B1(n15173), .B2(n13156), .ZN(
        n4312) );
  AOI221_X1 U4962 ( .B1(n13219), .B2(n614), .C1(n13216), .C2(n15728), .A(n4251), .ZN(n4244) );
  OAI22_X1 U4963 ( .A1(n14850), .A2(n13213), .B1(n14818), .B2(n13210), .ZN(
        n4251) );
  AOI221_X1 U4964 ( .B1(n13165), .B2(n6019), .C1(n13162), .C2(n6051), .A(n4259), .ZN(n4252) );
  OAI22_X1 U4965 ( .A1(n15140), .A2(n13159), .B1(n15172), .B2(n13156), .ZN(
        n4259) );
  AOI221_X1 U4966 ( .B1(n13219), .B2(n612), .C1(n13216), .C2(n15727), .A(n4214), .ZN(n4207) );
  OAI22_X1 U4967 ( .A1(n14849), .A2(n13213), .B1(n14817), .B2(n13210), .ZN(
        n4214) );
  AOI221_X1 U4968 ( .B1(n13165), .B2(n6020), .C1(n13162), .C2(n6052), .A(n4222), .ZN(n4215) );
  OAI22_X1 U4969 ( .A1(n15139), .A2(n13159), .B1(n15171), .B2(n13156), .ZN(
        n4222) );
  AOI221_X1 U4970 ( .B1(n13219), .B2(n610), .C1(n13216), .C2(n15726), .A(n4177), .ZN(n4170) );
  OAI22_X1 U4971 ( .A1(n14848), .A2(n13213), .B1(n14816), .B2(n13210), .ZN(
        n4177) );
  AOI221_X1 U4972 ( .B1(n13165), .B2(n6021), .C1(n13162), .C2(n6053), .A(n4185), .ZN(n4178) );
  OAI22_X1 U4973 ( .A1(n15138), .A2(n13159), .B1(n15170), .B2(n13156), .ZN(
        n4185) );
  AOI221_X1 U4974 ( .B1(n13219), .B2(n608), .C1(n13216), .C2(n15725), .A(n4140), .ZN(n4133) );
  OAI22_X1 U4975 ( .A1(n14847), .A2(n13213), .B1(n14815), .B2(n13210), .ZN(
        n4140) );
  AOI221_X1 U4976 ( .B1(n13165), .B2(n6022), .C1(n13162), .C2(n6054), .A(n4148), .ZN(n4141) );
  OAI22_X1 U4977 ( .A1(n15137), .A2(n13159), .B1(n15169), .B2(n13156), .ZN(
        n4148) );
  AOI221_X1 U4978 ( .B1(n13219), .B2(n606), .C1(n13216), .C2(n15724), .A(n4103), .ZN(n4096) );
  OAI22_X1 U4979 ( .A1(n14846), .A2(n13213), .B1(n14814), .B2(n13210), .ZN(
        n4103) );
  AOI221_X1 U4980 ( .B1(n13165), .B2(n6023), .C1(n13162), .C2(n6055), .A(n4111), .ZN(n4104) );
  OAI22_X1 U4981 ( .A1(n15136), .A2(n13159), .B1(n15168), .B2(n13156), .ZN(
        n4111) );
  AOI221_X1 U4982 ( .B1(n13219), .B2(n604), .C1(n13216), .C2(n15723), .A(n4066), .ZN(n4059) );
  OAI22_X1 U4983 ( .A1(n14845), .A2(n13213), .B1(n14813), .B2(n13210), .ZN(
        n4066) );
  AOI221_X1 U4984 ( .B1(n13165), .B2(n6024), .C1(n13162), .C2(n6056), .A(n4074), .ZN(n4067) );
  OAI22_X1 U4985 ( .A1(n15135), .A2(n13159), .B1(n15167), .B2(n13156), .ZN(
        n4074) );
  AOI221_X1 U4986 ( .B1(n13219), .B2(n602), .C1(n13216), .C2(n15722), .A(n4029), .ZN(n4022) );
  OAI22_X1 U4987 ( .A1(n14844), .A2(n13213), .B1(n14812), .B2(n13210), .ZN(
        n4029) );
  AOI221_X1 U4988 ( .B1(n13165), .B2(n6025), .C1(n13162), .C2(n6057), .A(n4037), .ZN(n4030) );
  OAI22_X1 U4989 ( .A1(n15134), .A2(n13159), .B1(n15166), .B2(n13156), .ZN(
        n4037) );
  AOI221_X1 U4990 ( .B1(n13219), .B2(n600), .C1(n13216), .C2(n15721), .A(n3992), .ZN(n3985) );
  OAI22_X1 U4991 ( .A1(n14843), .A2(n13213), .B1(n14811), .B2(n13210), .ZN(
        n3992) );
  AOI221_X1 U4992 ( .B1(n13165), .B2(n6026), .C1(n13162), .C2(n6058), .A(n4000), .ZN(n3993) );
  OAI22_X1 U4993 ( .A1(n15133), .A2(n13159), .B1(n15165), .B2(n13156), .ZN(
        n4000) );
  AOI221_X1 U4994 ( .B1(n13219), .B2(n598), .C1(n13216), .C2(n15720), .A(n3955), .ZN(n3948) );
  OAI22_X1 U4995 ( .A1(n14842), .A2(n13213), .B1(n14810), .B2(n13210), .ZN(
        n3955) );
  AOI221_X1 U4996 ( .B1(n13165), .B2(n6027), .C1(n13162), .C2(n6059), .A(n3963), .ZN(n3956) );
  OAI22_X1 U4997 ( .A1(n15132), .A2(n13159), .B1(n15164), .B2(n13156), .ZN(
        n3963) );
  AOI221_X1 U4998 ( .B1(n13219), .B2(n596), .C1(n13216), .C2(n15719), .A(n3918), .ZN(n3911) );
  OAI22_X1 U4999 ( .A1(n14841), .A2(n13213), .B1(n14809), .B2(n13210), .ZN(
        n3918) );
  AOI221_X1 U5000 ( .B1(n13165), .B2(n6028), .C1(n13162), .C2(n6060), .A(n3926), .ZN(n3919) );
  OAI22_X1 U5001 ( .A1(n15131), .A2(n13159), .B1(n15163), .B2(n13156), .ZN(
        n3926) );
  AOI221_X1 U5002 ( .B1(n13219), .B2(n594), .C1(n13216), .C2(n15718), .A(n3881), .ZN(n3874) );
  OAI22_X1 U5003 ( .A1(n14840), .A2(n13213), .B1(n14808), .B2(n13210), .ZN(
        n3881) );
  AOI221_X1 U5004 ( .B1(n13165), .B2(n6029), .C1(n13162), .C2(n6061), .A(n3889), .ZN(n3882) );
  OAI22_X1 U5005 ( .A1(n15130), .A2(n13159), .B1(n15162), .B2(n13156), .ZN(
        n3889) );
  OAI22_X1 U5006 ( .A1(n13829), .A2(n13407), .B1(n6942), .B2(n13402), .ZN(
        n7770) );
  OAI22_X1 U5007 ( .A1(n13835), .A2(n13407), .B1(n6943), .B2(n13402), .ZN(
        n7771) );
  OAI22_X1 U5008 ( .A1(n13841), .A2(n13407), .B1(n6944), .B2(n13402), .ZN(
        n7772) );
  OAI22_X1 U5009 ( .A1(n13847), .A2(n13407), .B1(n6945), .B2(n13402), .ZN(
        n7773) );
  OAI22_X1 U5010 ( .A1(n13853), .A2(n13407), .B1(n6946), .B2(n13402), .ZN(
        n7774) );
  OAI22_X1 U5011 ( .A1(n13859), .A2(n13407), .B1(n6947), .B2(n13402), .ZN(
        n7775) );
  OAI22_X1 U5012 ( .A1(n13865), .A2(n13407), .B1(n6948), .B2(n13402), .ZN(
        n7776) );
  OAI22_X1 U5013 ( .A1(n13871), .A2(n13407), .B1(n6949), .B2(n13402), .ZN(
        n7777) );
  OAI22_X1 U5014 ( .A1(n13877), .A2(n13406), .B1(n6950), .B2(n13402), .ZN(
        n7778) );
  OAI22_X1 U5015 ( .A1(n13883), .A2(n13406), .B1(n6951), .B2(n13402), .ZN(
        n7779) );
  OAI22_X1 U5016 ( .A1(n13889), .A2(n13406), .B1(n6952), .B2(n13402), .ZN(
        n7780) );
  OAI22_X1 U5017 ( .A1(n13895), .A2(n13406), .B1(n6953), .B2(n13402), .ZN(
        n7781) );
  OAI22_X1 U5018 ( .A1(n13901), .A2(n13406), .B1(n6954), .B2(n13403), .ZN(
        n7782) );
  OAI22_X1 U5019 ( .A1(n13907), .A2(n13406), .B1(n6955), .B2(n13403), .ZN(
        n7783) );
  OAI22_X1 U5020 ( .A1(n13913), .A2(n13406), .B1(n6956), .B2(n13403), .ZN(
        n7784) );
  OAI22_X1 U5021 ( .A1(n13919), .A2(n13406), .B1(n6957), .B2(n13403), .ZN(
        n7785) );
  OAI22_X1 U5022 ( .A1(n13925), .A2(n13406), .B1(n6958), .B2(n13403), .ZN(
        n7786) );
  OAI22_X1 U5023 ( .A1(n13931), .A2(n13406), .B1(n6959), .B2(n13403), .ZN(
        n7787) );
  OAI22_X1 U5024 ( .A1(n13937), .A2(n13406), .B1(n6960), .B2(n13403), .ZN(
        n7788) );
  OAI22_X1 U5025 ( .A1(n13943), .A2(n13406), .B1(n6961), .B2(n13403), .ZN(
        n7789) );
  OAI22_X1 U5026 ( .A1(n13949), .A2(n13405), .B1(n6962), .B2(n13403), .ZN(
        n7790) );
  OAI22_X1 U5027 ( .A1(n13955), .A2(n13405), .B1(n6963), .B2(n13403), .ZN(
        n7791) );
  OAI22_X1 U5028 ( .A1(n13961), .A2(n13405), .B1(n6964), .B2(n13403), .ZN(
        n7792) );
  OAI22_X1 U5029 ( .A1(n13967), .A2(n13405), .B1(n6965), .B2(n13403), .ZN(
        n7793) );
  OAI22_X1 U5030 ( .A1(n13973), .A2(n13405), .B1(n6966), .B2(n13404), .ZN(
        n7794) );
  OAI22_X1 U5031 ( .A1(n13979), .A2(n13405), .B1(n6967), .B2(n13404), .ZN(
        n7795) );
  OAI22_X1 U5032 ( .A1(n13985), .A2(n13405), .B1(n6968), .B2(n13404), .ZN(
        n7796) );
  OAI22_X1 U5033 ( .A1(n13991), .A2(n13405), .B1(n6969), .B2(n13404), .ZN(
        n7797) );
  OAI22_X1 U5034 ( .A1(n13997), .A2(n13405), .B1(n6970), .B2(n13404), .ZN(
        n7798) );
  OAI22_X1 U5035 ( .A1(n14003), .A2(n13405), .B1(n6971), .B2(n13404), .ZN(
        n7799) );
  OAI22_X1 U5036 ( .A1(n14009), .A2(n13405), .B1(n6972), .B2(n13404), .ZN(
        n7800) );
  OAI22_X1 U5037 ( .A1(n14018), .A2(n13405), .B1(n6973), .B2(n13404), .ZN(
        n7801) );
  OAI22_X1 U5038 ( .A1(n13829), .A2(n13413), .B1(n7160), .B2(n13408), .ZN(
        n7802) );
  OAI22_X1 U5039 ( .A1(n13835), .A2(n13413), .B1(n7161), .B2(n13408), .ZN(
        n7803) );
  OAI22_X1 U5040 ( .A1(n13841), .A2(n13413), .B1(n7162), .B2(n13408), .ZN(
        n7804) );
  OAI22_X1 U5041 ( .A1(n13847), .A2(n13413), .B1(n7163), .B2(n13408), .ZN(
        n7805) );
  OAI22_X1 U5042 ( .A1(n13853), .A2(n13413), .B1(n7164), .B2(n13408), .ZN(
        n7806) );
  OAI22_X1 U5043 ( .A1(n13859), .A2(n13413), .B1(n7165), .B2(n13408), .ZN(
        n7807) );
  OAI22_X1 U5044 ( .A1(n13865), .A2(n13413), .B1(n7166), .B2(n13408), .ZN(
        n7808) );
  OAI22_X1 U5045 ( .A1(n13871), .A2(n13413), .B1(n7167), .B2(n13408), .ZN(
        n7809) );
  OAI22_X1 U5046 ( .A1(n13877), .A2(n13412), .B1(n7168), .B2(n13408), .ZN(
        n7810) );
  OAI22_X1 U5047 ( .A1(n13883), .A2(n13412), .B1(n7169), .B2(n13408), .ZN(
        n7811) );
  OAI22_X1 U5048 ( .A1(n13889), .A2(n13412), .B1(n7170), .B2(n13408), .ZN(
        n7812) );
  OAI22_X1 U5049 ( .A1(n13895), .A2(n13412), .B1(n7171), .B2(n13408), .ZN(
        n7813) );
  OAI22_X1 U5050 ( .A1(n13901), .A2(n13412), .B1(n7172), .B2(n13409), .ZN(
        n7814) );
  OAI22_X1 U5051 ( .A1(n13907), .A2(n13412), .B1(n7173), .B2(n13409), .ZN(
        n7815) );
  OAI22_X1 U5052 ( .A1(n13913), .A2(n13412), .B1(n7174), .B2(n13409), .ZN(
        n7816) );
  OAI22_X1 U5053 ( .A1(n13919), .A2(n13412), .B1(n7175), .B2(n13409), .ZN(
        n7817) );
  OAI22_X1 U5054 ( .A1(n13925), .A2(n13412), .B1(n7176), .B2(n13409), .ZN(
        n7818) );
  OAI22_X1 U5055 ( .A1(n13931), .A2(n13412), .B1(n7177), .B2(n13409), .ZN(
        n7819) );
  OAI22_X1 U5056 ( .A1(n13937), .A2(n13412), .B1(n7178), .B2(n13409), .ZN(
        n7820) );
  OAI22_X1 U5057 ( .A1(n13943), .A2(n13412), .B1(n7179), .B2(n13409), .ZN(
        n7821) );
  OAI22_X1 U5058 ( .A1(n13949), .A2(n13411), .B1(n7180), .B2(n13409), .ZN(
        n7822) );
  OAI22_X1 U5059 ( .A1(n13955), .A2(n13411), .B1(n7181), .B2(n13409), .ZN(
        n7823) );
  OAI22_X1 U5060 ( .A1(n13961), .A2(n13411), .B1(n7182), .B2(n13409), .ZN(
        n7824) );
  OAI22_X1 U5061 ( .A1(n13967), .A2(n13411), .B1(n7183), .B2(n13409), .ZN(
        n7825) );
  OAI22_X1 U5062 ( .A1(n13973), .A2(n13411), .B1(n7184), .B2(n13410), .ZN(
        n7826) );
  OAI22_X1 U5063 ( .A1(n13979), .A2(n13411), .B1(n7185), .B2(n13410), .ZN(
        n7827) );
  OAI22_X1 U5064 ( .A1(n13985), .A2(n13411), .B1(n7186), .B2(n13410), .ZN(
        n7828) );
  OAI22_X1 U5065 ( .A1(n13991), .A2(n13411), .B1(n7187), .B2(n13410), .ZN(
        n7829) );
  OAI22_X1 U5066 ( .A1(n13997), .A2(n13411), .B1(n7188), .B2(n13410), .ZN(
        n7830) );
  OAI22_X1 U5067 ( .A1(n14003), .A2(n13411), .B1(n7189), .B2(n13410), .ZN(
        n7831) );
  OAI22_X1 U5068 ( .A1(n14009), .A2(n13411), .B1(n7190), .B2(n13410), .ZN(
        n7832) );
  OAI22_X1 U5069 ( .A1(n14018), .A2(n13411), .B1(n7191), .B2(n13410), .ZN(
        n7833) );
  OAI22_X1 U5070 ( .A1(n13835), .A2(n13437), .B1(n7193), .B2(n13432), .ZN(
        n7931) );
  OAI22_X1 U5071 ( .A1(n13841), .A2(n13437), .B1(n7194), .B2(n13432), .ZN(
        n7932) );
  OAI22_X1 U5072 ( .A1(n13847), .A2(n13437), .B1(n7195), .B2(n13432), .ZN(
        n7933) );
  OAI22_X1 U5073 ( .A1(n13853), .A2(n13437), .B1(n7196), .B2(n13432), .ZN(
        n7934) );
  OAI22_X1 U5074 ( .A1(n13859), .A2(n13437), .B1(n7197), .B2(n13432), .ZN(
        n7935) );
  OAI22_X1 U5075 ( .A1(n13865), .A2(n13437), .B1(n7198), .B2(n13432), .ZN(
        n7936) );
  OAI22_X1 U5076 ( .A1(n13871), .A2(n13437), .B1(n7199), .B2(n13432), .ZN(
        n7937) );
  OAI22_X1 U5077 ( .A1(n13877), .A2(n13436), .B1(n7200), .B2(n13432), .ZN(
        n7938) );
  OAI22_X1 U5078 ( .A1(n13883), .A2(n13436), .B1(n7201), .B2(n13432), .ZN(
        n7939) );
  OAI22_X1 U5079 ( .A1(n13889), .A2(n13436), .B1(n7202), .B2(n13432), .ZN(
        n7940) );
  OAI22_X1 U5080 ( .A1(n13895), .A2(n13436), .B1(n7203), .B2(n13432), .ZN(
        n7941) );
  OAI22_X1 U5081 ( .A1(n13901), .A2(n13436), .B1(n7204), .B2(n13433), .ZN(
        n7942) );
  OAI22_X1 U5082 ( .A1(n13907), .A2(n13436), .B1(n7205), .B2(n13433), .ZN(
        n7943) );
  OAI22_X1 U5083 ( .A1(n13913), .A2(n13436), .B1(n7206), .B2(n13433), .ZN(
        n7944) );
  OAI22_X1 U5084 ( .A1(n13919), .A2(n13436), .B1(n7207), .B2(n13433), .ZN(
        n7945) );
  OAI22_X1 U5085 ( .A1(n13925), .A2(n13436), .B1(n7208), .B2(n13433), .ZN(
        n7946) );
  OAI22_X1 U5086 ( .A1(n13931), .A2(n13436), .B1(n7209), .B2(n13433), .ZN(
        n7947) );
  OAI22_X1 U5087 ( .A1(n13937), .A2(n13436), .B1(n7210), .B2(n13433), .ZN(
        n7948) );
  OAI22_X1 U5088 ( .A1(n13943), .A2(n13436), .B1(n7211), .B2(n13433), .ZN(
        n7949) );
  OAI22_X1 U5089 ( .A1(n13949), .A2(n13435), .B1(n7212), .B2(n13433), .ZN(
        n7950) );
  OAI22_X1 U5090 ( .A1(n13955), .A2(n13435), .B1(n7213), .B2(n13433), .ZN(
        n7951) );
  OAI22_X1 U5091 ( .A1(n13961), .A2(n13435), .B1(n7214), .B2(n13433), .ZN(
        n7952) );
  OAI22_X1 U5092 ( .A1(n13967), .A2(n13435), .B1(n7215), .B2(n13433), .ZN(
        n7953) );
  OAI22_X1 U5093 ( .A1(n13973), .A2(n13435), .B1(n7216), .B2(n13434), .ZN(
        n7954) );
  OAI22_X1 U5094 ( .A1(n13979), .A2(n13435), .B1(n7217), .B2(n13434), .ZN(
        n7955) );
  OAI22_X1 U5095 ( .A1(n13985), .A2(n13435), .B1(n7218), .B2(n13434), .ZN(
        n7956) );
  OAI22_X1 U5096 ( .A1(n13991), .A2(n13435), .B1(n7219), .B2(n13434), .ZN(
        n7957) );
  OAI22_X1 U5097 ( .A1(n13997), .A2(n13435), .B1(n7220), .B2(n13434), .ZN(
        n7958) );
  OAI22_X1 U5098 ( .A1(n14003), .A2(n13435), .B1(n7221), .B2(n13434), .ZN(
        n7959) );
  OAI22_X1 U5099 ( .A1(n14009), .A2(n13435), .B1(n7222), .B2(n13434), .ZN(
        n7960) );
  OAI22_X1 U5100 ( .A1(n14018), .A2(n13435), .B1(n7223), .B2(n13434), .ZN(
        n7961) );
  OAI22_X1 U5101 ( .A1(n14016), .A2(n13579), .B1(n13578), .B2(n12709), .ZN(
        n8729) );
  OAI22_X1 U5102 ( .A1(n14005), .A2(n13687), .B1(n13686), .B2(n14460), .ZN(
        n9304) );
  OAI22_X1 U5103 ( .A1(n14014), .A2(n13687), .B1(n13686), .B2(n14459), .ZN(
        n9305) );
  OAI22_X1 U5104 ( .A1(n13972), .A2(n13471), .B1(n13470), .B2(n12710), .ZN(
        n8146) );
  OAI22_X1 U5105 ( .A1(n13978), .A2(n13471), .B1(n13470), .B2(n12711), .ZN(
        n8147) );
  OAI22_X1 U5106 ( .A1(n13984), .A2(n13471), .B1(n13470), .B2(n12712), .ZN(
        n8148) );
  OAI22_X1 U5107 ( .A1(n13990), .A2(n13471), .B1(n13470), .B2(n12713), .ZN(
        n8149) );
  OAI22_X1 U5108 ( .A1(n13996), .A2(n13471), .B1(n13470), .B2(n12714), .ZN(
        n8150) );
  OAI22_X1 U5109 ( .A1(n14002), .A2(n13471), .B1(n13470), .B2(n12715), .ZN(
        n8151) );
  OAI22_X1 U5110 ( .A1(n14008), .A2(n13471), .B1(n13470), .B2(n12716), .ZN(
        n8152) );
  OAI22_X1 U5111 ( .A1(n14017), .A2(n13471), .B1(n13470), .B2(n12717), .ZN(
        n8153) );
  OAI22_X1 U5112 ( .A1(n13972), .A2(n13477), .B1(n13476), .B2(n12718), .ZN(
        n8178) );
  OAI22_X1 U5113 ( .A1(n13978), .A2(n13477), .B1(n13476), .B2(n12719), .ZN(
        n8179) );
  OAI22_X1 U5114 ( .A1(n13984), .A2(n13477), .B1(n13476), .B2(n12720), .ZN(
        n8180) );
  OAI22_X1 U5115 ( .A1(n13990), .A2(n13477), .B1(n13476), .B2(n12721), .ZN(
        n8181) );
  OAI22_X1 U5116 ( .A1(n13996), .A2(n13477), .B1(n13476), .B2(n12722), .ZN(
        n8182) );
  OAI22_X1 U5117 ( .A1(n14002), .A2(n13477), .B1(n13476), .B2(n12723), .ZN(
        n8183) );
  OAI22_X1 U5118 ( .A1(n14008), .A2(n13477), .B1(n13476), .B2(n12724), .ZN(
        n8184) );
  OAI22_X1 U5119 ( .A1(n14017), .A2(n13477), .B1(n13476), .B2(n12725), .ZN(
        n8185) );
  OAI22_X1 U5120 ( .A1(n14019), .A2(n13968), .B1(n6930), .B2(n14012), .ZN(
        n9970) );
  OAI22_X1 U5121 ( .A1(n14019), .A2(n13974), .B1(n6931), .B2(n14012), .ZN(
        n9971) );
  OAI22_X1 U5122 ( .A1(n14019), .A2(n13980), .B1(n6932), .B2(n14012), .ZN(
        n9972) );
  OAI22_X1 U5123 ( .A1(n14019), .A2(n13986), .B1(n6933), .B2(n14012), .ZN(
        n9973) );
  OAI22_X1 U5124 ( .A1(n14019), .A2(n13992), .B1(n6934), .B2(n14012), .ZN(
        n9974) );
  OAI22_X1 U5125 ( .A1(n14019), .A2(n13998), .B1(n6935), .B2(n14012), .ZN(
        n9975) );
  OAI22_X1 U5126 ( .A1(n14019), .A2(n14004), .B1(n6936), .B2(n14012), .ZN(
        n9976) );
  OAI22_X1 U5127 ( .A1(n14019), .A2(n14013), .B1(n6937), .B2(n14012), .ZN(
        n9977) );
  OAI22_X1 U5128 ( .A1(n13968), .A2(n13795), .B1(n5627), .B2(n13794), .ZN(
        n9874) );
  OAI22_X1 U5129 ( .A1(n13974), .A2(n13795), .B1(n5637), .B2(n13794), .ZN(
        n9875) );
  OAI22_X1 U5130 ( .A1(n13980), .A2(n13795), .B1(n5647), .B2(n13794), .ZN(
        n9876) );
  OAI22_X1 U5131 ( .A1(n13986), .A2(n13795), .B1(n5657), .B2(n13794), .ZN(
        n9877) );
  OAI22_X1 U5132 ( .A1(n13992), .A2(n13795), .B1(n5667), .B2(n13794), .ZN(
        n9878) );
  OAI22_X1 U5133 ( .A1(n13998), .A2(n13795), .B1(n5677), .B2(n13794), .ZN(
        n9879) );
  OAI22_X1 U5134 ( .A1(n14004), .A2(n13795), .B1(n5687), .B2(n13794), .ZN(
        n9880) );
  OAI22_X1 U5135 ( .A1(n14013), .A2(n13795), .B1(n5697), .B2(n13794), .ZN(
        n9881) );
  OAI22_X1 U5136 ( .A1(n13969), .A2(n13741), .B1(n5625), .B2(n13740), .ZN(
        n9586) );
  OAI22_X1 U5137 ( .A1(n13975), .A2(n13741), .B1(n5635), .B2(n13740), .ZN(
        n9587) );
  OAI22_X1 U5138 ( .A1(n13981), .A2(n13741), .B1(n5645), .B2(n13740), .ZN(
        n9588) );
  OAI22_X1 U5139 ( .A1(n13987), .A2(n13741), .B1(n5655), .B2(n13740), .ZN(
        n9589) );
  OAI22_X1 U5140 ( .A1(n13993), .A2(n13741), .B1(n5665), .B2(n13740), .ZN(
        n9590) );
  OAI22_X1 U5141 ( .A1(n13999), .A2(n13741), .B1(n5675), .B2(n13740), .ZN(
        n9591) );
  OAI22_X1 U5142 ( .A1(n14005), .A2(n13741), .B1(n5685), .B2(n13740), .ZN(
        n9592) );
  OAI22_X1 U5143 ( .A1(n14014), .A2(n13741), .B1(n5695), .B2(n13740), .ZN(
        n9593) );
  OAI22_X1 U5144 ( .A1(n13969), .A2(n13693), .B1(n5796), .B2(n13692), .ZN(
        n9330) );
  OAI22_X1 U5145 ( .A1(n13975), .A2(n13693), .B1(n5800), .B2(n13692), .ZN(
        n9331) );
  OAI22_X1 U5146 ( .A1(n13981), .A2(n13693), .B1(n5804), .B2(n13692), .ZN(
        n9332) );
  OAI22_X1 U5147 ( .A1(n13987), .A2(n13693), .B1(n5808), .B2(n13692), .ZN(
        n9333) );
  OAI22_X1 U5148 ( .A1(n13993), .A2(n13693), .B1(n5812), .B2(n13692), .ZN(
        n9334) );
  OAI22_X1 U5149 ( .A1(n13999), .A2(n13693), .B1(n5816), .B2(n13692), .ZN(
        n9335) );
  OAI22_X1 U5150 ( .A1(n14005), .A2(n13693), .B1(n5820), .B2(n13692), .ZN(
        n9336) );
  OAI22_X1 U5151 ( .A1(n14014), .A2(n13693), .B1(n5824), .B2(n13692), .ZN(
        n9337) );
  OAI22_X1 U5152 ( .A1(n13970), .A2(n13639), .B1(n5622), .B2(n13638), .ZN(
        n9042) );
  OAI22_X1 U5153 ( .A1(n13976), .A2(n13639), .B1(n5632), .B2(n13638), .ZN(
        n9043) );
  OAI22_X1 U5154 ( .A1(n13982), .A2(n13639), .B1(n5642), .B2(n13638), .ZN(
        n9044) );
  OAI22_X1 U5155 ( .A1(n13988), .A2(n13639), .B1(n5652), .B2(n13638), .ZN(
        n9045) );
  OAI22_X1 U5156 ( .A1(n13994), .A2(n13639), .B1(n5662), .B2(n13638), .ZN(
        n9046) );
  OAI22_X1 U5157 ( .A1(n14000), .A2(n13639), .B1(n5672), .B2(n13638), .ZN(
        n9047) );
  OAI22_X1 U5159 ( .A1(n14006), .A2(n13639), .B1(n5682), .B2(n13638), .ZN(
        n9048) );
  OAI22_X1 U5160 ( .A1(n14015), .A2(n13639), .B1(n5692), .B2(n13638), .ZN(
        n9049) );
  OAI22_X1 U5161 ( .A1(n13971), .A2(n13519), .B1(n976), .B2(n13518), .ZN(n8402) );
  OAI22_X1 U5162 ( .A1(n13977), .A2(n13519), .B1(n975), .B2(n13518), .ZN(n8403) );
  OAI22_X1 U5163 ( .A1(n13983), .A2(n13519), .B1(n974), .B2(n13518), .ZN(n8404) );
  OAI22_X1 U5164 ( .A1(n13989), .A2(n13519), .B1(n973), .B2(n13518), .ZN(n8405) );
  OAI22_X1 U5165 ( .A1(n13995), .A2(n13519), .B1(n972), .B2(n13518), .ZN(n8406) );
  OAI22_X1 U5166 ( .A1(n14001), .A2(n13519), .B1(n971), .B2(n13518), .ZN(n8407) );
  OAI22_X1 U5167 ( .A1(n14007), .A2(n13519), .B1(n970), .B2(n13518), .ZN(n8408) );
  OAI22_X1 U5168 ( .A1(n14016), .A2(n13519), .B1(n969), .B2(n13518), .ZN(n8409) );
  OAI22_X1 U5169 ( .A1(n13971), .A2(n13543), .B1(n640), .B2(n13542), .ZN(n8530) );
  OAI22_X1 U5170 ( .A1(n13977), .A2(n13543), .B1(n637), .B2(n13542), .ZN(n8531) );
  OAI22_X1 U5171 ( .A1(n13983), .A2(n13543), .B1(n634), .B2(n13542), .ZN(n8532) );
  OAI22_X1 U5172 ( .A1(n13989), .A2(n13543), .B1(n631), .B2(n13542), .ZN(n8533) );
  OAI22_X1 U5173 ( .A1(n13995), .A2(n13543), .B1(n628), .B2(n13542), .ZN(n8534) );
  OAI22_X1 U5174 ( .A1(n14001), .A2(n13543), .B1(n625), .B2(n13542), .ZN(n8535) );
  OAI22_X1 U5175 ( .A1(n14007), .A2(n13543), .B1(n622), .B2(n13542), .ZN(n8536) );
  OAI22_X1 U5176 ( .A1(n13968), .A2(n13789), .B1(n816), .B2(n13788), .ZN(n9842) );
  OAI22_X1 U5177 ( .A1(n13974), .A2(n13789), .B1(n815), .B2(n13788), .ZN(n9843) );
  OAI22_X1 U5178 ( .A1(n13980), .A2(n13789), .B1(n814), .B2(n13788), .ZN(n9844) );
  OAI22_X1 U5179 ( .A1(n13986), .A2(n13789), .B1(n813), .B2(n13788), .ZN(n9845) );
  OAI22_X1 U5180 ( .A1(n13992), .A2(n13789), .B1(n812), .B2(n13788), .ZN(n9846) );
  OAI22_X1 U5181 ( .A1(n13998), .A2(n13789), .B1(n811), .B2(n13788), .ZN(n9847) );
  OAI22_X1 U5182 ( .A1(n14004), .A2(n13789), .B1(n810), .B2(n13788), .ZN(n9848) );
  OAI22_X1 U5183 ( .A1(n14013), .A2(n13789), .B1(n809), .B2(n13788), .ZN(n9849) );
  OAI22_X1 U5184 ( .A1(n13969), .A2(n13735), .B1(n848), .B2(n13734), .ZN(n9554) );
  OAI22_X1 U5185 ( .A1(n13975), .A2(n13735), .B1(n847), .B2(n13734), .ZN(n9555) );
  OAI22_X1 U5186 ( .A1(n13981), .A2(n13735), .B1(n846), .B2(n13734), .ZN(n9556) );
  OAI22_X1 U5187 ( .A1(n13987), .A2(n13735), .B1(n845), .B2(n13734), .ZN(n9557) );
  OAI22_X1 U5188 ( .A1(n13993), .A2(n13735), .B1(n844), .B2(n13734), .ZN(n9558) );
  OAI22_X1 U5189 ( .A1(n13999), .A2(n13735), .B1(n843), .B2(n13734), .ZN(n9559) );
  OAI22_X1 U5190 ( .A1(n14005), .A2(n13735), .B1(n842), .B2(n13734), .ZN(n9560) );
  OAI22_X1 U5191 ( .A1(n14014), .A2(n13735), .B1(n841), .B2(n13734), .ZN(n9561) );
  OAI22_X1 U5192 ( .A1(n13969), .A2(n13681), .B1(n880), .B2(n13680), .ZN(n9266) );
  OAI22_X1 U5193 ( .A1(n13975), .A2(n13681), .B1(n879), .B2(n13680), .ZN(n9267) );
  OAI22_X1 U5194 ( .A1(n13981), .A2(n13681), .B1(n878), .B2(n13680), .ZN(n9268) );
  OAI22_X1 U5195 ( .A1(n13987), .A2(n13681), .B1(n877), .B2(n13680), .ZN(n9269) );
  OAI22_X1 U5196 ( .A1(n13993), .A2(n13681), .B1(n876), .B2(n13680), .ZN(n9270) );
  OAI22_X1 U5197 ( .A1(n13999), .A2(n13681), .B1(n875), .B2(n13680), .ZN(n9271) );
  OAI22_X1 U5198 ( .A1(n14005), .A2(n13681), .B1(n874), .B2(n13680), .ZN(n9272) );
  OAI22_X1 U5199 ( .A1(n14014), .A2(n13681), .B1(n873), .B2(n13680), .ZN(n9273) );
  OAI22_X1 U5200 ( .A1(n13970), .A2(n13633), .B1(n5623), .B2(n13632), .ZN(
        n9010) );
  OAI22_X1 U5201 ( .A1(n13976), .A2(n13633), .B1(n5633), .B2(n13632), .ZN(
        n9011) );
  OAI22_X1 U5202 ( .A1(n13982), .A2(n13633), .B1(n5643), .B2(n13632), .ZN(
        n9012) );
  OAI22_X1 U5203 ( .A1(n13988), .A2(n13633), .B1(n5653), .B2(n13632), .ZN(
        n9013) );
  OAI22_X1 U5204 ( .A1(n13994), .A2(n13633), .B1(n5663), .B2(n13632), .ZN(
        n9014) );
  OAI22_X1 U5205 ( .A1(n14000), .A2(n13633), .B1(n5673), .B2(n13632), .ZN(
        n9015) );
  OAI22_X1 U5206 ( .A1(n14006), .A2(n13633), .B1(n5683), .B2(n13632), .ZN(
        n9016) );
  OAI22_X1 U5207 ( .A1(n14015), .A2(n13633), .B1(n5693), .B2(n13632), .ZN(
        n9017) );
  OAI22_X1 U5208 ( .A1(n13970), .A2(n13627), .B1(n912), .B2(n13626), .ZN(n8978) );
  OAI22_X1 U5209 ( .A1(n13976), .A2(n13627), .B1(n911), .B2(n13626), .ZN(n8979) );
  OAI22_X1 U5210 ( .A1(n13982), .A2(n13627), .B1(n910), .B2(n13626), .ZN(n8980) );
  OAI22_X1 U5211 ( .A1(n13988), .A2(n13627), .B1(n909), .B2(n13626), .ZN(n8981) );
  OAI22_X1 U5212 ( .A1(n13994), .A2(n13627), .B1(n908), .B2(n13626), .ZN(n8982) );
  OAI22_X1 U5213 ( .A1(n14000), .A2(n13627), .B1(n907), .B2(n13626), .ZN(n8983) );
  OAI22_X1 U5214 ( .A1(n14006), .A2(n13627), .B1(n906), .B2(n13626), .ZN(n8984) );
  OAI22_X1 U5215 ( .A1(n14015), .A2(n13627), .B1(n905), .B2(n13626), .ZN(n8985) );
  OAI22_X1 U5216 ( .A1(n13971), .A2(n13573), .B1(n944), .B2(n13572), .ZN(n8690) );
  OAI22_X1 U5217 ( .A1(n13977), .A2(n13573), .B1(n943), .B2(n13572), .ZN(n8691) );
  OAI22_X1 U5218 ( .A1(n13983), .A2(n13573), .B1(n942), .B2(n13572), .ZN(n8692) );
  OAI22_X1 U5219 ( .A1(n13989), .A2(n13573), .B1(n941), .B2(n13572), .ZN(n8693) );
  OAI22_X1 U5220 ( .A1(n13995), .A2(n13573), .B1(n940), .B2(n13572), .ZN(n8694) );
  OAI22_X1 U5221 ( .A1(n14001), .A2(n13573), .B1(n939), .B2(n13572), .ZN(n8695) );
  OAI22_X1 U5222 ( .A1(n14007), .A2(n13573), .B1(n938), .B2(n13572), .ZN(n8696) );
  OAI22_X1 U5223 ( .A1(n14016), .A2(n13573), .B1(n937), .B2(n13572), .ZN(n8697) );
  OAI22_X1 U5224 ( .A1(n13972), .A2(n13465), .B1(n7248), .B2(n13464), .ZN(
        n8114) );
  OAI22_X1 U5225 ( .A1(n13978), .A2(n13465), .B1(n7249), .B2(n13464), .ZN(
        n8115) );
  OAI22_X1 U5226 ( .A1(n13984), .A2(n13465), .B1(n7250), .B2(n13464), .ZN(
        n8116) );
  OAI22_X1 U5227 ( .A1(n13990), .A2(n13465), .B1(n7251), .B2(n13464), .ZN(
        n8117) );
  OAI22_X1 U5228 ( .A1(n13996), .A2(n13465), .B1(n7252), .B2(n13464), .ZN(
        n8118) );
  OAI22_X1 U5229 ( .A1(n14002), .A2(n13465), .B1(n7253), .B2(n13464), .ZN(
        n8119) );
  OAI22_X1 U5230 ( .A1(n14008), .A2(n13465), .B1(n7254), .B2(n13464), .ZN(
        n8120) );
  OAI22_X1 U5231 ( .A1(n14017), .A2(n13465), .B1(n7255), .B2(n13464), .ZN(
        n8121) );
  OAI22_X1 U5232 ( .A1(n13972), .A2(n13513), .B1(n6974), .B2(n13512), .ZN(
        n8370) );
  OAI22_X1 U5233 ( .A1(n13978), .A2(n13513), .B1(n6975), .B2(n13512), .ZN(
        n8371) );
  OAI22_X1 U5234 ( .A1(n13984), .A2(n13513), .B1(n6976), .B2(n13512), .ZN(
        n8372) );
  OAI22_X1 U5235 ( .A1(n13990), .A2(n13513), .B1(n6977), .B2(n13512), .ZN(
        n8373) );
  OAI22_X1 U5236 ( .A1(n13996), .A2(n13513), .B1(n6978), .B2(n13512), .ZN(
        n8374) );
  OAI22_X1 U5237 ( .A1(n14002), .A2(n13513), .B1(n6979), .B2(n13512), .ZN(
        n8375) );
  OAI22_X1 U5238 ( .A1(n14008), .A2(n13513), .B1(n6980), .B2(n13512), .ZN(
        n8376) );
  OAI22_X1 U5239 ( .A1(n14017), .A2(n13513), .B1(n6981), .B2(n13512), .ZN(
        n8377) );
  OAI22_X1 U5240 ( .A1(n14016), .A2(n13543), .B1(n7257), .B2(n13542), .ZN(
        n8537) );
  OAI22_X1 U5241 ( .A1(n13970), .A2(n13621), .B1(n6982), .B2(n13620), .ZN(
        n8946) );
  OAI22_X1 U5242 ( .A1(n13976), .A2(n13621), .B1(n6983), .B2(n13620), .ZN(
        n8947) );
  OAI22_X1 U5243 ( .A1(n13982), .A2(n13621), .B1(n6984), .B2(n13620), .ZN(
        n8948) );
  OAI22_X1 U5244 ( .A1(n13988), .A2(n13621), .B1(n6985), .B2(n13620), .ZN(
        n8949) );
  OAI22_X1 U5245 ( .A1(n13994), .A2(n13621), .B1(n6986), .B2(n13620), .ZN(
        n8950) );
  OAI22_X1 U5246 ( .A1(n14000), .A2(n13621), .B1(n6987), .B2(n13620), .ZN(
        n8951) );
  OAI22_X1 U5247 ( .A1(n14006), .A2(n13621), .B1(n6988), .B2(n13620), .ZN(
        n8952) );
  OAI22_X1 U5248 ( .A1(n14015), .A2(n13621), .B1(n6989), .B2(n13620), .ZN(
        n8953) );
  OAI22_X1 U5249 ( .A1(n13969), .A2(n13675), .B1(n6990), .B2(n13674), .ZN(
        n9234) );
  OAI22_X1 U5250 ( .A1(n13975), .A2(n13675), .B1(n6991), .B2(n13674), .ZN(
        n9235) );
  OAI22_X1 U5251 ( .A1(n13981), .A2(n13675), .B1(n6992), .B2(n13674), .ZN(
        n9236) );
  OAI22_X1 U5253 ( .A1(n13987), .A2(n13675), .B1(n6993), .B2(n13674), .ZN(
        n9237) );
  OAI22_X1 U5254 ( .A1(n13993), .A2(n13675), .B1(n6994), .B2(n13674), .ZN(
        n9238) );
  OAI22_X1 U5255 ( .A1(n13999), .A2(n13675), .B1(n6995), .B2(n13674), .ZN(
        n9239) );
  OAI22_X1 U5256 ( .A1(n14005), .A2(n13675), .B1(n6996), .B2(n13674), .ZN(
        n9240) );
  OAI22_X1 U5257 ( .A1(n14014), .A2(n13675), .B1(n6997), .B2(n13674), .ZN(
        n9241) );
  OAI22_X1 U5258 ( .A1(n13969), .A2(n13729), .B1(n7006), .B2(n13728), .ZN(
        n9522) );
  OAI22_X1 U5259 ( .A1(n13975), .A2(n13729), .B1(n7007), .B2(n13728), .ZN(
        n9523) );
  OAI22_X1 U5260 ( .A1(n13981), .A2(n13729), .B1(n7008), .B2(n13728), .ZN(
        n9524) );
  OAI22_X1 U5261 ( .A1(n13987), .A2(n13729), .B1(n7009), .B2(n13728), .ZN(
        n9525) );
  OAI22_X1 U5262 ( .A1(n13993), .A2(n13729), .B1(n7010), .B2(n13728), .ZN(
        n9526) );
  OAI22_X1 U5263 ( .A1(n13999), .A2(n13729), .B1(n7011), .B2(n13728), .ZN(
        n9527) );
  OAI22_X1 U5264 ( .A1(n14005), .A2(n13729), .B1(n7012), .B2(n13728), .ZN(
        n9528) );
  OAI22_X1 U5265 ( .A1(n14014), .A2(n13729), .B1(n7013), .B2(n13728), .ZN(
        n9529) );
  OAI22_X1 U5266 ( .A1(n13969), .A2(n13753), .B1(n6786), .B2(n13752), .ZN(
        n9650) );
  OAI22_X1 U5267 ( .A1(n13975), .A2(n13753), .B1(n6787), .B2(n13752), .ZN(
        n9651) );
  OAI22_X1 U5268 ( .A1(n13981), .A2(n13753), .B1(n6788), .B2(n13752), .ZN(
        n9652) );
  OAI22_X1 U5269 ( .A1(n13987), .A2(n13753), .B1(n6789), .B2(n13752), .ZN(
        n9653) );
  OAI22_X1 U5270 ( .A1(n13993), .A2(n13753), .B1(n6790), .B2(n13752), .ZN(
        n9654) );
  OAI22_X1 U5271 ( .A1(n13999), .A2(n13753), .B1(n6791), .B2(n13752), .ZN(
        n9655) );
  OAI22_X1 U5272 ( .A1(n14005), .A2(n13753), .B1(n6792), .B2(n13752), .ZN(
        n9656) );
  OAI22_X1 U5273 ( .A1(n14014), .A2(n13753), .B1(n6793), .B2(n13752), .ZN(
        n9657) );
  OAI22_X1 U5274 ( .A1(n13968), .A2(n13759), .B1(n6914), .B2(n13758), .ZN(
        n9682) );
  OAI22_X1 U5275 ( .A1(n13974), .A2(n13759), .B1(n6915), .B2(n13758), .ZN(
        n9683) );
  OAI22_X1 U5276 ( .A1(n13980), .A2(n13759), .B1(n6916), .B2(n13758), .ZN(
        n9684) );
  OAI22_X1 U5277 ( .A1(n13986), .A2(n13759), .B1(n6917), .B2(n13758), .ZN(
        n9685) );
  OAI22_X1 U5278 ( .A1(n13992), .A2(n13759), .B1(n6918), .B2(n13758), .ZN(
        n9686) );
  OAI22_X1 U5279 ( .A1(n13998), .A2(n13759), .B1(n6919), .B2(n13758), .ZN(
        n9687) );
  OAI22_X1 U5280 ( .A1(n14004), .A2(n13759), .B1(n6920), .B2(n13758), .ZN(
        n9688) );
  OAI22_X1 U5281 ( .A1(n14013), .A2(n13759), .B1(n6921), .B2(n13758), .ZN(
        n9689) );
  OAI22_X1 U5282 ( .A1(n13968), .A2(n13783), .B1(n7014), .B2(n13782), .ZN(
        n9810) );
  OAI22_X1 U5283 ( .A1(n13974), .A2(n13783), .B1(n7015), .B2(n13782), .ZN(
        n9811) );
  OAI22_X1 U5284 ( .A1(n13980), .A2(n13783), .B1(n7016), .B2(n13782), .ZN(
        n9812) );
  OAI22_X1 U5285 ( .A1(n13986), .A2(n13783), .B1(n7017), .B2(n13782), .ZN(
        n9813) );
  OAI22_X1 U5286 ( .A1(n13992), .A2(n13783), .B1(n7018), .B2(n13782), .ZN(
        n9814) );
  OAI22_X1 U5287 ( .A1(n13998), .A2(n13783), .B1(n7019), .B2(n13782), .ZN(
        n9815) );
  OAI22_X1 U5288 ( .A1(n14004), .A2(n13783), .B1(n7020), .B2(n13782), .ZN(
        n9816) );
  OAI22_X1 U5289 ( .A1(n14013), .A2(n13783), .B1(n7021), .B2(n13782), .ZN(
        n9817) );
  OAI22_X1 U5290 ( .A1(n13968), .A2(n13807), .B1(n6802), .B2(n13806), .ZN(
        n9938) );
  OAI22_X1 U5291 ( .A1(n13974), .A2(n13807), .B1(n6803), .B2(n13806), .ZN(
        n9939) );
  OAI22_X1 U5292 ( .A1(n13980), .A2(n13807), .B1(n6804), .B2(n13806), .ZN(
        n9940) );
  OAI22_X1 U5293 ( .A1(n13986), .A2(n13807), .B1(n6805), .B2(n13806), .ZN(
        n9941) );
  OAI22_X1 U5294 ( .A1(n13992), .A2(n13807), .B1(n6806), .B2(n13806), .ZN(
        n9942) );
  OAI22_X1 U5295 ( .A1(n13998), .A2(n13807), .B1(n6807), .B2(n13806), .ZN(
        n9943) );
  OAI22_X1 U5296 ( .A1(n14004), .A2(n13807), .B1(n6808), .B2(n13806), .ZN(
        n9944) );
  OAI22_X1 U5297 ( .A1(n14013), .A2(n13807), .B1(n6809), .B2(n13806), .ZN(
        n9945) );
  OAI22_X1 U5298 ( .A1(n13971), .A2(n13579), .B1(n5795), .B2(n13578), .ZN(
        n8722) );
  OAI22_X1 U5299 ( .A1(n13977), .A2(n13579), .B1(n5799), .B2(n13578), .ZN(
        n8723) );
  OAI22_X1 U5300 ( .A1(n13983), .A2(n13579), .B1(n5803), .B2(n13578), .ZN(
        n8724) );
  OAI22_X1 U5301 ( .A1(n13989), .A2(n13579), .B1(n5807), .B2(n13578), .ZN(
        n8725) );
  OAI22_X1 U5302 ( .A1(n13995), .A2(n13579), .B1(n5811), .B2(n13578), .ZN(
        n8726) );
  OAI22_X1 U5303 ( .A1(n14001), .A2(n13579), .B1(n5815), .B2(n13578), .ZN(
        n8727) );
  OAI22_X1 U5304 ( .A1(n14007), .A2(n13579), .B1(n5819), .B2(n13578), .ZN(
        n8728) );
  OAI22_X1 U5305 ( .A1(n13969), .A2(n13687), .B1(n5797), .B2(n13686), .ZN(
        n9298) );
  OAI22_X1 U5306 ( .A1(n13975), .A2(n13687), .B1(n5801), .B2(n13686), .ZN(
        n9299) );
  OAI22_X1 U5307 ( .A1(n13981), .A2(n13687), .B1(n5805), .B2(n13686), .ZN(
        n9300) );
  OAI22_X1 U5308 ( .A1(n13987), .A2(n13687), .B1(n5809), .B2(n13686), .ZN(
        n9301) );
  OAI22_X1 U5309 ( .A1(n13993), .A2(n13687), .B1(n5813), .B2(n13686), .ZN(
        n9302) );
  OAI22_X1 U5310 ( .A1(n13999), .A2(n13687), .B1(n5817), .B2(n13686), .ZN(
        n9303) );
  OAI22_X1 U5311 ( .A1(n14020), .A2(n13896), .B1(n675), .B2(n14011), .ZN(n9958) );
  OAI22_X1 U5312 ( .A1(n14020), .A2(n13902), .B1(n672), .B2(n14011), .ZN(n9959) );
  OAI22_X1 U5313 ( .A1(n14020), .A2(n13908), .B1(n669), .B2(n14011), .ZN(n9960) );
  OAI22_X1 U5314 ( .A1(n14020), .A2(n13914), .B1(n666), .B2(n14011), .ZN(n9961) );
  OAI22_X1 U5315 ( .A1(n13896), .A2(n13760), .B1(n674), .B2(n13757), .ZN(n9670) );
  OAI22_X1 U5316 ( .A1(n13902), .A2(n13760), .B1(n671), .B2(n13757), .ZN(n9671) );
  OAI22_X1 U5317 ( .A1(n13908), .A2(n13760), .B1(n668), .B2(n13757), .ZN(n9672) );
  OAI22_X1 U5318 ( .A1(n13914), .A2(n13760), .B1(n665), .B2(n13757), .ZN(n9673) );
  OAI22_X1 U5319 ( .A1(n13920), .A2(n13760), .B1(n662), .B2(n13757), .ZN(n9674) );
  OAI22_X1 U5320 ( .A1(n13926), .A2(n13760), .B1(n659), .B2(n13757), .ZN(n9675) );
  OAI22_X1 U5321 ( .A1(n13932), .A2(n13760), .B1(n656), .B2(n13757), .ZN(n9676) );
  OAI22_X1 U5322 ( .A1(n13938), .A2(n13760), .B1(n653), .B2(n13757), .ZN(n9677) );
  OAI22_X1 U5323 ( .A1(n14021), .A2(n13824), .B1(n711), .B2(n14010), .ZN(n9946) );
  OAI22_X1 U5324 ( .A1(n14021), .A2(n13830), .B1(n708), .B2(n14010), .ZN(n9947) );
  OAI22_X1 U5325 ( .A1(n14021), .A2(n13836), .B1(n705), .B2(n14010), .ZN(n9948) );
  OAI22_X1 U5326 ( .A1(n14021), .A2(n13842), .B1(n702), .B2(n14010), .ZN(n9949) );
  OAI22_X1 U5327 ( .A1(n14021), .A2(n13848), .B1(n699), .B2(n14010), .ZN(n9950) );
  OAI22_X1 U5328 ( .A1(n14021), .A2(n13854), .B1(n696), .B2(n14010), .ZN(n9951) );
  OAI22_X1 U5329 ( .A1(n14021), .A2(n13860), .B1(n693), .B2(n14010), .ZN(n9952) );
  OAI22_X1 U5330 ( .A1(n14021), .A2(n13866), .B1(n690), .B2(n14010), .ZN(n9953) );
  OAI22_X1 U5331 ( .A1(n14020), .A2(n13872), .B1(n687), .B2(n14010), .ZN(n9954) );
  OAI22_X1 U5332 ( .A1(n14020), .A2(n13878), .B1(n684), .B2(n14010), .ZN(n9955) );
  OAI22_X1 U5333 ( .A1(n14020), .A2(n13884), .B1(n681), .B2(n14010), .ZN(n9956) );
  OAI22_X1 U5334 ( .A1(n14020), .A2(n13890), .B1(n678), .B2(n14010), .ZN(n9957) );
  OAI22_X1 U5335 ( .A1(n13824), .A2(n13797), .B1(n5387), .B2(n13792), .ZN(
        n9850) );
  OAI22_X1 U5336 ( .A1(n13830), .A2(n13797), .B1(n5397), .B2(n13792), .ZN(
        n9851) );
  OAI22_X1 U5337 ( .A1(n13836), .A2(n13797), .B1(n5407), .B2(n13792), .ZN(
        n9852) );
  OAI22_X1 U5338 ( .A1(n13842), .A2(n13797), .B1(n5417), .B2(n13792), .ZN(
        n9853) );
  OAI22_X1 U5339 ( .A1(n13848), .A2(n13797), .B1(n5427), .B2(n13792), .ZN(
        n9854) );
  OAI22_X1 U5340 ( .A1(n13854), .A2(n13797), .B1(n5437), .B2(n13792), .ZN(
        n9855) );
  OAI22_X1 U5341 ( .A1(n13860), .A2(n13797), .B1(n5447), .B2(n13792), .ZN(
        n9856) );
  OAI22_X1 U5342 ( .A1(n13866), .A2(n13797), .B1(n5457), .B2(n13792), .ZN(
        n9857) );
  OAI22_X1 U5343 ( .A1(n13872), .A2(n13796), .B1(n5467), .B2(n13792), .ZN(
        n9858) );
  OAI22_X1 U5344 ( .A1(n13878), .A2(n13796), .B1(n5477), .B2(n13792), .ZN(
        n9859) );
  OAI22_X1 U5345 ( .A1(n13884), .A2(n13796), .B1(n5487), .B2(n13792), .ZN(
        n9860) );
  OAI22_X1 U5346 ( .A1(n13890), .A2(n13796), .B1(n5497), .B2(n13792), .ZN(
        n9861) );
  OAI22_X1 U5347 ( .A1(n13896), .A2(n13796), .B1(n5507), .B2(n13793), .ZN(
        n9862) );
  OAI22_X1 U5348 ( .A1(n13902), .A2(n13796), .B1(n5517), .B2(n13793), .ZN(
        n9863) );
  OAI22_X1 U5349 ( .A1(n13908), .A2(n13796), .B1(n5527), .B2(n13793), .ZN(
        n9864) );
  OAI22_X1 U5350 ( .A1(n13914), .A2(n13796), .B1(n5537), .B2(n13793), .ZN(
        n9865) );
  OAI22_X1 U5351 ( .A1(n13920), .A2(n13796), .B1(n5547), .B2(n13793), .ZN(
        n9866) );
  OAI22_X1 U5352 ( .A1(n13926), .A2(n13796), .B1(n5557), .B2(n13793), .ZN(
        n9867) );
  OAI22_X1 U5353 ( .A1(n13932), .A2(n13796), .B1(n5567), .B2(n13793), .ZN(
        n9868) );
  OAI22_X1 U5354 ( .A1(n13938), .A2(n13796), .B1(n5577), .B2(n13793), .ZN(
        n9869) );
  OAI22_X1 U5355 ( .A1(n13944), .A2(n13795), .B1(n5587), .B2(n13793), .ZN(
        n9870) );
  OAI22_X1 U5356 ( .A1(n13950), .A2(n13795), .B1(n5597), .B2(n13793), .ZN(
        n9871) );
  OAI22_X1 U5357 ( .A1(n13956), .A2(n13795), .B1(n5607), .B2(n13793), .ZN(
        n9872) );
  OAI22_X1 U5358 ( .A1(n13962), .A2(n13795), .B1(n5617), .B2(n13793), .ZN(
        n9873) );
  OAI22_X1 U5359 ( .A1(n13824), .A2(n13761), .B1(n710), .B2(n13756), .ZN(n9658) );
  OAI22_X1 U5360 ( .A1(n13830), .A2(n13761), .B1(n707), .B2(n13756), .ZN(n9659) );
  OAI22_X1 U5361 ( .A1(n13836), .A2(n13761), .B1(n704), .B2(n13756), .ZN(n9660) );
  OAI22_X1 U5362 ( .A1(n13842), .A2(n13761), .B1(n701), .B2(n13756), .ZN(n9661) );
  OAI22_X1 U5363 ( .A1(n13848), .A2(n13761), .B1(n698), .B2(n13756), .ZN(n9662) );
  OAI22_X1 U5364 ( .A1(n13854), .A2(n13761), .B1(n695), .B2(n13756), .ZN(n9663) );
  OAI22_X1 U5365 ( .A1(n13860), .A2(n13761), .B1(n692), .B2(n13756), .ZN(n9664) );
  OAI22_X1 U5366 ( .A1(n13866), .A2(n13761), .B1(n689), .B2(n13756), .ZN(n9665) );
  OAI22_X1 U5367 ( .A1(n13872), .A2(n13760), .B1(n686), .B2(n13756), .ZN(n9666) );
  OAI22_X1 U5368 ( .A1(n13878), .A2(n13760), .B1(n683), .B2(n13756), .ZN(n9667) );
  OAI22_X1 U5369 ( .A1(n13884), .A2(n13760), .B1(n680), .B2(n13756), .ZN(n9668) );
  OAI22_X1 U5370 ( .A1(n13890), .A2(n13760), .B1(n677), .B2(n13756), .ZN(n9669) );
  OAI22_X1 U5371 ( .A1(n13824), .A2(n13743), .B1(n5385), .B2(n13738), .ZN(
        n9562) );
  OAI22_X1 U5372 ( .A1(n13831), .A2(n13743), .B1(n5395), .B2(n13738), .ZN(
        n9563) );
  OAI22_X1 U5373 ( .A1(n13837), .A2(n13743), .B1(n5405), .B2(n13738), .ZN(
        n9564) );
  OAI22_X1 U5374 ( .A1(n13843), .A2(n13743), .B1(n5415), .B2(n13738), .ZN(
        n9565) );
  OAI22_X1 U5375 ( .A1(n13849), .A2(n13743), .B1(n5425), .B2(n13738), .ZN(
        n9566) );
  OAI22_X1 U5376 ( .A1(n13855), .A2(n13743), .B1(n5435), .B2(n13738), .ZN(
        n9567) );
  OAI22_X1 U5377 ( .A1(n13861), .A2(n13743), .B1(n5445), .B2(n13738), .ZN(
        n9568) );
  OAI22_X1 U5378 ( .A1(n13867), .A2(n13743), .B1(n5455), .B2(n13738), .ZN(
        n9569) );
  OAI22_X1 U5379 ( .A1(n13873), .A2(n13742), .B1(n5465), .B2(n13738), .ZN(
        n9570) );
  OAI22_X1 U5380 ( .A1(n13879), .A2(n13742), .B1(n5475), .B2(n13738), .ZN(
        n9571) );
  OAI22_X1 U5381 ( .A1(n13885), .A2(n13742), .B1(n5485), .B2(n13738), .ZN(
        n9572) );
  OAI22_X1 U5382 ( .A1(n13891), .A2(n13742), .B1(n5495), .B2(n13738), .ZN(
        n9573) );
  OAI22_X1 U5383 ( .A1(n13897), .A2(n13742), .B1(n5505), .B2(n13739), .ZN(
        n9574) );
  OAI22_X1 U5384 ( .A1(n13903), .A2(n13742), .B1(n5515), .B2(n13739), .ZN(
        n9575) );
  OAI22_X1 U5385 ( .A1(n13909), .A2(n13742), .B1(n5525), .B2(n13739), .ZN(
        n9576) );
  OAI22_X1 U5386 ( .A1(n13915), .A2(n13742), .B1(n5535), .B2(n13739), .ZN(
        n9577) );
  OAI22_X1 U5387 ( .A1(n13921), .A2(n13742), .B1(n5545), .B2(n13739), .ZN(
        n9578) );
  OAI22_X1 U5388 ( .A1(n13927), .A2(n13742), .B1(n5555), .B2(n13739), .ZN(
        n9579) );
  OAI22_X1 U5389 ( .A1(n13933), .A2(n13742), .B1(n5565), .B2(n13739), .ZN(
        n9580) );
  OAI22_X1 U5390 ( .A1(n13939), .A2(n13742), .B1(n5575), .B2(n13739), .ZN(
        n9581) );
  OAI22_X1 U5391 ( .A1(n13945), .A2(n13741), .B1(n5585), .B2(n13739), .ZN(
        n9582) );
  OAI22_X1 U5392 ( .A1(n13951), .A2(n13741), .B1(n5595), .B2(n13739), .ZN(
        n9583) );
  OAI22_X1 U5393 ( .A1(n13957), .A2(n13741), .B1(n5605), .B2(n13739), .ZN(
        n9584) );
  OAI22_X1 U5394 ( .A1(n13963), .A2(n13741), .B1(n5615), .B2(n13739), .ZN(
        n9585) );
  OAI22_X1 U5395 ( .A1(n13944), .A2(n13759), .B1(n6938), .B2(n13757), .ZN(
        n9678) );
  OAI22_X1 U5396 ( .A1(n13950), .A2(n13759), .B1(n6939), .B2(n13757), .ZN(
        n9679) );
  OAI22_X1 U5397 ( .A1(n13956), .A2(n13759), .B1(n6940), .B2(n13757), .ZN(
        n9680) );
  OAI22_X1 U5398 ( .A1(n13962), .A2(n13759), .B1(n6941), .B2(n13757), .ZN(
        n9681) );
  OAI22_X1 U5399 ( .A1(n14020), .A2(n13920), .B1(n6922), .B2(n14011), .ZN(
        n9962) );
  OAI22_X1 U5400 ( .A1(n14020), .A2(n13926), .B1(n6923), .B2(n14011), .ZN(
        n9963) );
  OAI22_X1 U5401 ( .A1(n14020), .A2(n13932), .B1(n6924), .B2(n14011), .ZN(
        n9964) );
  OAI22_X1 U5402 ( .A1(n14020), .A2(n13938), .B1(n6925), .B2(n14011), .ZN(
        n9965) );
  OAI22_X1 U5403 ( .A1(n14019), .A2(n13944), .B1(n6926), .B2(n14011), .ZN(
        n9966) );
  OAI22_X1 U5404 ( .A1(n14019), .A2(n13950), .B1(n6927), .B2(n14011), .ZN(
        n9967) );
  OAI22_X1 U5405 ( .A1(n14019), .A2(n13956), .B1(n6928), .B2(n14011), .ZN(
        n9968) );
  OAI22_X1 U5406 ( .A1(n14019), .A2(n13962), .B1(n6929), .B2(n14011), .ZN(
        n9969) );
  OAI22_X1 U5407 ( .A1(n13824), .A2(n13755), .B1(n6870), .B2(n13750), .ZN(
        n9626) );
  OAI22_X1 U5408 ( .A1(n13831), .A2(n13755), .B1(n6871), .B2(n13750), .ZN(
        n9627) );
  OAI22_X1 U5409 ( .A1(n13837), .A2(n13755), .B1(n6872), .B2(n13750), .ZN(
        n9628) );
  OAI22_X1 U5410 ( .A1(n13843), .A2(n13755), .B1(n6873), .B2(n13750), .ZN(
        n9629) );
  OAI22_X1 U5411 ( .A1(n13849), .A2(n13755), .B1(n6874), .B2(n13750), .ZN(
        n9630) );
  OAI22_X1 U5412 ( .A1(n13855), .A2(n13755), .B1(n6875), .B2(n13750), .ZN(
        n9631) );
  OAI22_X1 U5413 ( .A1(n13861), .A2(n13755), .B1(n6876), .B2(n13750), .ZN(
        n9632) );
  OAI22_X1 U5414 ( .A1(n13867), .A2(n13755), .B1(n6877), .B2(n13750), .ZN(
        n9633) );
  OAI22_X1 U5415 ( .A1(n13873), .A2(n13754), .B1(n6878), .B2(n13750), .ZN(
        n9634) );
  OAI22_X1 U5416 ( .A1(n13879), .A2(n13754), .B1(n6879), .B2(n13750), .ZN(
        n9635) );
  OAI22_X1 U5417 ( .A1(n13885), .A2(n13754), .B1(n6880), .B2(n13750), .ZN(
        n9636) );
  OAI22_X1 U5418 ( .A1(n13891), .A2(n13754), .B1(n6881), .B2(n13750), .ZN(
        n9637) );
  OAI22_X1 U5419 ( .A1(n13897), .A2(n13754), .B1(n6882), .B2(n13751), .ZN(
        n9638) );
  OAI22_X1 U5420 ( .A1(n13903), .A2(n13754), .B1(n6884), .B2(n13751), .ZN(
        n9639) );
  OAI22_X1 U5421 ( .A1(n13909), .A2(n13754), .B1(n6886), .B2(n13751), .ZN(
        n9640) );
  OAI22_X1 U5422 ( .A1(n13915), .A2(n13754), .B1(n6888), .B2(n13751), .ZN(
        n9641) );
  OAI22_X1 U5423 ( .A1(n13921), .A2(n13754), .B1(n6890), .B2(n13751), .ZN(
        n9642) );
  OAI22_X1 U5424 ( .A1(n13927), .A2(n13754), .B1(n6891), .B2(n13751), .ZN(
        n9643) );
  OAI22_X1 U5425 ( .A1(n13933), .A2(n13754), .B1(n6892), .B2(n13751), .ZN(
        n9644) );
  OAI22_X1 U5426 ( .A1(n13939), .A2(n13754), .B1(n6893), .B2(n13751), .ZN(
        n9645) );
  OAI22_X1 U5427 ( .A1(n13945), .A2(n13753), .B1(n6810), .B2(n13751), .ZN(
        n9646) );
  OAI22_X1 U5428 ( .A1(n13951), .A2(n13753), .B1(n6811), .B2(n13751), .ZN(
        n9647) );
  OAI22_X1 U5429 ( .A1(n13957), .A2(n13753), .B1(n6812), .B2(n13751), .ZN(
        n9648) );
  OAI22_X1 U5430 ( .A1(n13963), .A2(n13753), .B1(n6813), .B2(n13751), .ZN(
        n9649) );
  OAI22_X1 U5431 ( .A1(n13824), .A2(n13809), .B1(n6830), .B2(n13804), .ZN(
        n9914) );
  OAI22_X1 U5432 ( .A1(n13830), .A2(n13809), .B1(n6831), .B2(n13804), .ZN(
        n9915) );
  OAI22_X1 U5433 ( .A1(n13836), .A2(n13809), .B1(n6832), .B2(n13804), .ZN(
        n9916) );
  OAI22_X1 U5434 ( .A1(n13842), .A2(n13809), .B1(n6833), .B2(n13804), .ZN(
        n9917) );
  OAI22_X1 U5435 ( .A1(n13848), .A2(n13809), .B1(n6834), .B2(n13804), .ZN(
        n9918) );
  OAI22_X1 U5436 ( .A1(n13854), .A2(n13809), .B1(n6835), .B2(n13804), .ZN(
        n9919) );
  OAI22_X1 U5437 ( .A1(n13860), .A2(n13809), .B1(n6836), .B2(n13804), .ZN(
        n9920) );
  OAI22_X1 U5438 ( .A1(n13866), .A2(n13809), .B1(n6837), .B2(n13804), .ZN(
        n9921) );
  OAI22_X1 U5439 ( .A1(n13872), .A2(n13808), .B1(n6838), .B2(n13804), .ZN(
        n9922) );
  OAI22_X1 U5440 ( .A1(n13878), .A2(n13808), .B1(n6839), .B2(n13804), .ZN(
        n9923) );
  OAI22_X1 U5441 ( .A1(n13884), .A2(n13808), .B1(n6840), .B2(n13804), .ZN(
        n9924) );
  OAI22_X1 U5442 ( .A1(n13890), .A2(n13808), .B1(n6841), .B2(n13804), .ZN(
        n9925) );
  OAI22_X1 U5443 ( .A1(n13896), .A2(n13808), .B1(n6883), .B2(n13805), .ZN(
        n9926) );
  OAI22_X1 U5444 ( .A1(n13902), .A2(n13808), .B1(n6885), .B2(n13805), .ZN(
        n9927) );
  OAI22_X1 U5445 ( .A1(n13908), .A2(n13808), .B1(n6887), .B2(n13805), .ZN(
        n9928) );
  OAI22_X1 U5446 ( .A1(n13914), .A2(n13808), .B1(n6889), .B2(n13805), .ZN(
        n9929) );
  OAI22_X1 U5447 ( .A1(n13920), .A2(n13808), .B1(n6794), .B2(n13805), .ZN(
        n9930) );
  OAI22_X1 U5448 ( .A1(n13926), .A2(n13808), .B1(n6795), .B2(n13805), .ZN(
        n9931) );
  OAI22_X1 U5449 ( .A1(n13932), .A2(n13808), .B1(n6796), .B2(n13805), .ZN(
        n9932) );
  OAI22_X1 U5450 ( .A1(n13938), .A2(n13808), .B1(n6797), .B2(n13805), .ZN(
        n9933) );
  OAI22_X1 U5451 ( .A1(n13944), .A2(n13807), .B1(n6798), .B2(n13805), .ZN(
        n9934) );
  OAI22_X1 U5452 ( .A1(n13950), .A2(n13807), .B1(n6799), .B2(n13805), .ZN(
        n9935) );
  OAI22_X1 U5453 ( .A1(n13956), .A2(n13807), .B1(n6800), .B2(n13805), .ZN(
        n9936) );
  OAI22_X1 U5454 ( .A1(n13962), .A2(n13807), .B1(n6801), .B2(n13805), .ZN(
        n9937) );
  OAI22_X1 U5455 ( .A1(n13939), .A2(n13694), .B1(n5776), .B2(n13691), .ZN(
        n9325) );
  OAI22_X1 U5456 ( .A1(n13824), .A2(n13791), .B1(n840), .B2(n13786), .ZN(n9818) );
  OAI22_X1 U5457 ( .A1(n13830), .A2(n13791), .B1(n839), .B2(n13786), .ZN(n9819) );
  OAI22_X1 U5458 ( .A1(n13836), .A2(n13791), .B1(n838), .B2(n13786), .ZN(n9820) );
  OAI22_X1 U5459 ( .A1(n13842), .A2(n13791), .B1(n837), .B2(n13786), .ZN(n9821) );
  OAI22_X1 U5460 ( .A1(n13848), .A2(n13791), .B1(n836), .B2(n13786), .ZN(n9822) );
  OAI22_X1 U5461 ( .A1(n13854), .A2(n13791), .B1(n835), .B2(n13786), .ZN(n9823) );
  OAI22_X1 U5462 ( .A1(n13860), .A2(n13791), .B1(n834), .B2(n13786), .ZN(n9824) );
  OAI22_X1 U5463 ( .A1(n13866), .A2(n13791), .B1(n833), .B2(n13786), .ZN(n9825) );
  OAI22_X1 U5464 ( .A1(n13872), .A2(n13790), .B1(n832), .B2(n13786), .ZN(n9826) );
  OAI22_X1 U5465 ( .A1(n13878), .A2(n13790), .B1(n831), .B2(n13786), .ZN(n9827) );
  OAI22_X1 U5466 ( .A1(n13884), .A2(n13790), .B1(n830), .B2(n13786), .ZN(n9828) );
  OAI22_X1 U5467 ( .A1(n13890), .A2(n13790), .B1(n829), .B2(n13786), .ZN(n9829) );
  OAI22_X1 U5468 ( .A1(n13896), .A2(n13790), .B1(n828), .B2(n13787), .ZN(n9830) );
  OAI22_X1 U5469 ( .A1(n13902), .A2(n13790), .B1(n827), .B2(n13787), .ZN(n9831) );
  OAI22_X1 U5470 ( .A1(n13908), .A2(n13790), .B1(n826), .B2(n13787), .ZN(n9832) );
  OAI22_X1 U5471 ( .A1(n13914), .A2(n13790), .B1(n825), .B2(n13787), .ZN(n9833) );
  OAI22_X1 U5472 ( .A1(n13920), .A2(n13790), .B1(n824), .B2(n13787), .ZN(n9834) );
  OAI22_X1 U5473 ( .A1(n13926), .A2(n13790), .B1(n823), .B2(n13787), .ZN(n9835) );
  OAI22_X1 U5474 ( .A1(n13932), .A2(n13790), .B1(n822), .B2(n13787), .ZN(n9836) );
  OAI22_X1 U5475 ( .A1(n13938), .A2(n13790), .B1(n821), .B2(n13787), .ZN(n9837) );
  OAI22_X1 U5476 ( .A1(n13944), .A2(n13789), .B1(n820), .B2(n13787), .ZN(n9838) );
  OAI22_X1 U5477 ( .A1(n13950), .A2(n13789), .B1(n819), .B2(n13787), .ZN(n9839) );
  OAI22_X1 U5478 ( .A1(n13956), .A2(n13789), .B1(n818), .B2(n13787), .ZN(n9840) );
  OAI22_X1 U5479 ( .A1(n13962), .A2(n13789), .B1(n817), .B2(n13787), .ZN(n9841) );
  OAI22_X1 U5480 ( .A1(n13825), .A2(n13737), .B1(n872), .B2(n13732), .ZN(n9530) );
  OAI22_X1 U5481 ( .A1(n13831), .A2(n13737), .B1(n871), .B2(n13732), .ZN(n9531) );
  OAI22_X1 U5482 ( .A1(n13837), .A2(n13737), .B1(n870), .B2(n13732), .ZN(n9532) );
  OAI22_X1 U5483 ( .A1(n13843), .A2(n13737), .B1(n869), .B2(n13732), .ZN(n9533) );
  OAI22_X1 U5484 ( .A1(n13849), .A2(n13737), .B1(n868), .B2(n13732), .ZN(n9534) );
  OAI22_X1 U5485 ( .A1(n13855), .A2(n13737), .B1(n867), .B2(n13732), .ZN(n9535) );
  OAI22_X1 U5486 ( .A1(n13861), .A2(n13737), .B1(n866), .B2(n13732), .ZN(n9536) );
  OAI22_X1 U5487 ( .A1(n13867), .A2(n13737), .B1(n865), .B2(n13732), .ZN(n9537) );
  OAI22_X1 U5488 ( .A1(n13873), .A2(n13736), .B1(n864), .B2(n13732), .ZN(n9538) );
  OAI22_X1 U5489 ( .A1(n13879), .A2(n13736), .B1(n863), .B2(n13732), .ZN(n9539) );
  OAI22_X1 U5490 ( .A1(n13885), .A2(n13736), .B1(n862), .B2(n13732), .ZN(n9540) );
  OAI22_X1 U5491 ( .A1(n13891), .A2(n13736), .B1(n861), .B2(n13732), .ZN(n9541) );
  OAI22_X1 U5492 ( .A1(n13897), .A2(n13736), .B1(n860), .B2(n13733), .ZN(n9542) );
  OAI22_X1 U5493 ( .A1(n13903), .A2(n13736), .B1(n859), .B2(n13733), .ZN(n9543) );
  OAI22_X1 U5494 ( .A1(n13909), .A2(n13736), .B1(n858), .B2(n13733), .ZN(n9544) );
  OAI22_X1 U5495 ( .A1(n13915), .A2(n13736), .B1(n857), .B2(n13733), .ZN(n9545) );
  OAI22_X1 U5496 ( .A1(n13921), .A2(n13736), .B1(n856), .B2(n13733), .ZN(n9546) );
  OAI22_X1 U5497 ( .A1(n13927), .A2(n13736), .B1(n855), .B2(n13733), .ZN(n9547) );
  OAI22_X1 U5498 ( .A1(n13933), .A2(n13736), .B1(n854), .B2(n13733), .ZN(n9548) );
  OAI22_X1 U5499 ( .A1(n13939), .A2(n13736), .B1(n853), .B2(n13733), .ZN(n9549) );
  OAI22_X1 U5500 ( .A1(n13945), .A2(n13735), .B1(n852), .B2(n13733), .ZN(n9550) );
  OAI22_X1 U5501 ( .A1(n13951), .A2(n13735), .B1(n851), .B2(n13733), .ZN(n9551) );
  OAI22_X1 U5502 ( .A1(n13957), .A2(n13735), .B1(n850), .B2(n13733), .ZN(n9552) );
  OAI22_X1 U5503 ( .A1(n13963), .A2(n13735), .B1(n849), .B2(n13733), .ZN(n9553) );
  OAI22_X1 U5504 ( .A1(n13945), .A2(n13693), .B1(n5780), .B2(n13691), .ZN(
        n9326) );
  OAI22_X1 U5505 ( .A1(n13951), .A2(n13693), .B1(n5784), .B2(n13691), .ZN(
        n9327) );
  OAI22_X1 U5506 ( .A1(n13957), .A2(n13693), .B1(n5788), .B2(n13691), .ZN(
        n9328) );
  OAI22_X1 U5507 ( .A1(n13963), .A2(n13693), .B1(n5792), .B2(n13691), .ZN(
        n9329) );
  OAI22_X1 U5508 ( .A1(n13825), .A2(n13689), .B1(n5701), .B2(n13684), .ZN(
        n9274) );
  OAI22_X1 U5509 ( .A1(n13831), .A2(n13689), .B1(n5705), .B2(n13684), .ZN(
        n9275) );
  OAI22_X1 U5510 ( .A1(n13837), .A2(n13689), .B1(n5709), .B2(n13684), .ZN(
        n9276) );
  OAI22_X1 U5511 ( .A1(n13843), .A2(n13689), .B1(n5713), .B2(n13684), .ZN(
        n9277) );
  OAI22_X1 U5512 ( .A1(n13849), .A2(n13689), .B1(n5717), .B2(n13684), .ZN(
        n9278) );
  OAI22_X1 U5513 ( .A1(n13855), .A2(n13689), .B1(n5721), .B2(n13684), .ZN(
        n9279) );
  OAI22_X1 U5514 ( .A1(n13861), .A2(n13689), .B1(n5725), .B2(n13684), .ZN(
        n9280) );
  OAI22_X1 U5515 ( .A1(n13867), .A2(n13689), .B1(n5729), .B2(n13684), .ZN(
        n9281) );
  OAI22_X1 U5516 ( .A1(n13873), .A2(n13688), .B1(n5733), .B2(n13684), .ZN(
        n9282) );
  OAI22_X1 U5517 ( .A1(n13879), .A2(n13688), .B1(n5737), .B2(n13684), .ZN(
        n9283) );
  OAI22_X1 U5518 ( .A1(n13885), .A2(n13688), .B1(n5741), .B2(n13684), .ZN(
        n9284) );
  OAI22_X1 U5519 ( .A1(n13891), .A2(n13688), .B1(n5745), .B2(n13684), .ZN(
        n9285) );
  OAI22_X1 U5520 ( .A1(n13897), .A2(n13688), .B1(n5749), .B2(n13685), .ZN(
        n9286) );
  OAI22_X1 U5521 ( .A1(n13903), .A2(n13688), .B1(n5753), .B2(n13685), .ZN(
        n9287) );
  OAI22_X1 U5522 ( .A1(n13909), .A2(n13688), .B1(n5757), .B2(n13685), .ZN(
        n9288) );
  OAI22_X1 U5523 ( .A1(n13915), .A2(n13688), .B1(n5761), .B2(n13685), .ZN(
        n9289) );
  OAI22_X1 U5524 ( .A1(n13921), .A2(n13688), .B1(n5765), .B2(n13685), .ZN(
        n9290) );
  OAI22_X1 U5525 ( .A1(n13927), .A2(n13688), .B1(n5769), .B2(n13685), .ZN(
        n9291) );
  OAI22_X1 U5526 ( .A1(n13933), .A2(n13688), .B1(n5773), .B2(n13685), .ZN(
        n9292) );
  OAI22_X1 U5527 ( .A1(n13939), .A2(n13688), .B1(n5777), .B2(n13685), .ZN(
        n9293) );
  OAI22_X1 U5528 ( .A1(n13945), .A2(n13687), .B1(n5781), .B2(n13685), .ZN(
        n9294) );
  OAI22_X1 U5529 ( .A1(n13951), .A2(n13687), .B1(n5785), .B2(n13685), .ZN(
        n9295) );
  OAI22_X1 U5530 ( .A1(n13957), .A2(n13687), .B1(n5789), .B2(n13685), .ZN(
        n9296) );
  OAI22_X1 U5531 ( .A1(n13963), .A2(n13687), .B1(n5793), .B2(n13685), .ZN(
        n9297) );
  OAI22_X1 U5532 ( .A1(n13825), .A2(n13683), .B1(n904), .B2(n13678), .ZN(n9242) );
  OAI22_X1 U5533 ( .A1(n13831), .A2(n13683), .B1(n903), .B2(n13678), .ZN(n9243) );
  OAI22_X1 U5534 ( .A1(n13837), .A2(n13683), .B1(n902), .B2(n13678), .ZN(n9244) );
  OAI22_X1 U5535 ( .A1(n13843), .A2(n13683), .B1(n901), .B2(n13678), .ZN(n9245) );
  OAI22_X1 U5536 ( .A1(n13849), .A2(n13683), .B1(n900), .B2(n13678), .ZN(n9246) );
  OAI22_X1 U5537 ( .A1(n13855), .A2(n13683), .B1(n899), .B2(n13678), .ZN(n9247) );
  OAI22_X1 U5538 ( .A1(n13861), .A2(n13683), .B1(n898), .B2(n13678), .ZN(n9248) );
  OAI22_X1 U5539 ( .A1(n13867), .A2(n13683), .B1(n897), .B2(n13678), .ZN(n9249) );
  OAI22_X1 U5540 ( .A1(n13873), .A2(n13682), .B1(n896), .B2(n13678), .ZN(n9250) );
  OAI22_X1 U5541 ( .A1(n13879), .A2(n13682), .B1(n895), .B2(n13678), .ZN(n9251) );
  OAI22_X1 U5542 ( .A1(n13885), .A2(n13682), .B1(n894), .B2(n13678), .ZN(n9252) );
  OAI22_X1 U5543 ( .A1(n13891), .A2(n13682), .B1(n893), .B2(n13678), .ZN(n9253) );
  OAI22_X1 U5544 ( .A1(n13897), .A2(n13682), .B1(n892), .B2(n13679), .ZN(n9254) );
  OAI22_X1 U5545 ( .A1(n13903), .A2(n13682), .B1(n891), .B2(n13679), .ZN(n9255) );
  OAI22_X1 U5546 ( .A1(n13909), .A2(n13682), .B1(n890), .B2(n13679), .ZN(n9256) );
  OAI22_X1 U5547 ( .A1(n13915), .A2(n13682), .B1(n889), .B2(n13679), .ZN(n9257) );
  OAI22_X1 U5548 ( .A1(n13921), .A2(n13682), .B1(n888), .B2(n13679), .ZN(n9258) );
  OAI22_X1 U5549 ( .A1(n13927), .A2(n13682), .B1(n887), .B2(n13679), .ZN(n9259) );
  OAI22_X1 U5550 ( .A1(n13933), .A2(n13682), .B1(n886), .B2(n13679), .ZN(n9260) );
  OAI22_X1 U5551 ( .A1(n13939), .A2(n13682), .B1(n885), .B2(n13679), .ZN(n9261) );
  OAI22_X1 U5552 ( .A1(n13945), .A2(n13681), .B1(n884), .B2(n13679), .ZN(n9262) );
  OAI22_X1 U5553 ( .A1(n13951), .A2(n13681), .B1(n883), .B2(n13679), .ZN(n9263) );
  OAI22_X1 U5554 ( .A1(n13957), .A2(n13681), .B1(n882), .B2(n13679), .ZN(n9264) );
  OAI22_X1 U5555 ( .A1(n13963), .A2(n13681), .B1(n881), .B2(n13679), .ZN(n9265) );
  OAI22_X1 U5556 ( .A1(n13874), .A2(n13640), .B1(n5462), .B2(n13636), .ZN(
        n9026) );
  OAI22_X1 U5557 ( .A1(n13880), .A2(n13640), .B1(n5472), .B2(n13636), .ZN(
        n9027) );
  OAI22_X1 U5558 ( .A1(n13886), .A2(n13640), .B1(n5482), .B2(n13636), .ZN(
        n9028) );
  OAI22_X1 U5559 ( .A1(n13892), .A2(n13640), .B1(n5492), .B2(n13636), .ZN(
        n9029) );
  OAI22_X1 U5560 ( .A1(n13898), .A2(n13640), .B1(n5502), .B2(n13637), .ZN(
        n9030) );
  OAI22_X1 U5561 ( .A1(n13904), .A2(n13640), .B1(n5512), .B2(n13637), .ZN(
        n9031) );
  OAI22_X1 U5562 ( .A1(n13910), .A2(n13640), .B1(n5522), .B2(n13637), .ZN(
        n9032) );
  OAI22_X1 U5563 ( .A1(n13916), .A2(n13640), .B1(n5532), .B2(n13637), .ZN(
        n9033) );
  OAI22_X1 U5564 ( .A1(n13922), .A2(n13640), .B1(n5542), .B2(n13637), .ZN(
        n9034) );
  OAI22_X1 U5565 ( .A1(n13928), .A2(n13640), .B1(n5552), .B2(n13637), .ZN(
        n9035) );
  OAI22_X1 U5566 ( .A1(n13934), .A2(n13640), .B1(n5562), .B2(n13637), .ZN(
        n9036) );
  OAI22_X1 U5567 ( .A1(n13940), .A2(n13640), .B1(n5572), .B2(n13637), .ZN(
        n9037) );
  OAI22_X1 U5568 ( .A1(n13946), .A2(n13639), .B1(n5582), .B2(n13637), .ZN(
        n9038) );
  OAI22_X1 U5569 ( .A1(n13952), .A2(n13639), .B1(n5592), .B2(n13637), .ZN(
        n9039) );
  OAI22_X1 U5570 ( .A1(n13958), .A2(n13639), .B1(n5602), .B2(n13637), .ZN(
        n9040) );
  OAI22_X1 U5571 ( .A1(n13964), .A2(n13639), .B1(n5612), .B2(n13637), .ZN(
        n9041) );
  OAI22_X1 U5572 ( .A1(n13826), .A2(n13635), .B1(n5383), .B2(n13630), .ZN(
        n8986) );
  OAI22_X1 U5573 ( .A1(n13832), .A2(n13635), .B1(n5393), .B2(n13630), .ZN(
        n8987) );
  OAI22_X1 U5574 ( .A1(n13838), .A2(n13635), .B1(n5403), .B2(n13630), .ZN(
        n8988) );
  OAI22_X1 U5575 ( .A1(n13844), .A2(n13635), .B1(n5413), .B2(n13630), .ZN(
        n8989) );
  OAI22_X1 U5576 ( .A1(n13850), .A2(n13635), .B1(n5423), .B2(n13630), .ZN(
        n8990) );
  OAI22_X1 U5577 ( .A1(n13856), .A2(n13635), .B1(n5433), .B2(n13630), .ZN(
        n8991) );
  OAI22_X1 U5578 ( .A1(n13862), .A2(n13635), .B1(n5443), .B2(n13630), .ZN(
        n8992) );
  OAI22_X1 U5579 ( .A1(n13868), .A2(n13635), .B1(n5453), .B2(n13630), .ZN(
        n8993) );
  OAI22_X1 U5580 ( .A1(n13874), .A2(n13634), .B1(n5463), .B2(n13630), .ZN(
        n8994) );
  OAI22_X1 U5581 ( .A1(n13880), .A2(n13634), .B1(n5473), .B2(n13630), .ZN(
        n8995) );
  OAI22_X1 U5582 ( .A1(n13886), .A2(n13634), .B1(n5483), .B2(n13630), .ZN(
        n8996) );
  OAI22_X1 U5583 ( .A1(n13892), .A2(n13634), .B1(n5493), .B2(n13630), .ZN(
        n8997) );
  OAI22_X1 U5584 ( .A1(n13898), .A2(n13634), .B1(n5503), .B2(n13631), .ZN(
        n8998) );
  OAI22_X1 U5585 ( .A1(n13904), .A2(n13634), .B1(n5513), .B2(n13631), .ZN(
        n8999) );
  OAI22_X1 U5586 ( .A1(n13910), .A2(n13634), .B1(n5523), .B2(n13631), .ZN(
        n9000) );
  OAI22_X1 U5587 ( .A1(n13916), .A2(n13634), .B1(n5533), .B2(n13631), .ZN(
        n9001) );
  OAI22_X1 U5588 ( .A1(n13922), .A2(n13634), .B1(n5543), .B2(n13631), .ZN(
        n9002) );
  OAI22_X1 U5589 ( .A1(n13928), .A2(n13634), .B1(n5553), .B2(n13631), .ZN(
        n9003) );
  OAI22_X1 U5590 ( .A1(n13934), .A2(n13634), .B1(n5563), .B2(n13631), .ZN(
        n9004) );
  OAI22_X1 U5591 ( .A1(n13940), .A2(n13634), .B1(n5573), .B2(n13631), .ZN(
        n9005) );
  OAI22_X1 U5592 ( .A1(n13946), .A2(n13633), .B1(n5583), .B2(n13631), .ZN(
        n9006) );
  OAI22_X1 U5593 ( .A1(n13952), .A2(n13633), .B1(n5593), .B2(n13631), .ZN(
        n9007) );
  OAI22_X1 U5594 ( .A1(n13958), .A2(n13633), .B1(n5603), .B2(n13631), .ZN(
        n9008) );
  OAI22_X1 U5595 ( .A1(n13964), .A2(n13633), .B1(n5613), .B2(n13631), .ZN(
        n9009) );
  OAI22_X1 U5596 ( .A1(n13826), .A2(n13629), .B1(n936), .B2(n13624), .ZN(n8954) );
  OAI22_X1 U5597 ( .A1(n13832), .A2(n13629), .B1(n935), .B2(n13624), .ZN(n8955) );
  OAI22_X1 U5598 ( .A1(n13838), .A2(n13629), .B1(n934), .B2(n13624), .ZN(n8956) );
  OAI22_X1 U5599 ( .A1(n13844), .A2(n13629), .B1(n933), .B2(n13624), .ZN(n8957) );
  OAI22_X1 U5600 ( .A1(n13850), .A2(n13629), .B1(n932), .B2(n13624), .ZN(n8958) );
  OAI22_X1 U5601 ( .A1(n13856), .A2(n13629), .B1(n931), .B2(n13624), .ZN(n8959) );
  OAI22_X1 U5602 ( .A1(n13862), .A2(n13629), .B1(n930), .B2(n13624), .ZN(n8960) );
  OAI22_X1 U5603 ( .A1(n13868), .A2(n13629), .B1(n929), .B2(n13624), .ZN(n8961) );
  OAI22_X1 U5604 ( .A1(n13874), .A2(n13628), .B1(n928), .B2(n13624), .ZN(n8962) );
  OAI22_X1 U5605 ( .A1(n13880), .A2(n13628), .B1(n927), .B2(n13624), .ZN(n8963) );
  OAI22_X1 U5606 ( .A1(n13886), .A2(n13628), .B1(n926), .B2(n13624), .ZN(n8964) );
  OAI22_X1 U5607 ( .A1(n13892), .A2(n13628), .B1(n925), .B2(n13624), .ZN(n8965) );
  OAI22_X1 U5608 ( .A1(n13898), .A2(n13628), .B1(n924), .B2(n13625), .ZN(n8966) );
  OAI22_X1 U5609 ( .A1(n13904), .A2(n13628), .B1(n923), .B2(n13625), .ZN(n8967) );
  OAI22_X1 U5610 ( .A1(n13910), .A2(n13628), .B1(n922), .B2(n13625), .ZN(n8968) );
  OAI22_X1 U5611 ( .A1(n13916), .A2(n13628), .B1(n921), .B2(n13625), .ZN(n8969) );
  OAI22_X1 U5612 ( .A1(n13922), .A2(n13628), .B1(n920), .B2(n13625), .ZN(n8970) );
  OAI22_X1 U5613 ( .A1(n13928), .A2(n13628), .B1(n919), .B2(n13625), .ZN(n8971) );
  OAI22_X1 U5614 ( .A1(n13934), .A2(n13628), .B1(n918), .B2(n13625), .ZN(n8972) );
  OAI22_X1 U5615 ( .A1(n13940), .A2(n13628), .B1(n917), .B2(n13625), .ZN(n8973) );
  OAI22_X1 U5616 ( .A1(n13946), .A2(n13627), .B1(n916), .B2(n13625), .ZN(n8974) );
  OAI22_X1 U5617 ( .A1(n13952), .A2(n13627), .B1(n915), .B2(n13625), .ZN(n8975) );
  OAI22_X1 U5618 ( .A1(n13958), .A2(n13627), .B1(n914), .B2(n13625), .ZN(n8976) );
  OAI22_X1 U5619 ( .A1(n13964), .A2(n13627), .B1(n913), .B2(n13625), .ZN(n8977) );
  OAI22_X1 U5620 ( .A1(n13947), .A2(n13585), .B1(n5778), .B2(n13582), .ZN(
        n8750) );
  OAI22_X1 U5621 ( .A1(n13953), .A2(n13585), .B1(n5782), .B2(n13582), .ZN(
        n8751) );
  OAI22_X1 U5622 ( .A1(n13959), .A2(n13585), .B1(n5786), .B2(n13582), .ZN(
        n8752) );
  OAI22_X1 U5623 ( .A1(n13965), .A2(n13585), .B1(n5790), .B2(n13582), .ZN(
        n8753) );
  OAI22_X1 U5624 ( .A1(n13971), .A2(n13585), .B1(n5794), .B2(n13582), .ZN(
        n8754) );
  OAI22_X1 U5625 ( .A1(n13977), .A2(n13585), .B1(n5798), .B2(n13582), .ZN(
        n8755) );
  OAI22_X1 U5626 ( .A1(n13983), .A2(n13585), .B1(n5802), .B2(n13582), .ZN(
        n8756) );
  OAI22_X1 U5627 ( .A1(n13989), .A2(n13585), .B1(n5806), .B2(n13582), .ZN(
        n8757) );
  OAI22_X1 U5628 ( .A1(n13995), .A2(n13585), .B1(n5810), .B2(n13582), .ZN(
        n8758) );
  OAI22_X1 U5629 ( .A1(n14001), .A2(n13585), .B1(n5814), .B2(n13582), .ZN(
        n8759) );
  OAI22_X1 U5630 ( .A1(n14007), .A2(n13585), .B1(n5818), .B2(n13582), .ZN(
        n8760) );
  OAI22_X1 U5631 ( .A1(n14016), .A2(n13585), .B1(n5822), .B2(n13582), .ZN(
        n8761) );
  OAI22_X1 U5632 ( .A1(n13827), .A2(n13581), .B1(n5699), .B2(n13576), .ZN(
        n8698) );
  OAI22_X1 U5633 ( .A1(n13833), .A2(n13581), .B1(n5703), .B2(n13576), .ZN(
        n8699) );
  OAI22_X1 U5634 ( .A1(n13839), .A2(n13581), .B1(n5707), .B2(n13576), .ZN(
        n8700) );
  OAI22_X1 U5635 ( .A1(n13845), .A2(n13581), .B1(n5711), .B2(n13576), .ZN(
        n8701) );
  OAI22_X1 U5636 ( .A1(n13851), .A2(n13581), .B1(n5715), .B2(n13576), .ZN(
        n8702) );
  OAI22_X1 U5637 ( .A1(n13857), .A2(n13581), .B1(n5719), .B2(n13576), .ZN(
        n8703) );
  OAI22_X1 U5638 ( .A1(n13863), .A2(n13581), .B1(n5723), .B2(n13576), .ZN(
        n8704) );
  OAI22_X1 U5639 ( .A1(n13869), .A2(n13581), .B1(n5727), .B2(n13576), .ZN(
        n8705) );
  OAI22_X1 U5640 ( .A1(n13875), .A2(n13580), .B1(n5731), .B2(n13576), .ZN(
        n8706) );
  OAI22_X1 U5641 ( .A1(n13881), .A2(n13580), .B1(n5735), .B2(n13576), .ZN(
        n8707) );
  OAI22_X1 U5642 ( .A1(n13887), .A2(n13580), .B1(n5739), .B2(n13576), .ZN(
        n8708) );
  OAI22_X1 U5643 ( .A1(n13893), .A2(n13580), .B1(n5743), .B2(n13576), .ZN(
        n8709) );
  OAI22_X1 U5644 ( .A1(n13899), .A2(n13580), .B1(n5747), .B2(n13577), .ZN(
        n8710) );
  OAI22_X1 U5645 ( .A1(n13905), .A2(n13580), .B1(n5751), .B2(n13577), .ZN(
        n8711) );
  OAI22_X1 U5646 ( .A1(n13911), .A2(n13580), .B1(n5755), .B2(n13577), .ZN(
        n8712) );
  OAI22_X1 U5647 ( .A1(n13917), .A2(n13580), .B1(n5759), .B2(n13577), .ZN(
        n8713) );
  OAI22_X1 U5648 ( .A1(n13923), .A2(n13580), .B1(n5763), .B2(n13577), .ZN(
        n8714) );
  OAI22_X1 U5649 ( .A1(n13929), .A2(n13580), .B1(n5767), .B2(n13577), .ZN(
        n8715) );
  OAI22_X1 U5650 ( .A1(n13935), .A2(n13580), .B1(n5771), .B2(n13577), .ZN(
        n8716) );
  OAI22_X1 U5651 ( .A1(n13941), .A2(n13580), .B1(n5775), .B2(n13577), .ZN(
        n8717) );
  OAI22_X1 U5652 ( .A1(n13947), .A2(n13579), .B1(n5779), .B2(n13577), .ZN(
        n8718) );
  OAI22_X1 U5653 ( .A1(n13953), .A2(n13579), .B1(n5783), .B2(n13577), .ZN(
        n8719) );
  OAI22_X1 U5654 ( .A1(n13959), .A2(n13579), .B1(n5787), .B2(n13577), .ZN(
        n8720) );
  OAI22_X1 U5655 ( .A1(n13965), .A2(n13579), .B1(n5791), .B2(n13577), .ZN(
        n8721) );
  OAI22_X1 U5656 ( .A1(n13827), .A2(n13575), .B1(n968), .B2(n13570), .ZN(n8666) );
  OAI22_X1 U5657 ( .A1(n13833), .A2(n13575), .B1(n967), .B2(n13570), .ZN(n8667) );
  OAI22_X1 U5658 ( .A1(n13839), .A2(n13575), .B1(n966), .B2(n13570), .ZN(n8668) );
  OAI22_X1 U5659 ( .A1(n13845), .A2(n13575), .B1(n965), .B2(n13570), .ZN(n8669) );
  OAI22_X1 U5660 ( .A1(n13851), .A2(n13575), .B1(n964), .B2(n13570), .ZN(n8670) );
  OAI22_X1 U5661 ( .A1(n13857), .A2(n13575), .B1(n963), .B2(n13570), .ZN(n8671) );
  OAI22_X1 U5662 ( .A1(n13863), .A2(n13575), .B1(n962), .B2(n13570), .ZN(n8672) );
  OAI22_X1 U5663 ( .A1(n13869), .A2(n13575), .B1(n961), .B2(n13570), .ZN(n8673) );
  OAI22_X1 U5664 ( .A1(n13875), .A2(n13574), .B1(n960), .B2(n13570), .ZN(n8674) );
  OAI22_X1 U5665 ( .A1(n13881), .A2(n13574), .B1(n959), .B2(n13570), .ZN(n8675) );
  OAI22_X1 U5666 ( .A1(n13887), .A2(n13574), .B1(n958), .B2(n13570), .ZN(n8676) );
  OAI22_X1 U5667 ( .A1(n13893), .A2(n13574), .B1(n957), .B2(n13570), .ZN(n8677) );
  OAI22_X1 U5668 ( .A1(n13899), .A2(n13574), .B1(n956), .B2(n13571), .ZN(n8678) );
  OAI22_X1 U5669 ( .A1(n13905), .A2(n13574), .B1(n955), .B2(n13571), .ZN(n8679) );
  OAI22_X1 U5670 ( .A1(n13911), .A2(n13574), .B1(n954), .B2(n13571), .ZN(n8680) );
  OAI22_X1 U5671 ( .A1(n13917), .A2(n13574), .B1(n953), .B2(n13571), .ZN(n8681) );
  OAI22_X1 U5672 ( .A1(n13923), .A2(n13574), .B1(n952), .B2(n13571), .ZN(n8682) );
  OAI22_X1 U5673 ( .A1(n13929), .A2(n13574), .B1(n951), .B2(n13571), .ZN(n8683) );
  OAI22_X1 U5674 ( .A1(n13935), .A2(n13574), .B1(n950), .B2(n13571), .ZN(n8684) );
  OAI22_X1 U5675 ( .A1(n13941), .A2(n13574), .B1(n949), .B2(n13571), .ZN(n8685) );
  OAI22_X1 U5676 ( .A1(n13947), .A2(n13573), .B1(n948), .B2(n13571), .ZN(n8686) );
  OAI22_X1 U5677 ( .A1(n13953), .A2(n13573), .B1(n947), .B2(n13571), .ZN(n8687) );
  OAI22_X1 U5678 ( .A1(n13959), .A2(n13573), .B1(n946), .B2(n13571), .ZN(n8688) );
  OAI22_X1 U5679 ( .A1(n13965), .A2(n13573), .B1(n945), .B2(n13571), .ZN(n8689) );
  OAI22_X1 U5680 ( .A1(n13827), .A2(n13545), .B1(n712), .B2(n13540), .ZN(n8506) );
  OAI22_X1 U5681 ( .A1(n13833), .A2(n13545), .B1(n709), .B2(n13540), .ZN(n8507) );
  OAI22_X1 U5682 ( .A1(n13839), .A2(n13545), .B1(n706), .B2(n13540), .ZN(n8508) );
  OAI22_X1 U5683 ( .A1(n13845), .A2(n13545), .B1(n703), .B2(n13540), .ZN(n8509) );
  OAI22_X1 U5684 ( .A1(n13851), .A2(n13545), .B1(n700), .B2(n13540), .ZN(n8510) );
  OAI22_X1 U5685 ( .A1(n13857), .A2(n13545), .B1(n697), .B2(n13540), .ZN(n8511) );
  OAI22_X1 U5686 ( .A1(n13863), .A2(n13545), .B1(n694), .B2(n13540), .ZN(n8512) );
  OAI22_X1 U5687 ( .A1(n13869), .A2(n13545), .B1(n691), .B2(n13540), .ZN(n8513) );
  OAI22_X1 U5688 ( .A1(n13875), .A2(n13544), .B1(n688), .B2(n13540), .ZN(n8514) );
  OAI22_X1 U5689 ( .A1(n13881), .A2(n13544), .B1(n685), .B2(n13540), .ZN(n8515) );
  OAI22_X1 U5690 ( .A1(n13887), .A2(n13544), .B1(n682), .B2(n13540), .ZN(n8516) );
  OAI22_X1 U5691 ( .A1(n13893), .A2(n13544), .B1(n679), .B2(n13540), .ZN(n8517) );
  OAI22_X1 U5692 ( .A1(n13899), .A2(n13544), .B1(n676), .B2(n13541), .ZN(n8518) );
  OAI22_X1 U5693 ( .A1(n13905), .A2(n13544), .B1(n673), .B2(n13541), .ZN(n8519) );
  OAI22_X1 U5694 ( .A1(n13911), .A2(n13544), .B1(n670), .B2(n13541), .ZN(n8520) );
  OAI22_X1 U5695 ( .A1(n13917), .A2(n13544), .B1(n667), .B2(n13541), .ZN(n8521) );
  OAI22_X1 U5696 ( .A1(n13923), .A2(n13544), .B1(n664), .B2(n13541), .ZN(n8522) );
  OAI22_X1 U5697 ( .A1(n13929), .A2(n13544), .B1(n661), .B2(n13541), .ZN(n8523) );
  OAI22_X1 U5698 ( .A1(n13935), .A2(n13544), .B1(n658), .B2(n13541), .ZN(n8524) );
  OAI22_X1 U5699 ( .A1(n13941), .A2(n13544), .B1(n655), .B2(n13541), .ZN(n8525) );
  OAI22_X1 U5700 ( .A1(n13947), .A2(n13543), .B1(n652), .B2(n13541), .ZN(n8526) );
  OAI22_X1 U5701 ( .A1(n13953), .A2(n13543), .B1(n649), .B2(n13541), .ZN(n8527) );
  OAI22_X1 U5702 ( .A1(n13959), .A2(n13543), .B1(n646), .B2(n13541), .ZN(n8528) );
  OAI22_X1 U5703 ( .A1(n13965), .A2(n13543), .B1(n643), .B2(n13541), .ZN(n8529) );
  OAI22_X1 U5704 ( .A1(n13875), .A2(n13520), .B1(n992), .B2(n13516), .ZN(n8386) );
  OAI22_X1 U5705 ( .A1(n13881), .A2(n13520), .B1(n991), .B2(n13516), .ZN(n8387) );
  OAI22_X1 U5706 ( .A1(n13887), .A2(n13520), .B1(n990), .B2(n13516), .ZN(n8388) );
  OAI22_X1 U5707 ( .A1(n13893), .A2(n13520), .B1(n989), .B2(n13516), .ZN(n8389) );
  OAI22_X1 U5708 ( .A1(n13899), .A2(n13520), .B1(n988), .B2(n13517), .ZN(n8390) );
  OAI22_X1 U5709 ( .A1(n13905), .A2(n13520), .B1(n987), .B2(n13517), .ZN(n8391) );
  OAI22_X1 U5710 ( .A1(n13911), .A2(n13520), .B1(n986), .B2(n13517), .ZN(n8392) );
  OAI22_X1 U5711 ( .A1(n13917), .A2(n13520), .B1(n985), .B2(n13517), .ZN(n8393) );
  OAI22_X1 U5712 ( .A1(n13923), .A2(n13520), .B1(n984), .B2(n13517), .ZN(n8394) );
  OAI22_X1 U5713 ( .A1(n13929), .A2(n13520), .B1(n983), .B2(n13517), .ZN(n8395) );
  OAI22_X1 U5714 ( .A1(n13935), .A2(n13520), .B1(n982), .B2(n13517), .ZN(n8396) );
  OAI22_X1 U5715 ( .A1(n13941), .A2(n13520), .B1(n981), .B2(n13517), .ZN(n8397) );
  OAI22_X1 U5716 ( .A1(n13947), .A2(n13519), .B1(n980), .B2(n13517), .ZN(n8398) );
  OAI22_X1 U5717 ( .A1(n13953), .A2(n13519), .B1(n979), .B2(n13517), .ZN(n8399) );
  OAI22_X1 U5718 ( .A1(n13959), .A2(n13519), .B1(n978), .B2(n13517), .ZN(n8400) );
  OAI22_X1 U5719 ( .A1(n13965), .A2(n13519), .B1(n977), .B2(n13517), .ZN(n8401) );
  OAI22_X1 U5720 ( .A1(n13868), .A2(n13641), .B1(n5452), .B2(n13636), .ZN(
        n9025) );
  OAI22_X1 U5721 ( .A1(n13833), .A2(n13521), .B1(n999), .B2(n13516), .ZN(n8379) );
  OAI22_X1 U5722 ( .A1(n13839), .A2(n13521), .B1(n998), .B2(n13516), .ZN(n8380) );
  OAI22_X1 U5723 ( .A1(n13845), .A2(n13521), .B1(n997), .B2(n13516), .ZN(n8381) );
  OAI22_X1 U5724 ( .A1(n13851), .A2(n13521), .B1(n996), .B2(n13516), .ZN(n8382) );
  OAI22_X1 U5725 ( .A1(n13857), .A2(n13521), .B1(n995), .B2(n13516), .ZN(n8383) );
  OAI22_X1 U5726 ( .A1(n13863), .A2(n13521), .B1(n994), .B2(n13516), .ZN(n8384) );
  OAI22_X1 U5727 ( .A1(n13869), .A2(n13521), .B1(n993), .B2(n13516), .ZN(n8385) );
  OAI22_X1 U5728 ( .A1(n13828), .A2(n13437), .B1(n7192), .B2(n13432), .ZN(
        n7930) );
  OAI22_X1 U5729 ( .A1(n13828), .A2(n13467), .B1(n7224), .B2(n13462), .ZN(
        n8090) );
  OAI22_X1 U5730 ( .A1(n13834), .A2(n13467), .B1(n7225), .B2(n13462), .ZN(
        n8091) );
  OAI22_X1 U5731 ( .A1(n13840), .A2(n13467), .B1(n7226), .B2(n13462), .ZN(
        n8092) );
  OAI22_X1 U5732 ( .A1(n13846), .A2(n13467), .B1(n7227), .B2(n13462), .ZN(
        n8093) );
  OAI22_X1 U5733 ( .A1(n13852), .A2(n13467), .B1(n7228), .B2(n13462), .ZN(
        n8094) );
  OAI22_X1 U5734 ( .A1(n13858), .A2(n13467), .B1(n7229), .B2(n13462), .ZN(
        n8095) );
  OAI22_X1 U5735 ( .A1(n13864), .A2(n13467), .B1(n7230), .B2(n13462), .ZN(
        n8096) );
  OAI22_X1 U5736 ( .A1(n13870), .A2(n13467), .B1(n7231), .B2(n13462), .ZN(
        n8097) );
  OAI22_X1 U5737 ( .A1(n13876), .A2(n13466), .B1(n7232), .B2(n13462), .ZN(
        n8098) );
  OAI22_X1 U5738 ( .A1(n13882), .A2(n13466), .B1(n7233), .B2(n13462), .ZN(
        n8099) );
  OAI22_X1 U5739 ( .A1(n13888), .A2(n13466), .B1(n7234), .B2(n13462), .ZN(
        n8100) );
  OAI22_X1 U5740 ( .A1(n13894), .A2(n13466), .B1(n7235), .B2(n13462), .ZN(
        n8101) );
  OAI22_X1 U5741 ( .A1(n13900), .A2(n13466), .B1(n7236), .B2(n13463), .ZN(
        n8102) );
  OAI22_X1 U5742 ( .A1(n13906), .A2(n13466), .B1(n7237), .B2(n13463), .ZN(
        n8103) );
  OAI22_X1 U5743 ( .A1(n13912), .A2(n13466), .B1(n7238), .B2(n13463), .ZN(
        n8104) );
  OAI22_X1 U5744 ( .A1(n13918), .A2(n13466), .B1(n7239), .B2(n13463), .ZN(
        n8105) );
  OAI22_X1 U5745 ( .A1(n13924), .A2(n13466), .B1(n7240), .B2(n13463), .ZN(
        n8106) );
  OAI22_X1 U5746 ( .A1(n13930), .A2(n13466), .B1(n7241), .B2(n13463), .ZN(
        n8107) );
  OAI22_X1 U5747 ( .A1(n13936), .A2(n13466), .B1(n7242), .B2(n13463), .ZN(
        n8108) );
  OAI22_X1 U5748 ( .A1(n13942), .A2(n13466), .B1(n7243), .B2(n13463), .ZN(
        n8109) );
  OAI22_X1 U5749 ( .A1(n13948), .A2(n13465), .B1(n7244), .B2(n13463), .ZN(
        n8110) );
  OAI22_X1 U5750 ( .A1(n13954), .A2(n13465), .B1(n7245), .B2(n13463), .ZN(
        n8111) );
  OAI22_X1 U5751 ( .A1(n13960), .A2(n13465), .B1(n7246), .B2(n13463), .ZN(
        n8112) );
  OAI22_X1 U5752 ( .A1(n13966), .A2(n13465), .B1(n7247), .B2(n13463), .ZN(
        n8113) );
  OAI22_X1 U5753 ( .A1(n13827), .A2(n13515), .B1(n7022), .B2(n13510), .ZN(
        n8346) );
  OAI22_X1 U5754 ( .A1(n13834), .A2(n13515), .B1(n7023), .B2(n13510), .ZN(
        n8347) );
  OAI22_X1 U5755 ( .A1(n13840), .A2(n13515), .B1(n7024), .B2(n13510), .ZN(
        n8348) );
  OAI22_X1 U5756 ( .A1(n13846), .A2(n13515), .B1(n7025), .B2(n13510), .ZN(
        n8349) );
  OAI22_X1 U5757 ( .A1(n13852), .A2(n13515), .B1(n7026), .B2(n13510), .ZN(
        n8350) );
  OAI22_X1 U5758 ( .A1(n13858), .A2(n13515), .B1(n7027), .B2(n13510), .ZN(
        n8351) );
  OAI22_X1 U5759 ( .A1(n13864), .A2(n13515), .B1(n7028), .B2(n13510), .ZN(
        n8352) );
  OAI22_X1 U5760 ( .A1(n13870), .A2(n13515), .B1(n7029), .B2(n13510), .ZN(
        n8353) );
  OAI22_X1 U5761 ( .A1(n13876), .A2(n13514), .B1(n7030), .B2(n13510), .ZN(
        n8354) );
  OAI22_X1 U5762 ( .A1(n13882), .A2(n13514), .B1(n7031), .B2(n13510), .ZN(
        n8355) );
  OAI22_X1 U5763 ( .A1(n13888), .A2(n13514), .B1(n7032), .B2(n13510), .ZN(
        n8356) );
  OAI22_X1 U5764 ( .A1(n13894), .A2(n13514), .B1(n7033), .B2(n13510), .ZN(
        n8357) );
  OAI22_X1 U5765 ( .A1(n13900), .A2(n13514), .B1(n7034), .B2(n13511), .ZN(
        n8358) );
  OAI22_X1 U5766 ( .A1(n13906), .A2(n13514), .B1(n7035), .B2(n13511), .ZN(
        n8359) );
  OAI22_X1 U5767 ( .A1(n13912), .A2(n13514), .B1(n7036), .B2(n13511), .ZN(
        n8360) );
  OAI22_X1 U5768 ( .A1(n13918), .A2(n13514), .B1(n7037), .B2(n13511), .ZN(
        n8361) );
  OAI22_X1 U5769 ( .A1(n13924), .A2(n13514), .B1(n7038), .B2(n13511), .ZN(
        n8362) );
  OAI22_X1 U5770 ( .A1(n13930), .A2(n13514), .B1(n7039), .B2(n13511), .ZN(
        n8363) );
  OAI22_X1 U5771 ( .A1(n13936), .A2(n13514), .B1(n7040), .B2(n13511), .ZN(
        n8364) );
  OAI22_X1 U5772 ( .A1(n13942), .A2(n13514), .B1(n7041), .B2(n13511), .ZN(
        n8365) );
  OAI22_X1 U5773 ( .A1(n13948), .A2(n13513), .B1(n7042), .B2(n13511), .ZN(
        n8366) );
  OAI22_X1 U5774 ( .A1(n13954), .A2(n13513), .B1(n7043), .B2(n13511), .ZN(
        n8367) );
  OAI22_X1 U5775 ( .A1(n13960), .A2(n13513), .B1(n7044), .B2(n13511), .ZN(
        n8368) );
  OAI22_X1 U5776 ( .A1(n13966), .A2(n13513), .B1(n7045), .B2(n13511), .ZN(
        n8369) );
  OAI22_X1 U5777 ( .A1(n13827), .A2(n13521), .B1(n7256), .B2(n13516), .ZN(
        n8378) );
  OAI22_X1 U5778 ( .A1(n13826), .A2(n13623), .B1(n7046), .B2(n13618), .ZN(
        n8922) );
  OAI22_X1 U5779 ( .A1(n13832), .A2(n13623), .B1(n7047), .B2(n13618), .ZN(
        n8923) );
  OAI22_X1 U5780 ( .A1(n13838), .A2(n13623), .B1(n7048), .B2(n13618), .ZN(
        n8924) );
  OAI22_X1 U5781 ( .A1(n13844), .A2(n13623), .B1(n7049), .B2(n13618), .ZN(
        n8925) );
  OAI22_X1 U5782 ( .A1(n13850), .A2(n13623), .B1(n7050), .B2(n13618), .ZN(
        n8926) );
  OAI22_X1 U5783 ( .A1(n13856), .A2(n13623), .B1(n7051), .B2(n13618), .ZN(
        n8927) );
  OAI22_X1 U5784 ( .A1(n13862), .A2(n13623), .B1(n7052), .B2(n13618), .ZN(
        n8928) );
  OAI22_X1 U5785 ( .A1(n13868), .A2(n13623), .B1(n7053), .B2(n13618), .ZN(
        n8929) );
  OAI22_X1 U5786 ( .A1(n13874), .A2(n13622), .B1(n7054), .B2(n13618), .ZN(
        n8930) );
  OAI22_X1 U5787 ( .A1(n13880), .A2(n13622), .B1(n7055), .B2(n13618), .ZN(
        n8931) );
  OAI22_X1 U5788 ( .A1(n13886), .A2(n13622), .B1(n7056), .B2(n13618), .ZN(
        n8932) );
  OAI22_X1 U5789 ( .A1(n13892), .A2(n13622), .B1(n7057), .B2(n13618), .ZN(
        n8933) );
  OAI22_X1 U5790 ( .A1(n13898), .A2(n13622), .B1(n7058), .B2(n13619), .ZN(
        n8934) );
  OAI22_X1 U5791 ( .A1(n13904), .A2(n13622), .B1(n7059), .B2(n13619), .ZN(
        n8935) );
  OAI22_X1 U5792 ( .A1(n13910), .A2(n13622), .B1(n7060), .B2(n13619), .ZN(
        n8936) );
  OAI22_X1 U5793 ( .A1(n13916), .A2(n13622), .B1(n7061), .B2(n13619), .ZN(
        n8937) );
  OAI22_X1 U5794 ( .A1(n13922), .A2(n13622), .B1(n7062), .B2(n13619), .ZN(
        n8938) );
  OAI22_X1 U5795 ( .A1(n13928), .A2(n13622), .B1(n7063), .B2(n13619), .ZN(
        n8939) );
  OAI22_X1 U5796 ( .A1(n13934), .A2(n13622), .B1(n7064), .B2(n13619), .ZN(
        n8940) );
  OAI22_X1 U5797 ( .A1(n13940), .A2(n13622), .B1(n7065), .B2(n13619), .ZN(
        n8941) );
  OAI22_X1 U5798 ( .A1(n13946), .A2(n13621), .B1(n7066), .B2(n13619), .ZN(
        n8942) );
  OAI22_X1 U5799 ( .A1(n13952), .A2(n13621), .B1(n7067), .B2(n13619), .ZN(
        n8943) );
  OAI22_X1 U5800 ( .A1(n13958), .A2(n13621), .B1(n7068), .B2(n13619), .ZN(
        n8944) );
  OAI22_X1 U5801 ( .A1(n13964), .A2(n13621), .B1(n7069), .B2(n13619), .ZN(
        n8945) );
  OAI22_X1 U5802 ( .A1(n13826), .A2(n13641), .B1(n7153), .B2(n13636), .ZN(
        n9018) );
  OAI22_X1 U5803 ( .A1(n13832), .A2(n13641), .B1(n7154), .B2(n13636), .ZN(
        n9019) );
  OAI22_X1 U5804 ( .A1(n13838), .A2(n13641), .B1(n7155), .B2(n13636), .ZN(
        n9020) );
  OAI22_X1 U5805 ( .A1(n13844), .A2(n13641), .B1(n7156), .B2(n13636), .ZN(
        n9021) );
  OAI22_X1 U5806 ( .A1(n13850), .A2(n13641), .B1(n7157), .B2(n13636), .ZN(
        n9022) );
  OAI22_X1 U5807 ( .A1(n13856), .A2(n13641), .B1(n7158), .B2(n13636), .ZN(
        n9023) );
  OAI22_X1 U5808 ( .A1(n13862), .A2(n13641), .B1(n7159), .B2(n13636), .ZN(
        n9024) );
  OAI22_X1 U5809 ( .A1(n13825), .A2(n13677), .B1(n7070), .B2(n13672), .ZN(
        n9210) );
  OAI22_X1 U5810 ( .A1(n13831), .A2(n13677), .B1(n7071), .B2(n13672), .ZN(
        n9211) );
  OAI22_X1 U5811 ( .A1(n13837), .A2(n13677), .B1(n7072), .B2(n13672), .ZN(
        n9212) );
  OAI22_X1 U5812 ( .A1(n13843), .A2(n13677), .B1(n7073), .B2(n13672), .ZN(
        n9213) );
  OAI22_X1 U5813 ( .A1(n13849), .A2(n13677), .B1(n7074), .B2(n13672), .ZN(
        n9214) );
  OAI22_X1 U5814 ( .A1(n13855), .A2(n13677), .B1(n7075), .B2(n13672), .ZN(
        n9215) );
  OAI22_X1 U5815 ( .A1(n13861), .A2(n13677), .B1(n7076), .B2(n13672), .ZN(
        n9216) );
  OAI22_X1 U5816 ( .A1(n13867), .A2(n13677), .B1(n7077), .B2(n13672), .ZN(
        n9217) );
  OAI22_X1 U5817 ( .A1(n13873), .A2(n13676), .B1(n7078), .B2(n13672), .ZN(
        n9218) );
  OAI22_X1 U5818 ( .A1(n13879), .A2(n13676), .B1(n7079), .B2(n13672), .ZN(
        n9219) );
  OAI22_X1 U5819 ( .A1(n13885), .A2(n13676), .B1(n7080), .B2(n13672), .ZN(
        n9220) );
  OAI22_X1 U5820 ( .A1(n13891), .A2(n13676), .B1(n7081), .B2(n13672), .ZN(
        n9221) );
  OAI22_X1 U5821 ( .A1(n13897), .A2(n13676), .B1(n7082), .B2(n13673), .ZN(
        n9222) );
  OAI22_X1 U5822 ( .A1(n13903), .A2(n13676), .B1(n7083), .B2(n13673), .ZN(
        n9223) );
  OAI22_X1 U5823 ( .A1(n13909), .A2(n13676), .B1(n7084), .B2(n13673), .ZN(
        n9224) );
  OAI22_X1 U5824 ( .A1(n13915), .A2(n13676), .B1(n7085), .B2(n13673), .ZN(
        n9225) );
  OAI22_X1 U5825 ( .A1(n13921), .A2(n13676), .B1(n7086), .B2(n13673), .ZN(
        n9226) );
  OAI22_X1 U5826 ( .A1(n13927), .A2(n13676), .B1(n7087), .B2(n13673), .ZN(
        n9227) );
  OAI22_X1 U5827 ( .A1(n13933), .A2(n13676), .B1(n7088), .B2(n13673), .ZN(
        n9228) );
  OAI22_X1 U5828 ( .A1(n13939), .A2(n13676), .B1(n7089), .B2(n13673), .ZN(
        n9229) );
  OAI22_X1 U5829 ( .A1(n13945), .A2(n13675), .B1(n7090), .B2(n13673), .ZN(
        n9230) );
  OAI22_X1 U5830 ( .A1(n13951), .A2(n13675), .B1(n7091), .B2(n13673), .ZN(
        n9231) );
  OAI22_X1 U5831 ( .A1(n13957), .A2(n13675), .B1(n7092), .B2(n13673), .ZN(
        n9232) );
  OAI22_X1 U5832 ( .A1(n13963), .A2(n13675), .B1(n7093), .B2(n13673), .ZN(
        n9233) );
  OAI22_X1 U5833 ( .A1(n13825), .A2(n13695), .B1(n6998), .B2(n13690), .ZN(
        n9306) );
  OAI22_X1 U5834 ( .A1(n13831), .A2(n13695), .B1(n6999), .B2(n13690), .ZN(
        n9307) );
  OAI22_X1 U5835 ( .A1(n13837), .A2(n13695), .B1(n7000), .B2(n13690), .ZN(
        n9308) );
  OAI22_X1 U5836 ( .A1(n13843), .A2(n13695), .B1(n7001), .B2(n13690), .ZN(
        n9309) );
  OAI22_X1 U5837 ( .A1(n13849), .A2(n13695), .B1(n7002), .B2(n13690), .ZN(
        n9310) );
  OAI22_X1 U5838 ( .A1(n13855), .A2(n13695), .B1(n7003), .B2(n13690), .ZN(
        n9311) );
  OAI22_X1 U5839 ( .A1(n13861), .A2(n13695), .B1(n7004), .B2(n13690), .ZN(
        n9312) );
  OAI22_X1 U5840 ( .A1(n13867), .A2(n13695), .B1(n7005), .B2(n13690), .ZN(
        n9313) );
  OAI22_X1 U5841 ( .A1(n13873), .A2(n13694), .B1(n7094), .B2(n13690), .ZN(
        n9314) );
  OAI22_X1 U5842 ( .A1(n13879), .A2(n13694), .B1(n7095), .B2(n13690), .ZN(
        n9315) );
  OAI22_X1 U5843 ( .A1(n13885), .A2(n13694), .B1(n7096), .B2(n13690), .ZN(
        n9316) );
  OAI22_X1 U5844 ( .A1(n13891), .A2(n13694), .B1(n7097), .B2(n13690), .ZN(
        n9317) );
  OAI22_X1 U5845 ( .A1(n13897), .A2(n13694), .B1(n7098), .B2(n13691), .ZN(
        n9318) );
  OAI22_X1 U5846 ( .A1(n13903), .A2(n13694), .B1(n7099), .B2(n13691), .ZN(
        n9319) );
  OAI22_X1 U5847 ( .A1(n13909), .A2(n13694), .B1(n7100), .B2(n13691), .ZN(
        n9320) );
  OAI22_X1 U5848 ( .A1(n13915), .A2(n13694), .B1(n7101), .B2(n13691), .ZN(
        n9321) );
  OAI22_X1 U5849 ( .A1(n13921), .A2(n13694), .B1(n7102), .B2(n13691), .ZN(
        n9322) );
  OAI22_X1 U5850 ( .A1(n13927), .A2(n13694), .B1(n7103), .B2(n13691), .ZN(
        n9323) );
  OAI22_X1 U5851 ( .A1(n13933), .A2(n13694), .B1(n7104), .B2(n13691), .ZN(
        n9324) );
  OAI22_X1 U5852 ( .A1(n13825), .A2(n13731), .B1(n7105), .B2(n13726), .ZN(
        n9498) );
  OAI22_X1 U5853 ( .A1(n13831), .A2(n13731), .B1(n7106), .B2(n13726), .ZN(
        n9499) );
  OAI22_X1 U5854 ( .A1(n13837), .A2(n13731), .B1(n7107), .B2(n13726), .ZN(
        n9500) );
  OAI22_X1 U5855 ( .A1(n13843), .A2(n13731), .B1(n7108), .B2(n13726), .ZN(
        n9501) );
  OAI22_X1 U5856 ( .A1(n13849), .A2(n13731), .B1(n7109), .B2(n13726), .ZN(
        n9502) );
  OAI22_X1 U5857 ( .A1(n13855), .A2(n13731), .B1(n7110), .B2(n13726), .ZN(
        n9503) );
  OAI22_X1 U5858 ( .A1(n13861), .A2(n13731), .B1(n7111), .B2(n13726), .ZN(
        n9504) );
  OAI22_X1 U5859 ( .A1(n13867), .A2(n13731), .B1(n7112), .B2(n13726), .ZN(
        n9505) );
  OAI22_X1 U5860 ( .A1(n13873), .A2(n13730), .B1(n7113), .B2(n13726), .ZN(
        n9506) );
  OAI22_X1 U5861 ( .A1(n13879), .A2(n13730), .B1(n7114), .B2(n13726), .ZN(
        n9507) );
  OAI22_X1 U5862 ( .A1(n13885), .A2(n13730), .B1(n7115), .B2(n13726), .ZN(
        n9508) );
  OAI22_X1 U5863 ( .A1(n13891), .A2(n13730), .B1(n7116), .B2(n13726), .ZN(
        n9509) );
  OAI22_X1 U5864 ( .A1(n13897), .A2(n13730), .B1(n7117), .B2(n13727), .ZN(
        n9510) );
  OAI22_X1 U5865 ( .A1(n13903), .A2(n13730), .B1(n7118), .B2(n13727), .ZN(
        n9511) );
  OAI22_X1 U5866 ( .A1(n13909), .A2(n13730), .B1(n7119), .B2(n13727), .ZN(
        n9512) );
  OAI22_X1 U5867 ( .A1(n13915), .A2(n13730), .B1(n7120), .B2(n13727), .ZN(
        n9513) );
  OAI22_X1 U5868 ( .A1(n13921), .A2(n13730), .B1(n7121), .B2(n13727), .ZN(
        n9514) );
  OAI22_X1 U5869 ( .A1(n13927), .A2(n13730), .B1(n7122), .B2(n13727), .ZN(
        n9515) );
  OAI22_X1 U5870 ( .A1(n13933), .A2(n13730), .B1(n7123), .B2(n13727), .ZN(
        n9516) );
  OAI22_X1 U5871 ( .A1(n13939), .A2(n13730), .B1(n7124), .B2(n13727), .ZN(
        n9517) );
  OAI22_X1 U5872 ( .A1(n13945), .A2(n13729), .B1(n7125), .B2(n13727), .ZN(
        n9518) );
  OAI22_X1 U5873 ( .A1(n13951), .A2(n13729), .B1(n7126), .B2(n13727), .ZN(
        n9519) );
  OAI22_X1 U5874 ( .A1(n13957), .A2(n13729), .B1(n7127), .B2(n13727), .ZN(
        n9520) );
  OAI22_X1 U5875 ( .A1(n13963), .A2(n13729), .B1(n7128), .B2(n13727), .ZN(
        n9521) );
  OAI22_X1 U5876 ( .A1(n13824), .A2(n13785), .B1(n7129), .B2(n13780), .ZN(
        n9786) );
  OAI22_X1 U5877 ( .A1(n13830), .A2(n13785), .B1(n7130), .B2(n13780), .ZN(
        n9787) );
  OAI22_X1 U5878 ( .A1(n13836), .A2(n13785), .B1(n7131), .B2(n13780), .ZN(
        n9788) );
  OAI22_X1 U5879 ( .A1(n13842), .A2(n13785), .B1(n7132), .B2(n13780), .ZN(
        n9789) );
  OAI22_X1 U5880 ( .A1(n13848), .A2(n13785), .B1(n7133), .B2(n13780), .ZN(
        n9790) );
  OAI22_X1 U5881 ( .A1(n13854), .A2(n13785), .B1(n7134), .B2(n13780), .ZN(
        n9791) );
  OAI22_X1 U5882 ( .A1(n13860), .A2(n13785), .B1(n7135), .B2(n13780), .ZN(
        n9792) );
  OAI22_X1 U5883 ( .A1(n13866), .A2(n13785), .B1(n7136), .B2(n13780), .ZN(
        n9793) );
  OAI22_X1 U5884 ( .A1(n13872), .A2(n13784), .B1(n7137), .B2(n13780), .ZN(
        n9794) );
  OAI22_X1 U5885 ( .A1(n13878), .A2(n13784), .B1(n7138), .B2(n13780), .ZN(
        n9795) );
  OAI22_X1 U5886 ( .A1(n13884), .A2(n13784), .B1(n7139), .B2(n13780), .ZN(
        n9796) );
  OAI22_X1 U5887 ( .A1(n13890), .A2(n13784), .B1(n7140), .B2(n13780), .ZN(
        n9797) );
  OAI22_X1 U5888 ( .A1(n13896), .A2(n13784), .B1(n7141), .B2(n13781), .ZN(
        n9798) );
  OAI22_X1 U5889 ( .A1(n13902), .A2(n13784), .B1(n7142), .B2(n13781), .ZN(
        n9799) );
  OAI22_X1 U5890 ( .A1(n13908), .A2(n13784), .B1(n7143), .B2(n13781), .ZN(
        n9800) );
  OAI22_X1 U5891 ( .A1(n13914), .A2(n13784), .B1(n7144), .B2(n13781), .ZN(
        n9801) );
  OAI22_X1 U5892 ( .A1(n13920), .A2(n13784), .B1(n7145), .B2(n13781), .ZN(
        n9802) );
  OAI22_X1 U5893 ( .A1(n13926), .A2(n13784), .B1(n7146), .B2(n13781), .ZN(
        n9803) );
  OAI22_X1 U5894 ( .A1(n13932), .A2(n13784), .B1(n7147), .B2(n13781), .ZN(
        n9804) );
  OAI22_X1 U5895 ( .A1(n13938), .A2(n13784), .B1(n7148), .B2(n13781), .ZN(
        n9805) );
  OAI22_X1 U5896 ( .A1(n13944), .A2(n13783), .B1(n7149), .B2(n13781), .ZN(
        n9806) );
  OAI22_X1 U5897 ( .A1(n13950), .A2(n13783), .B1(n7150), .B2(n13781), .ZN(
        n9807) );
  OAI22_X1 U5898 ( .A1(n13956), .A2(n13783), .B1(n7151), .B2(n13781), .ZN(
        n9808) );
  OAI22_X1 U5899 ( .A1(n13962), .A2(n13783), .B1(n7152), .B2(n13781), .ZN(
        n9809) );
  OAI22_X1 U5900 ( .A1(n13828), .A2(n13473), .B1(n13468), .B2(n12726), .ZN(
        n8122) );
  OAI22_X1 U5901 ( .A1(n13834), .A2(n13473), .B1(n13468), .B2(n12727), .ZN(
        n8123) );
  OAI22_X1 U5902 ( .A1(n13840), .A2(n13473), .B1(n13468), .B2(n12728), .ZN(
        n8124) );
  OAI22_X1 U5903 ( .A1(n13846), .A2(n13473), .B1(n13468), .B2(n12729), .ZN(
        n8125) );
  OAI22_X1 U5904 ( .A1(n13852), .A2(n13473), .B1(n13468), .B2(n12730), .ZN(
        n8126) );
  OAI22_X1 U5905 ( .A1(n13858), .A2(n13473), .B1(n13468), .B2(n12731), .ZN(
        n8127) );
  OAI22_X1 U5906 ( .A1(n13864), .A2(n13473), .B1(n13468), .B2(n12732), .ZN(
        n8128) );
  OAI22_X1 U5907 ( .A1(n13870), .A2(n13473), .B1(n13468), .B2(n12733), .ZN(
        n8129) );
  OAI22_X1 U5908 ( .A1(n13876), .A2(n13472), .B1(n13468), .B2(n12734), .ZN(
        n8130) );
  OAI22_X1 U5909 ( .A1(n13882), .A2(n13472), .B1(n13468), .B2(n12735), .ZN(
        n8131) );
  OAI22_X1 U5910 ( .A1(n13888), .A2(n13472), .B1(n13468), .B2(n12736), .ZN(
        n8132) );
  OAI22_X1 U5911 ( .A1(n13894), .A2(n13472), .B1(n13468), .B2(n12737), .ZN(
        n8133) );
  OAI22_X1 U5912 ( .A1(n13900), .A2(n13472), .B1(n13469), .B2(n12738), .ZN(
        n8134) );
  OAI22_X1 U5913 ( .A1(n13906), .A2(n13472), .B1(n13469), .B2(n12739), .ZN(
        n8135) );
  OAI22_X1 U5914 ( .A1(n13912), .A2(n13472), .B1(n13469), .B2(n12740), .ZN(
        n8136) );
  OAI22_X1 U5915 ( .A1(n13918), .A2(n13472), .B1(n13469), .B2(n12741), .ZN(
        n8137) );
  OAI22_X1 U5916 ( .A1(n13924), .A2(n13472), .B1(n13469), .B2(n12742), .ZN(
        n8138) );
  OAI22_X1 U5917 ( .A1(n13930), .A2(n13472), .B1(n13469), .B2(n12743), .ZN(
        n8139) );
  OAI22_X1 U5918 ( .A1(n13936), .A2(n13472), .B1(n13469), .B2(n12744), .ZN(
        n8140) );
  OAI22_X1 U5919 ( .A1(n13942), .A2(n13472), .B1(n13469), .B2(n12745), .ZN(
        n8141) );
  OAI22_X1 U5920 ( .A1(n13948), .A2(n13471), .B1(n13469), .B2(n12746), .ZN(
        n8142) );
  OAI22_X1 U5921 ( .A1(n13954), .A2(n13471), .B1(n13469), .B2(n12747), .ZN(
        n8143) );
  OAI22_X1 U5922 ( .A1(n13960), .A2(n13471), .B1(n13469), .B2(n12748), .ZN(
        n8144) );
  OAI22_X1 U5923 ( .A1(n13966), .A2(n13471), .B1(n13469), .B2(n12749), .ZN(
        n8145) );
  OAI22_X1 U5924 ( .A1(n13828), .A2(n13479), .B1(n13474), .B2(n12750), .ZN(
        n8154) );
  OAI22_X1 U5925 ( .A1(n13834), .A2(n13479), .B1(n13474), .B2(n12751), .ZN(
        n8155) );
  OAI22_X1 U5926 ( .A1(n13840), .A2(n13479), .B1(n13474), .B2(n12752), .ZN(
        n8156) );
  OAI22_X1 U5927 ( .A1(n13846), .A2(n13479), .B1(n13474), .B2(n12753), .ZN(
        n8157) );
  OAI22_X1 U5928 ( .A1(n13852), .A2(n13479), .B1(n13474), .B2(n12754), .ZN(
        n8158) );
  OAI22_X1 U5929 ( .A1(n13858), .A2(n13479), .B1(n13474), .B2(n12755), .ZN(
        n8159) );
  OAI22_X1 U5930 ( .A1(n13864), .A2(n13479), .B1(n13474), .B2(n12756), .ZN(
        n8160) );
  OAI22_X1 U5931 ( .A1(n13870), .A2(n13479), .B1(n13474), .B2(n12757), .ZN(
        n8161) );
  OAI22_X1 U5932 ( .A1(n13876), .A2(n13478), .B1(n13474), .B2(n12758), .ZN(
        n8162) );
  OAI22_X1 U5933 ( .A1(n13882), .A2(n13478), .B1(n13474), .B2(n12759), .ZN(
        n8163) );
  OAI22_X1 U5934 ( .A1(n13888), .A2(n13478), .B1(n13474), .B2(n12760), .ZN(
        n8164) );
  OAI22_X1 U5935 ( .A1(n13894), .A2(n13478), .B1(n13474), .B2(n12761), .ZN(
        n8165) );
  OAI22_X1 U5936 ( .A1(n13900), .A2(n13478), .B1(n13475), .B2(n12762), .ZN(
        n8166) );
  OAI22_X1 U5937 ( .A1(n13906), .A2(n13478), .B1(n13475), .B2(n12763), .ZN(
        n8167) );
  OAI22_X1 U5938 ( .A1(n13912), .A2(n13478), .B1(n13475), .B2(n12764), .ZN(
        n8168) );
  OAI22_X1 U5939 ( .A1(n13918), .A2(n13478), .B1(n13475), .B2(n12765), .ZN(
        n8169) );
  OAI22_X1 U5940 ( .A1(n13924), .A2(n13478), .B1(n13475), .B2(n12766), .ZN(
        n8170) );
  OAI22_X1 U5941 ( .A1(n13930), .A2(n13478), .B1(n13475), .B2(n12767), .ZN(
        n8171) );
  OAI22_X1 U5942 ( .A1(n13936), .A2(n13478), .B1(n13475), .B2(n12768), .ZN(
        n8172) );
  OAI22_X1 U5943 ( .A1(n13942), .A2(n13478), .B1(n13475), .B2(n12769), .ZN(
        n8173) );
  OAI22_X1 U5944 ( .A1(n13948), .A2(n13477), .B1(n13475), .B2(n12770), .ZN(
        n8174) );
  OAI22_X1 U5945 ( .A1(n13954), .A2(n13477), .B1(n13475), .B2(n12771), .ZN(
        n8175) );
  OAI22_X1 U5946 ( .A1(n13960), .A2(n13477), .B1(n13475), .B2(n12772), .ZN(
        n8176) );
  OAI22_X1 U5947 ( .A1(n13966), .A2(n13477), .B1(n13475), .B2(n12773), .ZN(
        n8177) );
  NAND4_X1 U5948 ( .A1(n4624), .A2(n4625), .A3(n4626), .A4(n4627), .ZN(n4623)
         );
  AOI221_X1 U5949 ( .B1(n13101), .B2(n732), .C1(n13098), .C2(n15945), .A(n4631), .ZN(n4624) );
  AOI221_X1 U5950 ( .B1(n13128), .B2(n731), .C1(n13125), .C2(n15937), .A(n4629), .ZN(n4626) );
  AOI221_X1 U5951 ( .B1(n13116), .B2(n14082), .C1(n13113), .C2(n15604), .A(
        n4630), .ZN(n4625) );
  NAND4_X1 U5952 ( .A1(n4587), .A2(n4588), .A3(n4589), .A4(n4590), .ZN(n4586)
         );
  AOI221_X1 U5953 ( .B1(n13101), .B2(n729), .C1(n13098), .C2(n15944), .A(n4594), .ZN(n4587) );
  AOI221_X1 U5954 ( .B1(n13128), .B2(n728), .C1(n13125), .C2(n15936), .A(n4592), .ZN(n4589) );
  AOI221_X1 U5955 ( .B1(n13116), .B2(n14081), .C1(n13113), .C2(n15603), .A(
        n4593), .ZN(n4588) );
  NAND4_X1 U5956 ( .A1(n4550), .A2(n4551), .A3(n4552), .A4(n4553), .ZN(n4549)
         );
  AOI221_X1 U5957 ( .B1(n13101), .B2(n726), .C1(n13098), .C2(n15943), .A(n4557), .ZN(n4550) );
  AOI221_X1 U5958 ( .B1(n13128), .B2(n725), .C1(n13125), .C2(n15935), .A(n4555), .ZN(n4552) );
  AOI221_X1 U5959 ( .B1(n13116), .B2(n14080), .C1(n13113), .C2(n15602), .A(
        n4556), .ZN(n4551) );
  NAND4_X1 U5960 ( .A1(n4513), .A2(n4514), .A3(n4515), .A4(n4516), .ZN(n4512)
         );
  AOI221_X1 U5961 ( .B1(n13101), .B2(n723), .C1(n13098), .C2(n15942), .A(n4520), .ZN(n4513) );
  AOI221_X1 U5962 ( .B1(n13128), .B2(n722), .C1(n13125), .C2(n15934), .A(n4518), .ZN(n4515) );
  AOI221_X1 U5963 ( .B1(n13116), .B2(n14079), .C1(n13113), .C2(n15601), .A(
        n4519), .ZN(n4514) );
  NAND4_X1 U5964 ( .A1(n4476), .A2(n4477), .A3(n4478), .A4(n4479), .ZN(n4475)
         );
  AOI221_X1 U5965 ( .B1(n13101), .B2(n720), .C1(n13098), .C2(n15941), .A(n4483), .ZN(n4476) );
  AOI221_X1 U5966 ( .B1(n13128), .B2(n719), .C1(n13125), .C2(n15933), .A(n4481), .ZN(n4478) );
  AOI221_X1 U5967 ( .B1(n13116), .B2(n14078), .C1(n13113), .C2(n15600), .A(
        n4482), .ZN(n4477) );
  NAND4_X1 U5968 ( .A1(n4439), .A2(n4440), .A3(n4441), .A4(n4442), .ZN(n4438)
         );
  AOI221_X1 U5969 ( .B1(n13101), .B2(n717), .C1(n13098), .C2(n15940), .A(n4446), .ZN(n4439) );
  AOI221_X1 U5970 ( .B1(n13128), .B2(n716), .C1(n13125), .C2(n15932), .A(n4444), .ZN(n4441) );
  AOI221_X1 U5971 ( .B1(n13116), .B2(n14077), .C1(n13113), .C2(n15599), .A(
        n4445), .ZN(n4440) );
  NAND4_X1 U5972 ( .A1(n4330), .A2(n4331), .A3(n4332), .A4(n4333), .ZN(n4329)
         );
  AOI221_X1 U5973 ( .B1(n13101), .B2(n714), .C1(n13098), .C2(n15939), .A(n4353), .ZN(n4330) );
  AOI221_X1 U5974 ( .B1(n13128), .B2(n713), .C1(n13125), .C2(n15931), .A(n4342), .ZN(n4332) );
  AOI221_X1 U5975 ( .B1(n13116), .B2(n14076), .C1(n13113), .C2(n15598), .A(
        n4347), .ZN(n4331) );
  NAND4_X1 U5976 ( .A1(n5650), .A2(n5651), .A3(n5654), .A4(n5656), .ZN(n5649)
         );
  AOI221_X1 U5977 ( .B1(n13099), .B2(n807), .C1(n13096), .C2(n16030), .A(n5680), .ZN(n5650) );
  AOI221_X1 U5978 ( .B1(n13126), .B2(n806), .C1(n13123), .C2(n15994), .A(n5670), .ZN(n5654) );
  AOI221_X1 U5979 ( .B1(n13114), .B2(n14107), .C1(n13111), .C2(n15921), .A(
        n5678), .ZN(n5651) );
  NAND4_X1 U5980 ( .A1(n5589), .A2(n5590), .A3(n5591), .A4(n5594), .ZN(n5588)
         );
  AOI221_X1 U5981 ( .B1(n13099), .B2(n804), .C1(n13096), .C2(n16029), .A(n5600), .ZN(n5589) );
  AOI221_X1 U5982 ( .B1(n13126), .B2(n803), .C1(n13123), .C2(n15993), .A(n5598), .ZN(n5591) );
  AOI221_X1 U5983 ( .B1(n13114), .B2(n14106), .C1(n13111), .C2(n15920), .A(
        n5599), .ZN(n5590) );
  NAND4_X1 U5984 ( .A1(n5528), .A2(n5529), .A3(n5530), .A4(n5531), .ZN(n5526)
         );
  AOI221_X1 U5985 ( .B1(n13099), .B2(n801), .C1(n13096), .C2(n16028), .A(n5539), .ZN(n5528) );
  AOI221_X1 U5986 ( .B1(n13126), .B2(n800), .C1(n13123), .C2(n15992), .A(n5536), .ZN(n5530) );
  AOI221_X1 U5987 ( .B1(n13114), .B2(n14105), .C1(n13111), .C2(n15919), .A(
        n5538), .ZN(n5529) );
  NAND4_X1 U5988 ( .A1(n5466), .A2(n5468), .A3(n5469), .A4(n5470), .ZN(n5464)
         );
  AOI221_X1 U5989 ( .B1(n13099), .B2(n798), .C1(n13096), .C2(n16027), .A(n5478), .ZN(n5466) );
  AOI221_X1 U5990 ( .B1(n13126), .B2(n797), .C1(n13123), .C2(n15991), .A(n5474), .ZN(n5469) );
  AOI221_X1 U5991 ( .B1(n13114), .B2(n14104), .C1(n13111), .C2(n15918), .A(
        n5476), .ZN(n5468) );
  NAND4_X1 U5992 ( .A1(n5410), .A2(n5411), .A3(n5412), .A4(n5414), .ZN(n5409)
         );
  AOI221_X1 U5993 ( .B1(n13099), .B2(n795), .C1(n13096), .C2(n16026), .A(n5420), .ZN(n5410) );
  AOI221_X1 U5994 ( .B1(n13126), .B2(n794), .C1(n13123), .C2(n15990), .A(n5418), .ZN(n5412) );
  AOI221_X1 U5995 ( .B1(n13114), .B2(n14103), .C1(n13111), .C2(n15917), .A(
        n5419), .ZN(n5411) );
  NAND4_X1 U5996 ( .A1(n5364), .A2(n5365), .A3(n5366), .A4(n5367), .ZN(n5363)
         );
  AOI221_X1 U5997 ( .B1(n13099), .B2(n792), .C1(n13096), .C2(n16025), .A(n5371), .ZN(n5364) );
  AOI221_X1 U5998 ( .B1(n13126), .B2(n791), .C1(n13123), .C2(n15989), .A(n5369), .ZN(n5366) );
  AOI221_X1 U5999 ( .B1(n13114), .B2(n14102), .C1(n13111), .C2(n15916), .A(
        n5370), .ZN(n5365) );
  NAND4_X1 U6000 ( .A1(n5327), .A2(n5328), .A3(n5329), .A4(n5330), .ZN(n5326)
         );
  AOI221_X1 U6001 ( .B1(n13099), .B2(n789), .C1(n13096), .C2(n16024), .A(n5334), .ZN(n5327) );
  AOI221_X1 U6002 ( .B1(n13126), .B2(n788), .C1(n13123), .C2(n15988), .A(n5332), .ZN(n5329) );
  AOI221_X1 U6003 ( .B1(n13114), .B2(n14101), .C1(n13111), .C2(n15915), .A(
        n5333), .ZN(n5328) );
  NAND4_X1 U6004 ( .A1(n5290), .A2(n5291), .A3(n5292), .A4(n5293), .ZN(n5289)
         );
  AOI221_X1 U6005 ( .B1(n13099), .B2(n786), .C1(n13096), .C2(n16023), .A(n5297), .ZN(n5290) );
  AOI221_X1 U6006 ( .B1(n13126), .B2(n785), .C1(n13123), .C2(n15987), .A(n5295), .ZN(n5292) );
  AOI221_X1 U6007 ( .B1(n13114), .B2(n14100), .C1(n13111), .C2(n15914), .A(
        n5296), .ZN(n5291) );
  NAND4_X1 U6008 ( .A1(n5253), .A2(n5254), .A3(n5255), .A4(n5256), .ZN(n5252)
         );
  AOI221_X1 U6009 ( .B1(n13099), .B2(n783), .C1(n13096), .C2(n16022), .A(n5260), .ZN(n5253) );
  AOI221_X1 U6010 ( .B1(n13126), .B2(n782), .C1(n13123), .C2(n15986), .A(n5258), .ZN(n5255) );
  AOI221_X1 U6011 ( .B1(n13114), .B2(n14099), .C1(n13111), .C2(n15913), .A(
        n5259), .ZN(n5254) );
  NAND4_X1 U6012 ( .A1(n5216), .A2(n5217), .A3(n5218), .A4(n5219), .ZN(n5215)
         );
  AOI221_X1 U6013 ( .B1(n13099), .B2(n780), .C1(n13096), .C2(n16021), .A(n5223), .ZN(n5216) );
  AOI221_X1 U6014 ( .B1(n13126), .B2(n779), .C1(n13123), .C2(n15985), .A(n5221), .ZN(n5218) );
  AOI221_X1 U6015 ( .B1(n13114), .B2(n14098), .C1(n13111), .C2(n15912), .A(
        n5222), .ZN(n5217) );
  NAND4_X1 U6016 ( .A1(n5179), .A2(n5180), .A3(n5181), .A4(n5182), .ZN(n5178)
         );
  AOI221_X1 U6017 ( .B1(n13099), .B2(n777), .C1(n13096), .C2(n16020), .A(n5186), .ZN(n5179) );
  AOI221_X1 U6018 ( .B1(n13126), .B2(n776), .C1(n13123), .C2(n15984), .A(n5184), .ZN(n5181) );
  AOI221_X1 U6019 ( .B1(n13114), .B2(n14097), .C1(n13111), .C2(n15911), .A(
        n5185), .ZN(n5180) );
  NAND4_X1 U6020 ( .A1(n5142), .A2(n5143), .A3(n5144), .A4(n5145), .ZN(n5141)
         );
  AOI221_X1 U6021 ( .B1(n13099), .B2(n774), .C1(n13096), .C2(n16019), .A(n5149), .ZN(n5142) );
  AOI221_X1 U6022 ( .B1(n13126), .B2(n773), .C1(n13123), .C2(n15983), .A(n5147), .ZN(n5144) );
  AOI221_X1 U6023 ( .B1(n13114), .B2(n14096), .C1(n13111), .C2(n15910), .A(
        n5148), .ZN(n5143) );
  NAND4_X1 U6024 ( .A1(n5105), .A2(n5106), .A3(n5107), .A4(n5108), .ZN(n5104)
         );
  AOI221_X1 U6025 ( .B1(n13100), .B2(n771), .C1(n13097), .C2(n16018), .A(n5112), .ZN(n5105) );
  AOI221_X1 U6026 ( .B1(n13127), .B2(n770), .C1(n13124), .C2(n15982), .A(n5110), .ZN(n5107) );
  AOI221_X1 U6027 ( .B1(n13115), .B2(n14095), .C1(n13112), .C2(n15909), .A(
        n5111), .ZN(n5106) );
  NAND4_X1 U6028 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n5071), .ZN(n5067)
         );
  AOI221_X1 U6029 ( .B1(n13100), .B2(n768), .C1(n13097), .C2(n16017), .A(n5075), .ZN(n5068) );
  AOI221_X1 U6030 ( .B1(n13127), .B2(n767), .C1(n13124), .C2(n15981), .A(n5073), .ZN(n5070) );
  AOI221_X1 U6031 ( .B1(n13115), .B2(n14094), .C1(n13112), .C2(n15908), .A(
        n5074), .ZN(n5069) );
  NAND4_X1 U6032 ( .A1(n5031), .A2(n5032), .A3(n5033), .A4(n5034), .ZN(n5030)
         );
  AOI221_X1 U6033 ( .B1(n13100), .B2(n765), .C1(n13097), .C2(n16016), .A(n5038), .ZN(n5031) );
  AOI221_X1 U6034 ( .B1(n13127), .B2(n764), .C1(n13124), .C2(n15980), .A(n5036), .ZN(n5033) );
  AOI221_X1 U6035 ( .B1(n13115), .B2(n14093), .C1(n13112), .C2(n15907), .A(
        n5037), .ZN(n5032) );
  NAND4_X1 U6036 ( .A1(n4994), .A2(n4995), .A3(n4996), .A4(n4997), .ZN(n4993)
         );
  AOI221_X1 U6037 ( .B1(n13100), .B2(n762), .C1(n13097), .C2(n16015), .A(n5001), .ZN(n4994) );
  AOI221_X1 U6038 ( .B1(n13127), .B2(n761), .C1(n13124), .C2(n15979), .A(n4999), .ZN(n4996) );
  AOI221_X1 U6039 ( .B1(n13115), .B2(n14092), .C1(n13112), .C2(n15906), .A(
        n5000), .ZN(n4995) );
  NAND4_X1 U6040 ( .A1(n4957), .A2(n4958), .A3(n4959), .A4(n4960), .ZN(n4956)
         );
  AOI221_X1 U6041 ( .B1(n13100), .B2(n759), .C1(n13097), .C2(n16014), .A(n4964), .ZN(n4957) );
  AOI221_X1 U6042 ( .B1(n13127), .B2(n758), .C1(n13124), .C2(n15978), .A(n4962), .ZN(n4959) );
  AOI221_X1 U6043 ( .B1(n13115), .B2(n14091), .C1(n13112), .C2(n15905), .A(
        n4963), .ZN(n4958) );
  NAND4_X1 U6044 ( .A1(n4920), .A2(n4921), .A3(n4922), .A4(n4923), .ZN(n4919)
         );
  AOI221_X1 U6045 ( .B1(n13100), .B2(n756), .C1(n13097), .C2(n16013), .A(n4927), .ZN(n4920) );
  AOI221_X1 U6046 ( .B1(n13127), .B2(n755), .C1(n13124), .C2(n15977), .A(n4925), .ZN(n4922) );
  AOI221_X1 U6047 ( .B1(n13115), .B2(n14090), .C1(n13112), .C2(n15904), .A(
        n4926), .ZN(n4921) );
  NAND4_X1 U6048 ( .A1(n4883), .A2(n4884), .A3(n4885), .A4(n4886), .ZN(n4882)
         );
  AOI221_X1 U6049 ( .B1(n13100), .B2(n753), .C1(n13097), .C2(n16012), .A(n4890), .ZN(n4883) );
  AOI221_X1 U6050 ( .B1(n13127), .B2(n752), .C1(n13124), .C2(n15976), .A(n4888), .ZN(n4885) );
  AOI221_X1 U6051 ( .B1(n13115), .B2(n14089), .C1(n13112), .C2(n15903), .A(
        n4889), .ZN(n4884) );
  NAND4_X1 U6052 ( .A1(n4846), .A2(n4847), .A3(n4848), .A4(n4849), .ZN(n4845)
         );
  AOI221_X1 U6053 ( .B1(n13100), .B2(n750), .C1(n13097), .C2(n16011), .A(n4853), .ZN(n4846) );
  AOI221_X1 U6054 ( .B1(n13127), .B2(n749), .C1(n13124), .C2(n15975), .A(n4851), .ZN(n4848) );
  AOI221_X1 U6055 ( .B1(n13115), .B2(n14088), .C1(n13112), .C2(n15902), .A(
        n4852), .ZN(n4847) );
  NAND4_X1 U6056 ( .A1(n4809), .A2(n4810), .A3(n4811), .A4(n4812), .ZN(n4808)
         );
  AOI221_X1 U6057 ( .B1(n13100), .B2(n747), .C1(n13097), .C2(n16010), .A(n4816), .ZN(n4809) );
  AOI221_X1 U6058 ( .B1(n13127), .B2(n746), .C1(n13124), .C2(n15974), .A(n4814), .ZN(n4811) );
  AOI221_X1 U6059 ( .B1(n13115), .B2(n14087), .C1(n13112), .C2(n15901), .A(
        n4815), .ZN(n4810) );
  NAND4_X1 U6060 ( .A1(n4772), .A2(n4773), .A3(n4774), .A4(n4775), .ZN(n4771)
         );
  AOI221_X1 U6061 ( .B1(n13100), .B2(n744), .C1(n13097), .C2(n16009), .A(n4779), .ZN(n4772) );
  AOI221_X1 U6062 ( .B1(n13127), .B2(n743), .C1(n13124), .C2(n15973), .A(n4777), .ZN(n4774) );
  AOI221_X1 U6063 ( .B1(n13115), .B2(n14086), .C1(n13112), .C2(n15900), .A(
        n4778), .ZN(n4773) );
  NAND4_X1 U6064 ( .A1(n4735), .A2(n4736), .A3(n4737), .A4(n4738), .ZN(n4734)
         );
  AOI221_X1 U6065 ( .B1(n13100), .B2(n741), .C1(n13097), .C2(n16008), .A(n4742), .ZN(n4735) );
  AOI221_X1 U6066 ( .B1(n13127), .B2(n740), .C1(n13124), .C2(n15972), .A(n4740), .ZN(n4737) );
  AOI221_X1 U6067 ( .B1(n13115), .B2(n14085), .C1(n13112), .C2(n15899), .A(
        n4741), .ZN(n4736) );
  NAND4_X1 U6068 ( .A1(n4698), .A2(n4699), .A3(n4700), .A4(n4701), .ZN(n4697)
         );
  AOI221_X1 U6069 ( .B1(n13100), .B2(n738), .C1(n13097), .C2(n16007), .A(n4705), .ZN(n4698) );
  AOI221_X1 U6070 ( .B1(n13127), .B2(n737), .C1(n13124), .C2(n15971), .A(n4703), .ZN(n4700) );
  AOI221_X1 U6071 ( .B1(n13115), .B2(n14084), .C1(n13112), .C2(n15898), .A(
        n4704), .ZN(n4699) );
  NAND4_X1 U6072 ( .A1(n4661), .A2(n4662), .A3(n4663), .A4(n4664), .ZN(n4660)
         );
  AOI221_X1 U6073 ( .B1(n13101), .B2(n735), .C1(n13098), .C2(n15946), .A(n4668), .ZN(n4661) );
  AOI221_X1 U6074 ( .B1(n13128), .B2(n734), .C1(n13125), .C2(n15938), .A(n4666), .ZN(n4663) );
  AOI221_X1 U6075 ( .B1(n13116), .B2(n14083), .C1(n13113), .C2(n15605), .A(
        n4667), .ZN(n4662) );
  NAND4_X1 U6076 ( .A1(n3163), .A2(n3164), .A3(n3165), .A4(n3166), .ZN(n3153)
         );
  AOI221_X1 U6077 ( .B1(n13275), .B2(n15863), .C1(n13272), .C2(n99), .A(n3170), 
        .ZN(n3163) );
  AOI221_X1 U6078 ( .B1(n13302), .B2(n15575), .C1(n13299), .C2(n15791), .A(
        n3168), .ZN(n3165) );
  AOI221_X1 U6079 ( .B1(n13290), .B2(n14462), .C1(n13287), .C2(n15583), .A(
        n3169), .ZN(n3164) );
  NAND4_X1 U6080 ( .A1(n3072), .A2(n3073), .A3(n3074), .A4(n3075), .ZN(n3044)
         );
  AOI221_X1 U6081 ( .B1(n13275), .B2(n15862), .C1(n13272), .C2(n97), .A(n3095), 
        .ZN(n3072) );
  AOI221_X1 U6082 ( .B1(n13302), .B2(n15574), .C1(n13299), .C2(n15790), .A(
        n3084), .ZN(n3074) );
  AOI221_X1 U6083 ( .B1(n13290), .B2(n14461), .C1(n13287), .C2(n15582), .A(
        n3089), .ZN(n3073) );
  NAND4_X1 U6084 ( .A1(n4447), .A2(n4448), .A3(n4449), .A4(n4450), .ZN(n4437)
         );
  AOI221_X1 U6085 ( .B1(n13047), .B2(n15863), .C1(n13044), .C2(n99), .A(n4454), 
        .ZN(n4447) );
  AOI221_X1 U6086 ( .B1(n13074), .B2(n15791), .C1(n13071), .C2(n15575), .A(
        n4452), .ZN(n4449) );
  AOI221_X1 U6087 ( .B1(n13062), .B2(n14462), .C1(n13059), .C2(n15583), .A(
        n4453), .ZN(n4448) );
  NAND4_X1 U6088 ( .A1(n4356), .A2(n4357), .A3(n4358), .A4(n4359), .ZN(n4328)
         );
  AOI221_X1 U6089 ( .B1(n13047), .B2(n15862), .C1(n13044), .C2(n97), .A(n4379), 
        .ZN(n4356) );
  AOI221_X1 U6090 ( .B1(n13074), .B2(n15790), .C1(n13071), .C2(n15574), .A(
        n4368), .ZN(n4358) );
  AOI221_X1 U6091 ( .B1(n13062), .B2(n14461), .C1(n13059), .C2(n15582), .A(
        n4373), .ZN(n4357) );
  OAI21_X1 U6092 ( .B1(n13149), .B2(n1576), .A(n14026), .ZN(n7546) );
  OAI21_X1 U6093 ( .B1(n13149), .B2(n1545), .A(n14024), .ZN(n7608) );
  OAI21_X1 U6094 ( .B1(n13377), .B2(n1544), .A(n14024), .ZN(n7610) );
  OAI21_X1 U6095 ( .B1(n13377), .B2(n1513), .A(n14022), .ZN(n7672) );
  OAI21_X1 U6096 ( .B1(n13148), .B2(n1575), .A(n14026), .ZN(n7548) );
  OAI21_X1 U6097 ( .B1(n13148), .B2(n1574), .A(n14026), .ZN(n7550) );
  OAI21_X1 U6098 ( .B1(n13148), .B2(n1573), .A(n14026), .ZN(n7552) );
  OAI21_X1 U6099 ( .B1(n13148), .B2(n1572), .A(n14026), .ZN(n7554) );
  OAI21_X1 U6100 ( .B1(n13147), .B2(n1571), .A(n14026), .ZN(n7556) );
  OAI21_X1 U6101 ( .B1(n13147), .B2(n1570), .A(n14026), .ZN(n7558) );
  OAI21_X1 U6102 ( .B1(n13147), .B2(n1569), .A(n14026), .ZN(n7560) );
  OAI21_X1 U6103 ( .B1(n13147), .B2(n1568), .A(n14026), .ZN(n7562) );
  OAI21_X1 U6104 ( .B1(n13147), .B2(n1566), .A(n14026), .ZN(n7566) );
  OAI21_X1 U6105 ( .B1(n13147), .B2(n1564), .A(n14026), .ZN(n7570) );
  OAI21_X1 U6106 ( .B1(n13147), .B2(n1561), .A(n14025), .ZN(n7576) );
  OAI21_X1 U6107 ( .B1(n13147), .B2(n1560), .A(n14025), .ZN(n7578) );
  OAI21_X1 U6108 ( .B1(n13147), .B2(n1559), .A(n14025), .ZN(n7580) );
  OAI21_X1 U6109 ( .B1(n13147), .B2(n1558), .A(n14025), .ZN(n7582) );
  OAI21_X1 U6110 ( .B1(n13147), .B2(n1557), .A(n14025), .ZN(n7584) );
  OAI21_X1 U6111 ( .B1(n13147), .B2(n1556), .A(n14025), .ZN(n7586) );
  OAI21_X1 U6112 ( .B1(n13148), .B2(n1555), .A(n14025), .ZN(n7588) );
  OAI21_X1 U6113 ( .B1(n13147), .B2(n1554), .A(n14025), .ZN(n7590) );
  OAI21_X1 U6114 ( .B1(n13148), .B2(n1553), .A(n14025), .ZN(n7592) );
  OAI21_X1 U6115 ( .B1(n13148), .B2(n1552), .A(n14025), .ZN(n7594) );
  OAI21_X1 U6116 ( .B1(n13148), .B2(n1551), .A(n14025), .ZN(n7596) );
  OAI21_X1 U6117 ( .B1(n13148), .B2(n1550), .A(n14024), .ZN(n7598) );
  OAI21_X1 U6118 ( .B1(n13148), .B2(n1549), .A(n14024), .ZN(n7600) );
  OAI21_X1 U6119 ( .B1(n13148), .B2(n1548), .A(n14024), .ZN(n7602) );
  OAI21_X1 U6120 ( .B1(n13148), .B2(n1547), .A(n14024), .ZN(n7604) );
  OAI21_X1 U6121 ( .B1(n13148), .B2(n1546), .A(n14024), .ZN(n7606) );
  OAI21_X1 U6122 ( .B1(n13376), .B2(n1543), .A(n14024), .ZN(n7612) );
  OAI21_X1 U6123 ( .B1(n13376), .B2(n1542), .A(n14024), .ZN(n7614) );
  OAI21_X1 U6124 ( .B1(n13376), .B2(n1541), .A(n14024), .ZN(n7616) );
  OAI21_X1 U6125 ( .B1(n13376), .B2(n1540), .A(n14024), .ZN(n7618) );
  OAI21_X1 U6126 ( .B1(n13375), .B2(n1539), .A(n14024), .ZN(n7620) );
  OAI21_X1 U6127 ( .B1(n13375), .B2(n1538), .A(n14023), .ZN(n7622) );
  OAI21_X1 U6128 ( .B1(n13375), .B2(n1537), .A(n14023), .ZN(n7624) );
  OAI21_X1 U6129 ( .B1(n13375), .B2(n1536), .A(n14023), .ZN(n7626) );
  OAI21_X1 U6130 ( .B1(n13375), .B2(n1534), .A(n14023), .ZN(n7630) );
  OAI21_X1 U6131 ( .B1(n13375), .B2(n1532), .A(n14023), .ZN(n7634) );
  OAI21_X1 U6132 ( .B1(n13375), .B2(n1529), .A(n14023), .ZN(n7640) );
  OAI21_X1 U6133 ( .B1(n13375), .B2(n1528), .A(n14024), .ZN(n7642) );
  OAI21_X1 U6134 ( .B1(n13375), .B2(n1527), .A(n14023), .ZN(n7644) );
  OAI21_X1 U6135 ( .B1(n13375), .B2(n1526), .A(n14023), .ZN(n7646) );
  OAI21_X1 U6136 ( .B1(n13375), .B2(n1525), .A(n14022), .ZN(n7648) );
  OAI21_X1 U6137 ( .B1(n13375), .B2(n1524), .A(n14023), .ZN(n7650) );
  OAI21_X1 U6138 ( .B1(n13376), .B2(n1523), .A(n14022), .ZN(n7652) );
  OAI21_X1 U6139 ( .B1(n13375), .B2(n1522), .A(n14022), .ZN(n7654) );
  OAI21_X1 U6140 ( .B1(n13376), .B2(n1521), .A(n14022), .ZN(n7656) );
  OAI21_X1 U6141 ( .B1(n13376), .B2(n1520), .A(n14022), .ZN(n7658) );
  OAI21_X1 U6142 ( .B1(n13376), .B2(n1519), .A(n14022), .ZN(n7660) );
  OAI21_X1 U6143 ( .B1(n13376), .B2(n1518), .A(n14022), .ZN(n7662) );
  OAI21_X1 U6144 ( .B1(n13376), .B2(n1517), .A(n14022), .ZN(n7664) );
  OAI21_X1 U6145 ( .B1(n13376), .B2(n1516), .A(n14022), .ZN(n7666) );
  OAI21_X1 U6146 ( .B1(n13376), .B2(n1515), .A(n14022), .ZN(n7668) );
  OAI21_X1 U6147 ( .B1(n13376), .B2(n1514), .A(n14022), .ZN(n7670) );
  OAI21_X1 U6148 ( .B1(n13146), .B2(n1567), .A(n14026), .ZN(n7564) );
  OAI21_X1 U6149 ( .B1(n13146), .B2(n1565), .A(n14026), .ZN(n7568) );
  OAI21_X1 U6150 ( .B1(n13146), .B2(n1563), .A(n14025), .ZN(n7572) );
  OAI21_X1 U6151 ( .B1(n13146), .B2(n1562), .A(n14025), .ZN(n7574) );
  OAI21_X1 U6152 ( .B1(n13374), .B2(n1535), .A(n14023), .ZN(n7628) );
  OAI21_X1 U6153 ( .B1(n13374), .B2(n1533), .A(n14023), .ZN(n7632) );
  OAI21_X1 U6154 ( .B1(n13374), .B2(n1531), .A(n14023), .ZN(n7636) );
  OAI21_X1 U6155 ( .B1(n13374), .B2(n1530), .A(n14023), .ZN(n7638) );
  OAI22_X1 U6156 ( .A1(n13828), .A2(n13431), .B1(n13426), .B2(n12774), .ZN(
        n7898) );
  OAI22_X1 U6157 ( .A1(n13835), .A2(n13431), .B1(n13426), .B2(n12775), .ZN(
        n7899) );
  OAI22_X1 U6158 ( .A1(n13841), .A2(n13431), .B1(n13426), .B2(n12776), .ZN(
        n7900) );
  OAI22_X1 U6159 ( .A1(n13847), .A2(n13431), .B1(n13426), .B2(n12777), .ZN(
        n7901) );
  OAI22_X1 U6160 ( .A1(n13853), .A2(n13431), .B1(n13426), .B2(n12778), .ZN(
        n7902) );
  OAI22_X1 U6161 ( .A1(n13859), .A2(n13431), .B1(n13426), .B2(n12779), .ZN(
        n7903) );
  OAI22_X1 U6162 ( .A1(n13865), .A2(n13431), .B1(n13426), .B2(n12780), .ZN(
        n7904) );
  OAI22_X1 U6163 ( .A1(n13871), .A2(n13431), .B1(n13426), .B2(n12781), .ZN(
        n7905) );
  OAI22_X1 U6164 ( .A1(n13877), .A2(n13430), .B1(n13426), .B2(n12782), .ZN(
        n7906) );
  OAI22_X1 U6165 ( .A1(n13883), .A2(n13430), .B1(n13426), .B2(n12783), .ZN(
        n7907) );
  OAI22_X1 U6166 ( .A1(n13889), .A2(n13430), .B1(n13426), .B2(n12784), .ZN(
        n7908) );
  OAI22_X1 U6167 ( .A1(n13895), .A2(n13430), .B1(n13426), .B2(n12785), .ZN(
        n7909) );
  OAI22_X1 U6168 ( .A1(n13901), .A2(n13430), .B1(n13427), .B2(n12786), .ZN(
        n7910) );
  OAI22_X1 U6169 ( .A1(n13907), .A2(n13430), .B1(n13427), .B2(n12787), .ZN(
        n7911) );
  OAI22_X1 U6170 ( .A1(n13913), .A2(n13430), .B1(n13427), .B2(n12788), .ZN(
        n7912) );
  OAI22_X1 U6171 ( .A1(n13919), .A2(n13430), .B1(n13427), .B2(n12789), .ZN(
        n7913) );
  OAI22_X1 U6172 ( .A1(n13925), .A2(n13430), .B1(n13427), .B2(n12790), .ZN(
        n7914) );
  OAI22_X1 U6173 ( .A1(n13931), .A2(n13430), .B1(n13427), .B2(n12791), .ZN(
        n7915) );
  OAI22_X1 U6174 ( .A1(n13937), .A2(n13430), .B1(n13427), .B2(n12792), .ZN(
        n7916) );
  OAI22_X1 U6175 ( .A1(n13943), .A2(n13430), .B1(n13427), .B2(n12793), .ZN(
        n7917) );
  OAI22_X1 U6176 ( .A1(n13949), .A2(n13429), .B1(n13427), .B2(n12794), .ZN(
        n7918) );
  OAI22_X1 U6177 ( .A1(n13955), .A2(n13429), .B1(n13427), .B2(n12795), .ZN(
        n7919) );
  OAI22_X1 U6178 ( .A1(n13961), .A2(n13429), .B1(n13427), .B2(n12796), .ZN(
        n7920) );
  OAI22_X1 U6179 ( .A1(n13967), .A2(n13429), .B1(n13427), .B2(n12797), .ZN(
        n7921) );
  OAI22_X1 U6180 ( .A1(n13973), .A2(n13429), .B1(n13428), .B2(n12798), .ZN(
        n7922) );
  OAI22_X1 U6181 ( .A1(n13979), .A2(n13429), .B1(n13428), .B2(n12799), .ZN(
        n7923) );
  OAI22_X1 U6182 ( .A1(n13985), .A2(n13429), .B1(n13428), .B2(n12800), .ZN(
        n7924) );
  OAI22_X1 U6183 ( .A1(n13991), .A2(n13429), .B1(n13428), .B2(n12801), .ZN(
        n7925) );
  OAI22_X1 U6184 ( .A1(n13997), .A2(n13429), .B1(n13428), .B2(n12802), .ZN(
        n7926) );
  OAI22_X1 U6185 ( .A1(n14003), .A2(n13429), .B1(n13428), .B2(n12803), .ZN(
        n7927) );
  OAI22_X1 U6186 ( .A1(n14009), .A2(n13429), .B1(n13428), .B2(n12804), .ZN(
        n7928) );
  OAI22_X1 U6187 ( .A1(n14018), .A2(n13429), .B1(n13428), .B2(n12805), .ZN(
        n7929) );
  OAI22_X1 U6188 ( .A1(n13828), .A2(n13461), .B1(n13456), .B2(n12806), .ZN(
        n8058) );
  OAI22_X1 U6189 ( .A1(n13834), .A2(n13461), .B1(n13456), .B2(n12807), .ZN(
        n8059) );
  OAI22_X1 U6190 ( .A1(n13840), .A2(n13461), .B1(n13456), .B2(n12808), .ZN(
        n8060) );
  OAI22_X1 U6191 ( .A1(n13846), .A2(n13461), .B1(n13456), .B2(n12809), .ZN(
        n8061) );
  OAI22_X1 U6192 ( .A1(n13852), .A2(n13461), .B1(n13456), .B2(n12810), .ZN(
        n8062) );
  OAI22_X1 U6193 ( .A1(n13858), .A2(n13461), .B1(n13456), .B2(n12811), .ZN(
        n8063) );
  OAI22_X1 U6194 ( .A1(n13864), .A2(n13461), .B1(n13456), .B2(n12812), .ZN(
        n8064) );
  OAI22_X1 U6195 ( .A1(n13870), .A2(n13461), .B1(n13456), .B2(n12813), .ZN(
        n8065) );
  OAI22_X1 U6196 ( .A1(n13876), .A2(n13460), .B1(n13456), .B2(n12814), .ZN(
        n8066) );
  OAI22_X1 U6197 ( .A1(n13882), .A2(n13460), .B1(n13456), .B2(n12815), .ZN(
        n8067) );
  OAI22_X1 U6198 ( .A1(n13888), .A2(n13460), .B1(n13456), .B2(n12816), .ZN(
        n8068) );
  OAI22_X1 U6199 ( .A1(n13894), .A2(n13460), .B1(n13456), .B2(n12817), .ZN(
        n8069) );
  OAI22_X1 U6200 ( .A1(n13900), .A2(n13460), .B1(n13457), .B2(n12818), .ZN(
        n8070) );
  OAI22_X1 U6201 ( .A1(n13906), .A2(n13460), .B1(n13457), .B2(n12819), .ZN(
        n8071) );
  OAI22_X1 U6202 ( .A1(n13912), .A2(n13460), .B1(n13457), .B2(n12820), .ZN(
        n8072) );
  OAI22_X1 U6203 ( .A1(n13918), .A2(n13460), .B1(n13457), .B2(n12821), .ZN(
        n8073) );
  OAI22_X1 U6204 ( .A1(n13924), .A2(n13460), .B1(n13457), .B2(n12822), .ZN(
        n8074) );
  OAI22_X1 U6205 ( .A1(n13930), .A2(n13460), .B1(n13457), .B2(n12823), .ZN(
        n8075) );
  OAI22_X1 U6206 ( .A1(n13936), .A2(n13460), .B1(n13457), .B2(n12824), .ZN(
        n8076) );
  OAI22_X1 U6207 ( .A1(n13942), .A2(n13460), .B1(n13457), .B2(n12825), .ZN(
        n8077) );
  OAI22_X1 U6208 ( .A1(n13948), .A2(n13459), .B1(n13457), .B2(n12826), .ZN(
        n8078) );
  OAI22_X1 U6209 ( .A1(n13954), .A2(n13459), .B1(n13457), .B2(n12827), .ZN(
        n8079) );
  OAI22_X1 U6210 ( .A1(n13960), .A2(n13459), .B1(n13457), .B2(n12828), .ZN(
        n8080) );
  OAI22_X1 U6211 ( .A1(n13966), .A2(n13459), .B1(n13457), .B2(n12829), .ZN(
        n8081) );
  OAI22_X1 U6212 ( .A1(n13972), .A2(n13459), .B1(n13458), .B2(n12830), .ZN(
        n8082) );
  OAI22_X1 U6213 ( .A1(n13978), .A2(n13459), .B1(n13458), .B2(n12831), .ZN(
        n8083) );
  OAI22_X1 U6214 ( .A1(n13984), .A2(n13459), .B1(n13458), .B2(n12832), .ZN(
        n8084) );
  OAI22_X1 U6215 ( .A1(n13990), .A2(n13459), .B1(n13458), .B2(n12833), .ZN(
        n8085) );
  OAI22_X1 U6216 ( .A1(n13996), .A2(n13459), .B1(n13458), .B2(n12834), .ZN(
        n8086) );
  OAI22_X1 U6217 ( .A1(n14002), .A2(n13459), .B1(n13458), .B2(n12835), .ZN(
        n8087) );
  OAI22_X1 U6218 ( .A1(n14008), .A2(n13459), .B1(n13458), .B2(n12836), .ZN(
        n8088) );
  OAI22_X1 U6219 ( .A1(n14017), .A2(n13459), .B1(n13458), .B2(n12837), .ZN(
        n8089) );
  OAI22_X1 U6220 ( .A1(n13827), .A2(n13539), .B1(n13534), .B2(n12838), .ZN(
        n8474) );
  OAI22_X1 U6221 ( .A1(n13833), .A2(n13539), .B1(n13534), .B2(n12839), .ZN(
        n8475) );
  OAI22_X1 U6222 ( .A1(n13839), .A2(n13539), .B1(n13534), .B2(n12840), .ZN(
        n8476) );
  OAI22_X1 U6223 ( .A1(n13845), .A2(n13539), .B1(n13534), .B2(n12841), .ZN(
        n8477) );
  OAI22_X1 U6224 ( .A1(n13851), .A2(n13539), .B1(n13534), .B2(n12842), .ZN(
        n8478) );
  OAI22_X1 U6225 ( .A1(n13857), .A2(n13539), .B1(n13534), .B2(n12843), .ZN(
        n8479) );
  OAI22_X1 U6226 ( .A1(n13863), .A2(n13539), .B1(n13534), .B2(n12844), .ZN(
        n8480) );
  OAI22_X1 U6227 ( .A1(n13869), .A2(n13539), .B1(n13534), .B2(n12845), .ZN(
        n8481) );
  OAI22_X1 U6228 ( .A1(n13875), .A2(n13538), .B1(n13534), .B2(n12846), .ZN(
        n8482) );
  OAI22_X1 U6229 ( .A1(n13881), .A2(n13538), .B1(n13534), .B2(n12847), .ZN(
        n8483) );
  OAI22_X1 U6230 ( .A1(n13887), .A2(n13538), .B1(n13534), .B2(n12848), .ZN(
        n8484) );
  OAI22_X1 U6231 ( .A1(n13893), .A2(n13538), .B1(n13534), .B2(n12849), .ZN(
        n8485) );
  OAI22_X1 U6232 ( .A1(n13899), .A2(n13538), .B1(n13535), .B2(n12850), .ZN(
        n8486) );
  OAI22_X1 U6233 ( .A1(n13905), .A2(n13538), .B1(n13535), .B2(n12851), .ZN(
        n8487) );
  OAI22_X1 U6234 ( .A1(n13911), .A2(n13538), .B1(n13535), .B2(n12852), .ZN(
        n8488) );
  OAI22_X1 U6235 ( .A1(n13917), .A2(n13538), .B1(n13535), .B2(n12853), .ZN(
        n8489) );
  OAI22_X1 U6236 ( .A1(n13923), .A2(n13538), .B1(n13535), .B2(n12854), .ZN(
        n8490) );
  OAI22_X1 U6237 ( .A1(n13929), .A2(n13538), .B1(n13535), .B2(n12855), .ZN(
        n8491) );
  OAI22_X1 U6238 ( .A1(n13935), .A2(n13538), .B1(n13535), .B2(n12856), .ZN(
        n8492) );
  OAI22_X1 U6239 ( .A1(n13941), .A2(n13538), .B1(n13535), .B2(n12857), .ZN(
        n8493) );
  OAI22_X1 U6240 ( .A1(n13947), .A2(n13537), .B1(n13535), .B2(n12858), .ZN(
        n8494) );
  OAI22_X1 U6241 ( .A1(n13953), .A2(n13537), .B1(n13535), .B2(n12859), .ZN(
        n8495) );
  OAI22_X1 U6242 ( .A1(n13959), .A2(n13537), .B1(n13535), .B2(n12860), .ZN(
        n8496) );
  OAI22_X1 U6243 ( .A1(n13965), .A2(n13537), .B1(n13535), .B2(n12861), .ZN(
        n8497) );
  OAI22_X1 U6244 ( .A1(n13971), .A2(n13537), .B1(n13536), .B2(n12862), .ZN(
        n8498) );
  OAI22_X1 U6245 ( .A1(n13977), .A2(n13537), .B1(n13536), .B2(n12863), .ZN(
        n8499) );
  OAI22_X1 U6246 ( .A1(n13983), .A2(n13537), .B1(n13536), .B2(n12864), .ZN(
        n8500) );
  OAI22_X1 U6247 ( .A1(n13989), .A2(n13537), .B1(n13536), .B2(n12865), .ZN(
        n8501) );
  OAI22_X1 U6248 ( .A1(n13995), .A2(n13537), .B1(n13536), .B2(n12866), .ZN(
        n8502) );
  OAI22_X1 U6249 ( .A1(n14001), .A2(n13537), .B1(n13536), .B2(n12867), .ZN(
        n8503) );
  OAI22_X1 U6250 ( .A1(n14007), .A2(n13537), .B1(n13536), .B2(n12868), .ZN(
        n8504) );
  OAI22_X1 U6251 ( .A1(n14016), .A2(n13537), .B1(n13536), .B2(n12869), .ZN(
        n8505) );
  OAI22_X1 U6252 ( .A1(n13827), .A2(n13569), .B1(n13564), .B2(n12870), .ZN(
        n8634) );
  OAI22_X1 U6253 ( .A1(n13833), .A2(n13569), .B1(n13564), .B2(n12871), .ZN(
        n8635) );
  OAI22_X1 U6254 ( .A1(n13839), .A2(n13569), .B1(n13564), .B2(n12872), .ZN(
        n8636) );
  OAI22_X1 U6255 ( .A1(n13845), .A2(n13569), .B1(n13564), .B2(n12873), .ZN(
        n8637) );
  OAI22_X1 U6256 ( .A1(n13851), .A2(n13569), .B1(n13564), .B2(n12874), .ZN(
        n8638) );
  OAI22_X1 U6257 ( .A1(n13857), .A2(n13569), .B1(n13564), .B2(n12875), .ZN(
        n8639) );
  OAI22_X1 U6258 ( .A1(n13863), .A2(n13569), .B1(n13564), .B2(n12876), .ZN(
        n8640) );
  OAI22_X1 U6259 ( .A1(n13869), .A2(n13569), .B1(n13564), .B2(n12877), .ZN(
        n8641) );
  OAI22_X1 U6260 ( .A1(n13875), .A2(n13568), .B1(n13564), .B2(n12878), .ZN(
        n8642) );
  OAI22_X1 U6261 ( .A1(n13881), .A2(n13568), .B1(n13564), .B2(n12879), .ZN(
        n8643) );
  OAI22_X1 U6262 ( .A1(n13887), .A2(n13568), .B1(n13564), .B2(n12880), .ZN(
        n8644) );
  OAI22_X1 U6263 ( .A1(n13893), .A2(n13568), .B1(n13564), .B2(n12881), .ZN(
        n8645) );
  OAI22_X1 U6264 ( .A1(n13899), .A2(n13568), .B1(n13565), .B2(n12882), .ZN(
        n8646) );
  OAI22_X1 U6265 ( .A1(n13905), .A2(n13568), .B1(n13565), .B2(n12883), .ZN(
        n8647) );
  OAI22_X1 U6266 ( .A1(n13911), .A2(n13568), .B1(n13565), .B2(n12884), .ZN(
        n8648) );
  OAI22_X1 U6267 ( .A1(n13917), .A2(n13568), .B1(n13565), .B2(n12885), .ZN(
        n8649) );
  OAI22_X1 U6268 ( .A1(n13923), .A2(n13568), .B1(n13565), .B2(n12886), .ZN(
        n8650) );
  OAI22_X1 U6269 ( .A1(n13929), .A2(n13568), .B1(n13565), .B2(n12887), .ZN(
        n8651) );
  OAI22_X1 U6270 ( .A1(n13935), .A2(n13568), .B1(n13565), .B2(n12888), .ZN(
        n8652) );
  OAI22_X1 U6271 ( .A1(n13941), .A2(n13568), .B1(n13565), .B2(n12889), .ZN(
        n8653) );
  OAI22_X1 U6272 ( .A1(n13947), .A2(n13567), .B1(n13565), .B2(n12890), .ZN(
        n8654) );
  OAI22_X1 U6273 ( .A1(n13953), .A2(n13567), .B1(n13565), .B2(n12891), .ZN(
        n8655) );
  OAI22_X1 U6274 ( .A1(n13959), .A2(n13567), .B1(n13565), .B2(n12892), .ZN(
        n8656) );
  OAI22_X1 U6275 ( .A1(n13965), .A2(n13567), .B1(n13565), .B2(n12893), .ZN(
        n8657) );
  OAI22_X1 U6276 ( .A1(n13971), .A2(n13567), .B1(n13566), .B2(n12894), .ZN(
        n8658) );
  OAI22_X1 U6277 ( .A1(n13977), .A2(n13567), .B1(n13566), .B2(n12895), .ZN(
        n8659) );
  OAI22_X1 U6278 ( .A1(n13983), .A2(n13567), .B1(n13566), .B2(n12896), .ZN(
        n8660) );
  OAI22_X1 U6279 ( .A1(n13989), .A2(n13567), .B1(n13566), .B2(n12897), .ZN(
        n8661) );
  OAI22_X1 U6280 ( .A1(n13995), .A2(n13567), .B1(n13566), .B2(n12898), .ZN(
        n8662) );
  OAI22_X1 U6281 ( .A1(n14001), .A2(n13567), .B1(n13566), .B2(n12899), .ZN(
        n8663) );
  OAI22_X1 U6282 ( .A1(n14007), .A2(n13567), .B1(n13566), .B2(n12900), .ZN(
        n8664) );
  OAI22_X1 U6283 ( .A1(n14016), .A2(n13567), .B1(n13566), .B2(n12901), .ZN(
        n8665) );
  OAI22_X1 U6284 ( .A1(n13826), .A2(n13587), .B1(n13584), .B2(n12902), .ZN(
        n8730) );
  OAI22_X1 U6285 ( .A1(n13833), .A2(n13587), .B1(n13584), .B2(n12903), .ZN(
        n8731) );
  OAI22_X1 U6286 ( .A1(n13839), .A2(n13587), .B1(n13584), .B2(n12904), .ZN(
        n8732) );
  OAI22_X1 U6287 ( .A1(n13845), .A2(n13587), .B1(n13584), .B2(n12905), .ZN(
        n8733) );
  OAI22_X1 U6288 ( .A1(n13851), .A2(n13587), .B1(n13584), .B2(n12906), .ZN(
        n8734) );
  OAI22_X1 U6289 ( .A1(n13857), .A2(n13587), .B1(n13584), .B2(n12907), .ZN(
        n8735) );
  OAI22_X1 U6290 ( .A1(n13863), .A2(n13587), .B1(n13584), .B2(n12908), .ZN(
        n8736) );
  OAI22_X1 U6291 ( .A1(n13869), .A2(n13587), .B1(n13583), .B2(n12909), .ZN(
        n8737) );
  OAI22_X1 U6292 ( .A1(n13875), .A2(n13586), .B1(n13583), .B2(n12910), .ZN(
        n8738) );
  OAI22_X1 U6293 ( .A1(n13881), .A2(n13586), .B1(n13583), .B2(n12911), .ZN(
        n8739) );
  OAI22_X1 U6294 ( .A1(n13887), .A2(n13586), .B1(n13583), .B2(n12912), .ZN(
        n8740) );
  OAI22_X1 U6295 ( .A1(n13893), .A2(n13586), .B1(n13583), .B2(n12913), .ZN(
        n8741) );
  OAI22_X1 U6296 ( .A1(n13899), .A2(n13586), .B1(n13583), .B2(n12914), .ZN(
        n8742) );
  OAI22_X1 U6297 ( .A1(n13905), .A2(n13586), .B1(n13583), .B2(n12915), .ZN(
        n8743) );
  OAI22_X1 U6298 ( .A1(n13911), .A2(n13586), .B1(n13583), .B2(n12916), .ZN(
        n8744) );
  OAI22_X1 U6299 ( .A1(n13917), .A2(n13586), .B1(n13583), .B2(n12917), .ZN(
        n8745) );
  OAI22_X1 U6300 ( .A1(n13923), .A2(n13586), .B1(n13583), .B2(n12918), .ZN(
        n8746) );
  OAI22_X1 U6301 ( .A1(n13929), .A2(n13586), .B1(n13583), .B2(n12919), .ZN(
        n8747) );
  OAI22_X1 U6302 ( .A1(n13935), .A2(n13586), .B1(n13583), .B2(n12920), .ZN(
        n8748) );
  OAI22_X1 U6303 ( .A1(n13941), .A2(n13586), .B1(n13583), .B2(n12921), .ZN(
        n8749) );
  BUF_X1 U6304 ( .A(ENABLE), .Z(n14022) );
  BUF_X1 U6305 ( .A(ENABLE), .Z(n14026) );
  BUF_X1 U6306 ( .A(ENABLE), .Z(n14025) );
  BUF_X1 U6307 ( .A(ENABLE), .Z(n14024) );
  BUF_X1 U6308 ( .A(ENABLE), .Z(n14023) );
  NAND2_X1 U6309 ( .A1(DATAIN[0]), .A2(n13821), .ZN(n2865) );
  NAND2_X1 U6310 ( .A1(DATAIN[1]), .A2(n13821), .ZN(n2864) );
  NAND2_X1 U6311 ( .A1(DATAIN[2]), .A2(n13821), .ZN(n2863) );
  NAND2_X1 U6312 ( .A1(DATAIN[3]), .A2(n13821), .ZN(n2862) );
  NAND2_X1 U6313 ( .A1(DATAIN[4]), .A2(n13820), .ZN(n2861) );
  NAND2_X1 U6314 ( .A1(DATAIN[5]), .A2(n13820), .ZN(n2860) );
  NAND2_X1 U6315 ( .A1(DATAIN[6]), .A2(n13820), .ZN(n2859) );
  NAND2_X1 U6316 ( .A1(DATAIN[7]), .A2(n13820), .ZN(n2858) );
  NAND2_X1 U6317 ( .A1(DATAIN[8]), .A2(n13819), .ZN(n2857) );
  NAND2_X1 U6318 ( .A1(DATAIN[9]), .A2(n13819), .ZN(n2856) );
  NAND2_X1 U6319 ( .A1(DATAIN[10]), .A2(n13819), .ZN(n2855) );
  NAND2_X1 U6320 ( .A1(DATAIN[11]), .A2(n13819), .ZN(n2854) );
  NAND2_X1 U6321 ( .A1(DATAIN[12]), .A2(n13818), .ZN(n2853) );
  NAND2_X1 U6322 ( .A1(DATAIN[13]), .A2(n13818), .ZN(n2852) );
  NAND2_X1 U6323 ( .A1(DATAIN[14]), .A2(n13818), .ZN(n2851) );
  NAND2_X1 U6324 ( .A1(DATAIN[15]), .A2(n13818), .ZN(n2850) );
  NAND2_X1 U6325 ( .A1(DATAIN[16]), .A2(n13817), .ZN(n2849) );
  NAND2_X1 U6326 ( .A1(DATAIN[17]), .A2(n13817), .ZN(n2848) );
  NAND2_X1 U6327 ( .A1(DATAIN[18]), .A2(n13817), .ZN(n2847) );
  NAND2_X1 U6328 ( .A1(DATAIN[19]), .A2(n13817), .ZN(n2846) );
  NAND2_X1 U6329 ( .A1(DATAIN[20]), .A2(n13816), .ZN(n2845) );
  NAND2_X1 U6330 ( .A1(DATAIN[21]), .A2(n13816), .ZN(n2844) );
  NAND2_X1 U6331 ( .A1(DATAIN[22]), .A2(n13816), .ZN(n2843) );
  NAND2_X1 U6332 ( .A1(DATAIN[23]), .A2(n13816), .ZN(n2842) );
  NAND2_X1 U6333 ( .A1(DATAIN[24]), .A2(n13815), .ZN(n2841) );
  NAND2_X1 U6334 ( .A1(DATAIN[25]), .A2(n13815), .ZN(n2840) );
  NAND2_X1 U6335 ( .A1(DATAIN[26]), .A2(n13815), .ZN(n2839) );
  NAND2_X1 U6336 ( .A1(DATAIN[27]), .A2(n13815), .ZN(n2838) );
  NAND2_X1 U6337 ( .A1(DATAIN[28]), .A2(n13814), .ZN(n2837) );
  NAND2_X1 U6338 ( .A1(DATAIN[29]), .A2(n13814), .ZN(n2836) );
  NAND2_X1 U6339 ( .A1(DATAIN[30]), .A2(n13814), .ZN(n2835) );
  NAND2_X1 U6340 ( .A1(DATAIN[31]), .A2(n13814), .ZN(n2833) );
  INV_X1 U6341 ( .A(RESET), .ZN(n16063) );
  BUF_X1 U6342 ( .A(n2866), .Z(n13810) );
  NAND2_X1 U6343 ( .A1(WR), .A2(n14022), .ZN(n2866) );
  INV_X1 U6344 ( .A(RD2), .ZN(n16074) );
  INV_X1 U6345 ( .A(RD1), .ZN(n16073) );
  INV_X1 U6346 ( .A(WR), .ZN(n16075) );
  INV_X1 U6347 ( .A(DATAIN[28]), .ZN(n16079) );
  INV_X1 U6348 ( .A(DATAIN[29]), .ZN(n16078) );
  INV_X1 U6349 ( .A(DATAIN[30]), .ZN(n16077) );
  INV_X1 U6350 ( .A(DATAIN[31]), .ZN(n16076) );
  INV_X1 U6351 ( .A(DATAIN[0]), .ZN(n16107) );
  INV_X1 U6352 ( .A(DATAIN[1]), .ZN(n16106) );
  INV_X1 U6353 ( .A(DATAIN[2]), .ZN(n16105) );
  INV_X1 U6354 ( .A(DATAIN[3]), .ZN(n16104) );
  INV_X1 U6355 ( .A(DATAIN[4]), .ZN(n16103) );
  INV_X1 U6356 ( .A(DATAIN[5]), .ZN(n16102) );
  INV_X1 U6357 ( .A(DATAIN[6]), .ZN(n16101) );
  INV_X1 U6358 ( .A(DATAIN[7]), .ZN(n16100) );
  INV_X1 U6359 ( .A(DATAIN[8]), .ZN(n16099) );
  INV_X1 U6360 ( .A(DATAIN[9]), .ZN(n16098) );
  INV_X1 U6361 ( .A(DATAIN[10]), .ZN(n16097) );
  INV_X1 U6362 ( .A(DATAIN[11]), .ZN(n16096) );
  INV_X1 U6363 ( .A(DATAIN[12]), .ZN(n16095) );
  INV_X1 U6364 ( .A(DATAIN[13]), .ZN(n16094) );
  INV_X1 U6365 ( .A(DATAIN[14]), .ZN(n16093) );
  INV_X1 U6366 ( .A(DATAIN[15]), .ZN(n16092) );
  INV_X1 U6367 ( .A(DATAIN[16]), .ZN(n16091) );
  INV_X1 U6368 ( .A(DATAIN[17]), .ZN(n16090) );
  INV_X1 U6369 ( .A(DATAIN[18]), .ZN(n16089) );
  INV_X1 U6370 ( .A(DATAIN[19]), .ZN(n16088) );
  INV_X1 U6371 ( .A(DATAIN[20]), .ZN(n16087) );
  INV_X1 U6372 ( .A(DATAIN[21]), .ZN(n16086) );
  INV_X1 U6373 ( .A(DATAIN[22]), .ZN(n16085) );
  INV_X1 U6374 ( .A(DATAIN[23]), .ZN(n16084) );
  INV_X1 U6375 ( .A(DATAIN[24]), .ZN(n16083) );
  INV_X1 U6376 ( .A(DATAIN[25]), .ZN(n16082) );
  INV_X1 U6377 ( .A(DATAIN[26]), .ZN(n16081) );
  INV_X1 U6378 ( .A(DATAIN[27]), .ZN(n16080) );
  NOR3_X4 U6379 ( .A1(n16060), .A2(ADD_WR[6]), .A3(n16059), .ZN(n2982) );
  NOR3_X4 U6380 ( .A1(ADD_WR[4]), .A2(ADD_WR[6]), .A3(n16059), .ZN(n2949) );
  NOR3_X4 U6381 ( .A1(ADD_WR[5]), .A2(ADD_WR[6]), .A3(n16060), .ZN(n2916) );
  NOR3_X4 U6382 ( .A1(ADD_WR[5]), .A2(ADD_WR[6]), .A3(ADD_WR[4]), .ZN(n2868)
         );
  CLKBUF_X1 U6383 ( .A(n4325), .Z(n13149) );
  CLKBUF_X1 U6384 ( .A(n3041), .Z(n13377) );
  CLKBUF_X1 U6385 ( .A(n2865), .Z(n13829) );
  CLKBUF_X1 U6386 ( .A(n2864), .Z(n13835) );
  CLKBUF_X1 U6387 ( .A(n2863), .Z(n13841) );
  CLKBUF_X1 U6388 ( .A(n2862), .Z(n13847) );
  CLKBUF_X1 U6389 ( .A(n2861), .Z(n13853) );
  CLKBUF_X1 U6390 ( .A(n2860), .Z(n13859) );
  CLKBUF_X1 U6391 ( .A(n2859), .Z(n13865) );
  CLKBUF_X1 U6392 ( .A(n2858), .Z(n13871) );
  CLKBUF_X1 U6393 ( .A(n2857), .Z(n13877) );
  CLKBUF_X1 U6394 ( .A(n2856), .Z(n13883) );
  CLKBUF_X1 U6395 ( .A(n2855), .Z(n13889) );
  CLKBUF_X1 U6396 ( .A(n2854), .Z(n13895) );
  CLKBUF_X1 U6397 ( .A(n2853), .Z(n13901) );
  CLKBUF_X1 U6398 ( .A(n2852), .Z(n13907) );
  CLKBUF_X1 U6399 ( .A(n2851), .Z(n13913) );
  CLKBUF_X1 U6400 ( .A(n2850), .Z(n13919) );
  CLKBUF_X1 U6401 ( .A(n2849), .Z(n13925) );
  CLKBUF_X1 U6402 ( .A(n2848), .Z(n13931) );
  CLKBUF_X1 U6403 ( .A(n2847), .Z(n13937) );
  CLKBUF_X1 U6404 ( .A(n2846), .Z(n13943) );
  CLKBUF_X1 U6405 ( .A(n2845), .Z(n13949) );
  CLKBUF_X1 U6406 ( .A(n2844), .Z(n13955) );
  CLKBUF_X1 U6407 ( .A(n2843), .Z(n13961) );
  CLKBUF_X1 U6408 ( .A(n2842), .Z(n13967) );
  CLKBUF_X1 U6409 ( .A(n2841), .Z(n13973) );
  CLKBUF_X1 U6410 ( .A(n2840), .Z(n13979) );
  CLKBUF_X1 U6411 ( .A(n2839), .Z(n13985) );
  CLKBUF_X1 U6412 ( .A(n2838), .Z(n13991) );
  CLKBUF_X1 U6413 ( .A(n2837), .Z(n13997) );
  CLKBUF_X1 U6414 ( .A(n2836), .Z(n14003) );
  CLKBUF_X1 U6415 ( .A(n2835), .Z(n14009) );
  CLKBUF_X1 U6416 ( .A(n2833), .Z(n14018) );
  CLKBUF_X1 U6417 ( .A(ENABLE), .Z(n14027) );
endmodule


module registerFile_TLE ( clk, reset, enable, rd1, rd2, wr1, add_wr, add_rd1, 
        add_rd2, dataIn, dataOut1, dataOut2, fill, spill, call, ret, dataACK, 
        MMUStrobe );
  input [4:0] add_wr;
  input [4:0] add_rd1;
  input [4:0] add_rd2;
  input [31:0] dataIn;
  output [31:0] dataOut1;
  output [31:0] dataOut2;
  input clk, reset, enable, rd1, rd2, wr1, call, ret, MMUStrobe;
  output fill, spill, dataACK;

  wire   [3:0] cwp_s;
  wire   [6:0] add_wr_out_s;
  wire   [6:0] add_rd1_out_s;
  wire   [6:0] add_rd2_out_s;
  tri   [31:0] dataOut1;
  tri   [31:0] dataOut2;

  controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 contrU ( .clk(
        clk), .reset(reset), .enable(enable), .cwpOut(cwp_s), .call(call), 
        .ret(ret), .fill(fill), .spill(spill), .MMUStrobe(MMUStrobe), 
        .dataACK(dataACK) );
  translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 translU ( 
        .clk(clk), .reset(reset), .enable(enable), .rd1(rd1), .rd2(rd2), .wr(
        wr1), .add_wr(add_wr), .add_rd1(add_rd1), .add_rd2(add_rd2), .cwp(
        cwp_s), .add_wr_out(add_wr_out_s), .add_rd1_out(add_rd1_out_s), 
        .add_rd2_out(add_rd2_out_s) );
  physical_RF_NData32_NRegs72_NAddr7 physRF ( .CLK(clk), .RESET(reset), 
        .ENABLE(enable), .RD1(rd1), .RD2(rd2), .WR(wr1), .ADD_WR(add_wr_out_s), 
        .ADD_RD1(add_rd1_out_s), .ADD_RD2(add_rd2_out_s), .DATAIN(dataIn), 
        .OUT1(dataOut1), .OUT2(dataOut2) );
endmodule

