
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5 
   is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5.all;

entity 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
   is

   port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  SUM :
         out std_logic_vector (31 downto 0));

end controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0
   ;

architecture SYN_rpl of 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n2, n_1000, 
      n_1001 : std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => INC_DEC, CI => carry_31_port, CO =>
                           n_1000, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => INC_DEC, CI => carry_30_port, CO =>
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => INC_DEC, CI => carry_29_port, CO =>
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => INC_DEC, CI => carry_28_port, CO =>
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => INC_DEC, CI => carry_27_port, CO =>
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => INC_DEC, CI => carry_26_port, CO =>
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => INC_DEC, CI => carry_25_port, CO =>
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => INC_DEC, CI => carry_24_port, CO =>
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => INC_DEC, CI => carry_23_port, CO =>
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => INC_DEC, CI => carry_22_port, CO =>
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => INC_DEC, CI => carry_21_port, CO =>
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => INC_DEC, CI => carry_20_port, CO =>
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => INC_DEC, CI => carry_19_port, CO =>
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => INC_DEC, CI => carry_18_port, CO =>
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => INC_DEC, CI => carry_17_port, CO =>
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => INC_DEC, CI => carry_16_port, CO =>
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => INC_DEC, CI => carry_15_port, CO =>
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => INC_DEC, CI => carry_14_port, CO =>
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => INC_DEC, CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => INC_DEC, CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => INC_DEC, CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => INC_DEC, CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => INC_DEC, CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => INC_DEC, CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => INC_DEC, CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => INC_DEC, CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => INC_DEC, CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => INC_DEC, CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => INC_DEC, CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => INC_DEC, CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => INC_DEC, CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => INC_DEC, CI => n2, CO => carry_1_port
                           , S => n_1001);
   U1 : INV_X1 port map( A => INC_DEC, ZN => n2);
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5.all;

entity physical_RF_NData32_NRegs72_NAddr7 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (6 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end physical_RF_NData32_NRegs72_NAddr7;

architecture SYN_beh of physical_RF_NData32_NRegs72_NAddr7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
      n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, 
      n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, 
      n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, 
      n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, 
      n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, 
      n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, 
      n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, 
      n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, 
      n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, 
      n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, 
      n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, 
      n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, 
      n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, 
      n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, 
      n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, 
      n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, 
      n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, 
      n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, 
      n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, 
      n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, 
      n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, 
      n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, 
      n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, 
      n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, 
      n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, 
      n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, 
      n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, 
      n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, 
      n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, 
      n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, 
      n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, 
      n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
      n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, 
      n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, 
      n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, 
      n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, 
      n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, 
      n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, 
      n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, 
      n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, 
      n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, 
      n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, 
      n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, 
      n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
      n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, 
      n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, 
      n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, 
      n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
      n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, 
      n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, 
      n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, 
      n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, 
      n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, 
      n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, 
      n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, 
      n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, 
      n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, 
      n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, 
      n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, 
      n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, 
      n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, 
      n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, 
      n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, 
      n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, 
      n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, 
      n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, 
      n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, 
      n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, 
      n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, 
      n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, 
      n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, 
      n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, 
      n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, 
      n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, 
      n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, 
      n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, 
      n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, 
      n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, 
      n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, 
      n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, 
      n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, 
      n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, 
      n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, 
      n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
      n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, 
      n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, 
      n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, 
      n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, 
      n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, 
      n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
      n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, 
      n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, 
      n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, 
      n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, 
      n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, 
      n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, 
      n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, 
      n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
      n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, 
      n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, 
      n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, 
      n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, 
      n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, 
      n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, 
      n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, 
      n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, 
      n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, 
      n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, 
      n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, 
      n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, 
      n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, 
      n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, 
      n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, 
      n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, 
      n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, 
      n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, 
      n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, 
      n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
      n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, 
      n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
      n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
      n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, 
      n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
      n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, 
      n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, 
      n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, 
      n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, 
      n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, 
      n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, 
      n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, 
      n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, 
      n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, 
      n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, 
      n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, 
      n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, 
      n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, 
      n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, 
      n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, 
      n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, 
      n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, 
      n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, 
      n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, 
      n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
      n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, 
      n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, 
      n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
      n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
      n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
      n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, 
      n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, 
      n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, 
      n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
      n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, 
      n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, 
      n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, 
      n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, 
      n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, 
      n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, 
      n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, 
      n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, 
      n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
      n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, 
      n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, 
      n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, 
      n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, 
      n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, 
      n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, 
      n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, 
      n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, 
      n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, 
      n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, 
      n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, 
      n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, 
      n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, 
      n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, 
      n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, 
      n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, 
      n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, 
      n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, 
      n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, 
      n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, 
      n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
      n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, 
      n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, 
      n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, 
      n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
      n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, 
      n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, 
      n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, 
      n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
      n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, 
      n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, 
      n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, 
      n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
      n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, 
      n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, 
      n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, 
      n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, 
      n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, 
      n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, 
      n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, 
      n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, 
      n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, 
      n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, 
      n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, 
      n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, 
      n9976, n9977, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, 
      n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
      n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
      n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
      n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
      n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
      n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, 
      n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
      n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
      n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
      n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, 
      n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
      n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
      n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
      n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, 
      n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
      n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
      n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
      n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
      n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
      n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
      n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
      n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
      n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, 
      n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
      n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
      n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
      n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
      n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, 
      n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
      n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
      n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
      n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
      n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
      n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
      n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
      n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
      n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
      n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
      n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
      n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
      n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
      n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, 
      n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, 
      n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
      n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
      n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
      n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
      n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
      n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
      n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
      n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
      n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
      n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
      n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
      n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
      n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
      n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
      n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
      n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
      n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
      n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
      n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, 
      n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
      n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
      n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
      n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
      n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
      n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
      n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, 
      n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, 
      n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
      n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
      n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, 
      n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
      n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, 
      n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, 
      n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
      n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
      n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, 
      n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, 
      n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, 
      n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, 
      n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
      n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, 
      n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, 
      n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, 
      n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
      n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
      n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, 
      n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, 
      n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, 
      n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, 
      n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, 
      n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, 
      n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, 
      n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
      n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, 
      n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, 
      n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, 
      n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, 
      n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, 
      n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, 
      n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, 
      n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, 
      n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, 
      n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, 
      n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, 
      n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
      n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, 
      n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, 
      n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, 
      n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
      n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, 
      n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, 
      n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
      n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, 
      n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, 
      n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
      n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, 
      n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, 
      n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, 
      n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, 
      n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, 
      n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, 
      n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, 
      n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
      n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, 
      n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, 
      n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, 
      n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, 
      n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
      n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, 
      n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, 
      n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, 
      n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, 
      n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, 
      n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
      n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
      n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
      n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, 
      n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, 
      n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, 
      n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, 
      n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, 
      n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, 
      n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
      n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
      n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
      n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
      n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, 
      n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
      n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, 
      n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
      n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, 
      n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
      n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, 
      n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
      n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, 
      n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, 
      n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, 
      n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, 
      n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, 
      n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
      n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, 
      n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
      n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, 
      n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, 
      n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, 
      n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, 
      n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, 
      n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
      n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, 
      n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, 
      n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, 
      n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, 
      n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, 
      n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, 
      n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, 
      n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, 
      n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, 
      n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, 
      n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, 
      n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, 
      n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, 
      n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, 
      n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
      n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, 
      n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, 
      n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, 
      n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, 
      n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
      n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, 
      n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, 
      n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, 
      n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, 
      n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, 
      n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
      n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
      n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
      n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
      n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, 
      n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, 
      n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, 
      n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, 
      n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, 
      n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
      n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
      n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, 
      n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, 
      n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, 
      n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
      n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, 
      n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, 
      n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, 
      n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
      n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, 
      n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, 
      n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, 
      n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
      n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, 
      n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, 
      n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, 
      n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, 
      n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, 
      n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, 
      n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, 
      n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, 
      n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, 
      n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, 
      n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, 
      n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, 
      n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, 
      n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, 
      n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, 
      n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, 
      n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, 
      n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, 
      n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, 
      n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, 
      n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, 
      n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, 
      n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, 
      n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, 
      n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, 
      n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, 
      n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, 
      n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, 
      n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, 
      n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
      n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
      n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, 
      n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, 
      n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, 
      n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, 
      n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, 
      n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, 
      n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, 
      n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
      n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, 
      n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, 
      n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, 
      n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, 
      n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, 
      n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, 
      n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
      n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, 
      n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, 
      n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, 
      n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, 
      n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, 
      n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, 
      n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, 
      n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, 
      n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, 
      n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, 
      n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, 
      n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, 
      n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, 
      n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, 
      n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, 
      n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, 
      n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, 
      n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, 
      n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, 
      n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, 
      n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, 
      n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, 
      n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, 
      n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, 
      n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, 
      n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, 
      n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, 
      n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, 
      n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, 
      n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, 
      n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, 
      n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, 
      n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, 
      n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, 
      n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, 
      n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, 
      n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, 
      n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, 
      n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, 
      n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, 
      n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, 
      n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, 
      n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, 
      n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, 
      n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, 
      n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, 
      n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, 
      n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, 
      n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, 
      n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, 
      n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, 
      n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, 
      n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, 
      n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, 
      n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, 
      n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, 
      n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, 
      n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, 
      n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, 
      n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, 
      n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, 
      n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, 
      n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, 
      n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, 
      n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, 
      n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, 
      n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, 
      n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, 
      n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, 
      n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, 
      n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, 
      n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, 
      n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, 
      n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, 
      n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, 
      n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, 
      n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, 
      n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, 
      n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, 
      n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, 
      n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, 
      n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, 
      n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, 
      n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, 
      n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, 
      n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, 
      n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, 
      n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, 
      n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, 
      n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, 
      n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, 
      n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, 
      n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, 
      n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, 
      n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, 
      n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, 
      n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, 
      n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, 
      n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, 
      n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, 
      n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, 
      n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, 
      n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, 
      n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, 
      n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, 
      n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, 
      n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, 
      n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, 
      n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, 
      n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, 
      n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, 
      n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, 
      n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, 
      n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, 
      n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, 
      n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, 
      n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, 
      n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, 
      n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, 
      n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, 
      n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, 
      n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, 
      n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, 
      n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, 
      n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, 
      n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, 
      n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, 
      n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, 
      n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, 
      n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, 
      n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, 
      n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, 
      n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, 
      n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, 
      n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, 
      n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, 
      n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, 
      n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, 
      n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, 
      n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, 
      n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, 
      n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, 
      n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, 
      n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, 
      n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, 
      n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, 
      n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, 
      n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, 
      n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, 
      n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, 
      n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, 
      n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, 
      n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, 
      n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, 
      n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, 
      n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, 
      n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, 
      n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, 
      n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, 
      n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, 
      n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, 
      n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, 
      n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, 
      n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, 
      n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, 
      n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, 
      n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, 
      n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, 
      n6781, n6782, n6783, n6784, n6785, n_1002, n_1003, n_1004, n_1005, n_1006
      , n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015,
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n9977, CK => CLK, Q => n6657
                           , QN => n618);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n9976, CK => CLK, Q => n6656
                           , QN => n621);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n9975, CK => CLK, Q => n6655
                           , QN => n624);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n9974, CK => CLK, Q => n6654
                           , QN => n627);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n9973, CK => CLK, Q => n6653
                           , QN => n630);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n9972, CK => CLK, Q => n6652
                           , QN => n633);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n9971, CK => CLK, Q => n6651
                           , QN => n636);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n9970, CK => CLK, Q => n6650
                           , QN => n639);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n9969, CK => CLK, Q => n6649
                           , QN => n642);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n9968, CK => CLK, Q => n6648
                           , QN => n645);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n9967, CK => CLK, Q => n6647
                           , QN => n648);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n9966, CK => CLK, Q => n6646
                           , QN => n651);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n9965, CK => CLK, Q => n6645
                           , QN => n654);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n9964, CK => CLK, Q => n6644
                           , QN => n657);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n9963, CK => CLK, Q => n6643
                           , QN => n660);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n9962, CK => CLK, Q => n6642
                           , QN => n663);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n9961, CK => CLK, Q => n6641
                           , QN => n666);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n9960, CK => CLK, Q => n6640
                           , QN => n669);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n9959, CK => CLK, Q => n6639
                           , QN => n672);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n9958, CK => CLK, Q => n6638
                           , QN => n675);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n9957, CK => CLK, Q => n6637
                           , QN => n678);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n9956, CK => CLK, Q => n6636
                           , QN => n681);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n9955, CK => CLK, Q => n6635,
                           QN => n684);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n9954, CK => CLK, Q => n6634,
                           QN => n687);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n9953, CK => CLK, Q => n6633,
                           QN => n690);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n9952, CK => CLK, Q => n6632,
                           QN => n693);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n9951, CK => CLK, Q => n6631,
                           QN => n696);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n9950, CK => CLK, Q => n6630,
                           QN => n699);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n9949, CK => CLK, Q => n6629,
                           QN => n702);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n9948, CK => CLK, Q => n6628,
                           QN => n705);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n9947, CK => CLK, Q => n6627,
                           QN => n708);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n9946, CK => CLK, Q => n6626,
                           QN => n711);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n9945, CK => CLK, Q => n6625
                           , QN => n194);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n9944, CK => CLK, Q => n6624
                           , QN => n197);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n9943, CK => CLK, Q => n6623
                           , QN => n200);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n9942, CK => CLK, Q => n6622
                           , QN => n203);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n9941, CK => CLK, Q => n6621
                           , QN => n206);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n9940, CK => CLK, Q => n6620
                           , QN => n209);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n9939, CK => CLK, Q => n6619
                           , QN => n212);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n9938, CK => CLK, Q => n6618
                           , QN => n215);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n9937, CK => CLK, Q => n6617
                           , QN => n218);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n9936, CK => CLK, Q => n6616
                           , QN => n221);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n9935, CK => CLK, Q => n6615
                           , QN => n224);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n9934, CK => CLK, Q => n6614
                           , QN => n227);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n9933, CK => CLK, Q => n6613
                           , QN => n230);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n9932, CK => CLK, Q => n6612
                           , QN => n233);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n9931, CK => CLK, Q => n6611
                           , QN => n236);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n9930, CK => CLK, Q => n6610
                           , QN => n239);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n9929, CK => CLK, Q => n6609
                           , QN => n242);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n9928, CK => CLK, Q => n6608
                           , QN => n245);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n9927, CK => CLK, Q => n6607
                           , QN => n248);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n9926, CK => CLK, Q => n6606
                           , QN => n251);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n9925, CK => CLK, Q => n6605
                           , QN => n254);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n9924, CK => CLK, Q => n6604
                           , QN => n257);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n9923, CK => CLK, Q => n6603,
                           QN => n260);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n9922, CK => CLK, Q => n6602,
                           QN => n263);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n9921, CK => CLK, Q => n6601,
                           QN => n266);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n9920, CK => CLK, Q => n6600,
                           QN => n269);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n9919, CK => CLK, Q => n6599,
                           QN => n272);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n9918, CK => CLK, Q => n6598,
                           QN => n275);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n9917, CK => CLK, Q => n6597,
                           QN => n278);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n9916, CK => CLK, Q => n6596,
                           QN => n281);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n9915, CK => CLK, Q => n6595,
                           QN => n284);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n9914, CK => CLK, Q => n6594,
                           QN => n287);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n9913, CK => CLK, Q => n714,
                           QN => n5696);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n9912, CK => CLK, Q => n717,
                           QN => n5686);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n9911, CK => CLK, Q => n720,
                           QN => n5676);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n9910, CK => CLK, Q => n723,
                           QN => n5666);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n9909, CK => CLK, Q => n726,
                           QN => n5656);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n9908, CK => CLK, Q => n729,
                           QN => n5646);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n9907, CK => CLK, Q => n732,
                           QN => n5636);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n9906, CK => CLK, Q => n735,
                           QN => n5626);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n9905, CK => CLK, Q => n738,
                           QN => n5616);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n9904, CK => CLK, Q => n741,
                           QN => n5606);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n9903, CK => CLK, Q => n744,
                           QN => n5596);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n9902, CK => CLK, Q => n747,
                           QN => n5586);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n9901, CK => CLK, Q => n750,
                           QN => n5576);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n9900, CK => CLK, Q => n753,
                           QN => n5566);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n9899, CK => CLK, Q => n756,
                           QN => n5556);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n9898, CK => CLK, Q => n759,
                           QN => n5546);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n9897, CK => CLK, Q => n762,
                           QN => n5536);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n9896, CK => CLK, Q => n765,
                           QN => n5526);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n9895, CK => CLK, Q => n768,
                           QN => n5516);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n9894, CK => CLK, Q => n771,
                           QN => n5506);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n9893, CK => CLK, Q => n774,
                           QN => n5496);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n9892, CK => CLK, Q => n777,
                           QN => n5486);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n9891, CK => CLK, Q => n780, 
                           QN => n5476);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n9890, CK => CLK, Q => n783, 
                           QN => n5466);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n9889, CK => CLK, Q => n786, 
                           QN => n5456);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n9888, CK => CLK, Q => n789, 
                           QN => n5446);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n9887, CK => CLK, Q => n792, 
                           QN => n5436);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n9886, CK => CLK, Q => n795, 
                           QN => n5426);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n9885, CK => CLK, Q => n798, 
                           QN => n5416);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n9884, CK => CLK, Q => n801, 
                           QN => n5406);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n9883, CK => CLK, Q => n804, 
                           QN => n5396);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n9882, CK => CLK, Q => n807, 
                           QN => n5386);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n9881, CK => CLK, Q => n290,
                           QN => n5697);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n9880, CK => CLK, Q => n293,
                           QN => n5687);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n9879, CK => CLK, Q => n296,
                           QN => n5677);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n9878, CK => CLK, Q => n299,
                           QN => n5667);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n9877, CK => CLK, Q => n302,
                           QN => n5657);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n9876, CK => CLK, Q => n305,
                           QN => n5647);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n9875, CK => CLK, Q => n308,
                           QN => n5637);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n9874, CK => CLK, Q => n311,
                           QN => n5627);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n9873, CK => CLK, Q => n314,
                           QN => n5617);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n9872, CK => CLK, Q => n317,
                           QN => n5607);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n9871, CK => CLK, Q => n320,
                           QN => n5597);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n9870, CK => CLK, Q => n323,
                           QN => n5587);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n9869, CK => CLK, Q => n326,
                           QN => n5577);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n9868, CK => CLK, Q => n329,
                           QN => n5567);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n9867, CK => CLK, Q => n332,
                           QN => n5557);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n9866, CK => CLK, Q => n335,
                           QN => n5547);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n9865, CK => CLK, Q => n338,
                           QN => n5537);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n9864, CK => CLK, Q => n341,
                           QN => n5527);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n9863, CK => CLK, Q => n344,
                           QN => n5517);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n9862, CK => CLK, Q => n347,
                           QN => n5507);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n9861, CK => CLK, Q => n350,
                           QN => n5497);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n9860, CK => CLK, Q => n353,
                           QN => n5487);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n9859, CK => CLK, Q => n356, 
                           QN => n5477);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n9858, CK => CLK, Q => n359, 
                           QN => n5467);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n9857, CK => CLK, Q => n362, 
                           QN => n5457);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n9856, CK => CLK, Q => n365, 
                           QN => n5447);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n9855, CK => CLK, Q => n368, 
                           QN => n5437);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n9854, CK => CLK, Q => n371, 
                           QN => n5427);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n9853, CK => CLK, Q => n374, 
                           QN => n5417);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n9852, CK => CLK, Q => n377, 
                           QN => n5407);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n9851, CK => CLK, Q => n380, 
                           QN => n5397);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n9850, CK => CLK, Q => n383, 
                           QN => n5387);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n9849, CK => CLK, Q => n6593
                           , QN => n809);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n9848, CK => CLK, Q => n6592
                           , QN => n810);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n9847, CK => CLK, Q => n6591
                           , QN => n811);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n9846, CK => CLK, Q => n6590
                           , QN => n812);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n9845, CK => CLK, Q => n6589
                           , QN => n813);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n9844, CK => CLK, Q => n6588
                           , QN => n814);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n9843, CK => CLK, Q => n6587
                           , QN => n815);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n9842, CK => CLK, Q => n6586
                           , QN => n816);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n9841, CK => CLK, Q => n6585
                           , QN => n817);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n9840, CK => CLK, Q => n6584
                           , QN => n818);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n9839, CK => CLK, Q => n6583
                           , QN => n819);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n9838, CK => CLK, Q => n6582
                           , QN => n820);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n9837, CK => CLK, Q => n6581
                           , QN => n821);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n9836, CK => CLK, Q => n6580
                           , QN => n822);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n9835, CK => CLK, Q => n6579
                           , QN => n823);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n9834, CK => CLK, Q => n6578
                           , QN => n824);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n9833, CK => CLK, Q => n6577
                           , QN => n825);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n9832, CK => CLK, Q => n6576
                           , QN => n826);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n9831, CK => CLK, Q => n6575
                           , QN => n827);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n9830, CK => CLK, Q => n6574
                           , QN => n828);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n9829, CK => CLK, Q => n6573
                           , QN => n829);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n9828, CK => CLK, Q => n6572
                           , QN => n830);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n9827, CK => CLK, Q => n6571,
                           QN => n831);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n9826, CK => CLK, Q => n6570,
                           QN => n832);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n9825, CK => CLK, Q => n6569,
                           QN => n833);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n9824, CK => CLK, Q => n6568,
                           QN => n834);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n9823, CK => CLK, Q => n6567,
                           QN => n835);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n9822, CK => CLK, Q => n6566,
                           QN => n836);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n9821, CK => CLK, Q => n6565,
                           QN => n837);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n9820, CK => CLK, Q => n6564,
                           QN => n838);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n9819, CK => CLK, Q => n6563,
                           QN => n839);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n9818, CK => CLK, Q => n6562,
                           QN => n840);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n9817, CK => CLK, Q => n6561
                           , QN => n1161);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n9816, CK => CLK, Q => n6560
                           , QN => n1162);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n9815, CK => CLK, Q => n6559
                           , QN => n1163);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n9814, CK => CLK, Q => n6558
                           , QN => n1164);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n9813, CK => CLK, Q => n6557
                           , QN => n1165);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n9812, CK => CLK, Q => n6556
                           , QN => n1166);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n9811, CK => CLK, Q => n6555
                           , QN => n1167);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n9810, CK => CLK, Q => n6554
                           , QN => n1168);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n9809, CK => CLK, Q => n6553
                           , QN => n1169);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n9808, CK => CLK, Q => n6552
                           , QN => n1170);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n9807, CK => CLK, Q => n6551
                           , QN => n1171);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n9806, CK => CLK, Q => n6550
                           , QN => n1172);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n9805, CK => CLK, Q => n6549
                           , QN => n1173);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n9804, CK => CLK, Q => n6548
                           , QN => n1174);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n9803, CK => CLK, Q => n6547
                           , QN => n1175);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n9802, CK => CLK, Q => n6546
                           , QN => n1176);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n9801, CK => CLK, Q => n6545
                           , QN => n1177);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n9800, CK => CLK, Q => n6544
                           , QN => n1178);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n9799, CK => CLK, Q => n6543
                           , QN => n1179);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n9798, CK => CLK, Q => n6542
                           , QN => n1180);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n9797, CK => CLK, Q => n6541
                           , QN => n1181);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n9796, CK => CLK, Q => n6540
                           , QN => n1182);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n9795, CK => CLK, Q => n6539,
                           QN => n1183);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n9794, CK => CLK, Q => n6538,
                           QN => n1184);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n9793, CK => CLK, Q => n6537,
                           QN => n1185);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n9792, CK => CLK, Q => n6536,
                           QN => n1186);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n9791, CK => CLK, Q => n6535,
                           QN => n1187);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n9790, CK => CLK, Q => n6534,
                           QN => n1188);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n9789, CK => CLK, Q => n6533,
                           QN => n1189);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n9788, CK => CLK, Q => n6532,
                           QN => n1190);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n9787, CK => CLK, Q => n6531,
                           QN => n1191);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n9786, CK => CLK, Q => n6530,
                           QN => n1192);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n9785, CK => CLK, Q => 
                           n_1002, QN => n5377);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n9784, CK => CLK, Q => 
                           n_1003, QN => n5376);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n9783, CK => CLK, Q => 
                           n_1004, QN => n5375);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n9782, CK => CLK, Q => 
                           n_1005, QN => n5374);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n9781, CK => CLK, Q => 
                           n_1006, QN => n5373);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n9780, CK => CLK, Q => 
                           n_1007, QN => n5372);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n9779, CK => CLK, Q => 
                           n_1008, QN => n5371);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n9778, CK => CLK, Q => 
                           n_1009, QN => n5370);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n9777, CK => CLK, Q => 
                           n_1010, QN => n5369);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n9776, CK => CLK, Q => 
                           n_1011, QN => n5368);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n9775, CK => CLK, Q => 
                           n_1012, QN => n5367);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n9774, CK => CLK, Q => 
                           n_1013, QN => n5366);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n9773, CK => CLK, Q => 
                           n_1014, QN => n5365);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n9772, CK => CLK, Q => 
                           n_1015, QN => n5364);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n9771, CK => CLK, Q => 
                           n_1016, QN => n5363);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n9770, CK => CLK, Q => 
                           n_1017, QN => n5362);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n9769, CK => CLK, Q => 
                           n_1018, QN => n5361);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n9768, CK => CLK, Q => 
                           n_1019, QN => n5360);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n9767, CK => CLK, Q => 
                           n_1020, QN => n5359);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n9766, CK => CLK, Q => 
                           n_1021, QN => n5358);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n9765, CK => CLK, Q => 
                           n_1022, QN => n5357);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n9764, CK => CLK, Q => 
                           n_1023, QN => n5356);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n9763, CK => CLK, Q => n_1024
                           , QN => n5355);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n9762, CK => CLK, Q => n_1025
                           , QN => n5354);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n9761, CK => CLK, Q => n_1026
                           , QN => n5353);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n9760, CK => CLK, Q => n_1027
                           , QN => n5352);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n9759, CK => CLK, Q => n_1028
                           , QN => n5351);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n9758, CK => CLK, Q => n_1029
                           , QN => n5350);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n9757, CK => CLK, Q => n_1030
                           , QN => n5349);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n9756, CK => CLK, Q => n_1031
                           , QN => n5348);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n9755, CK => CLK, Q => n_1032
                           , QN => n5347);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n9754, CK => CLK, Q => n_1033
                           , QN => n5346);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n9753, CK => CLK, Q => 
                           n_1034, QN => n5345);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n9752, CK => CLK, Q => 
                           n_1035, QN => n5344);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n9751, CK => CLK, Q => 
                           n_1036, QN => n5343);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n9750, CK => CLK, Q => 
                           n_1037, QN => n5342);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n9749, CK => CLK, Q => 
                           n_1038, QN => n5341);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n9748, CK => CLK, Q => 
                           n_1039, QN => n5340);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n9747, CK => CLK, Q => 
                           n_1040, QN => n5339);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n9746, CK => CLK, Q => 
                           n_1041, QN => n5338);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n9745, CK => CLK, Q => 
                           n_1042, QN => n5337);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n9744, CK => CLK, Q => 
                           n_1043, QN => n5336);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n9743, CK => CLK, Q => 
                           n_1044, QN => n5335);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n9742, CK => CLK, Q => 
                           n_1045, QN => n5334);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n9741, CK => CLK, Q => 
                           n_1046, QN => n5333);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n9740, CK => CLK, Q => 
                           n_1047, QN => n5332);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n9739, CK => CLK, Q => 
                           n_1048, QN => n5331);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n9738, CK => CLK, Q => 
                           n_1049, QN => n5330);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n9737, CK => CLK, Q => 
                           n_1050, QN => n5329);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n9736, CK => CLK, Q => 
                           n_1051, QN => n5328);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n9735, CK => CLK, Q => 
                           n_1052, QN => n5327);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n9734, CK => CLK, Q => 
                           n_1053, QN => n5326);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n9733, CK => CLK, Q => 
                           n_1054, QN => n5325);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n9732, CK => CLK, Q => 
                           n_1055, QN => n5324);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n9731, CK => CLK, Q => n_1056
                           , QN => n5323);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n9730, CK => CLK, Q => n_1057
                           , QN => n5322);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n9729, CK => CLK, Q => n_1058
                           , QN => n5321);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n9728, CK => CLK, Q => n_1059
                           , QN => n5320);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n9727, CK => CLK, Q => n_1060
                           , QN => n5319);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n9726, CK => CLK, Q => n_1061
                           , QN => n5318);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n9725, CK => CLK, Q => n_1062
                           , QN => n5317);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n9724, CK => CLK, Q => n_1063
                           , QN => n5316);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n9723, CK => CLK, Q => n_1064
                           , QN => n5315);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n9722, CK => CLK, Q => n_1065
                           , QN => n5314);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n9721, CK => CLK, Q => 
                           n_1066, QN => n5313);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n9720, CK => CLK, Q => 
                           n_1067, QN => n5312);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n9719, CK => CLK, Q => 
                           n_1068, QN => n5311);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n9718, CK => CLK, Q => 
                           n_1069, QN => n5310);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n9717, CK => CLK, Q => 
                           n_1070, QN => n5309);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n9716, CK => CLK, Q => 
                           n_1071, QN => n5308);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n9715, CK => CLK, Q => 
                           n_1072, QN => n5307);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n9714, CK => CLK, Q => 
                           n_1073, QN => n5306);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n9713, CK => CLK, Q => 
                           n_1074, QN => n5305);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n9712, CK => CLK, Q => 
                           n_1075, QN => n5304);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n9711, CK => CLK, Q => 
                           n_1076, QN => n5303);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n9710, CK => CLK, Q => 
                           n_1077, QN => n5302);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n9709, CK => CLK, Q => 
                           n_1078, QN => n5301);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n9708, CK => CLK, Q => 
                           n_1079, QN => n5300);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n9707, CK => CLK, Q => 
                           n_1080, QN => n5299);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n9706, CK => CLK, Q => 
                           n_1081, QN => n5298);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n9705, CK => CLK, Q => 
                           n_1082, QN => n5297);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n9704, CK => CLK, Q => 
                           n_1083, QN => n5296);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n9703, CK => CLK, Q => 
                           n_1084, QN => n5295);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n9702, CK => CLK, Q => 
                           n_1085, QN => n5294);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n9701, CK => CLK, Q => 
                           n_1086, QN => n5293);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n9700, CK => CLK, Q => 
                           n_1087, QN => n5292);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n9699, CK => CLK, Q => n_1088
                           , QN => n5291);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n9698, CK => CLK, Q => n_1089
                           , QN => n5290);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n9697, CK => CLK, Q => n_1090
                           , QN => n5289);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n9696, CK => CLK, Q => n_1091
                           , QN => n5288);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n9695, CK => CLK, Q => n_1092
                           , QN => n5287);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n9694, CK => CLK, Q => n_1093
                           , QN => n5286);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n9693, CK => CLK, Q => n_1094
                           , QN => n5285);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n9692, CK => CLK, Q => n_1095
                           , QN => n5284);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n9691, CK => CLK, Q => n_1096
                           , QN => n5283);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n9690, CK => CLK, Q => n_1097
                           , QN => n5282);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n9689, CK => CLK, Q => n6529
                           , QN => n617);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n9688, CK => CLK, Q => n6528
                           , QN => n620);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n9687, CK => CLK, Q => n6527
                           , QN => n623);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n9686, CK => CLK, Q => n6526
                           , QN => n626);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n9685, CK => CLK, Q => n6525
                           , QN => n629);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n9684, CK => CLK, Q => n6524
                           , QN => n632);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n9683, CK => CLK, Q => n6523
                           , QN => n635);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n9682, CK => CLK, Q => n6522
                           , QN => n638);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n9681, CK => CLK, Q => n6521
                           , QN => n641);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n9680, CK => CLK, Q => n6520
                           , QN => n644);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n9679, CK => CLK, Q => n6519
                           , QN => n647);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n9678, CK => CLK, Q => n6518
                           , QN => n650);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n9677, CK => CLK, Q => n6517
                           , QN => n653);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n9676, CK => CLK, Q => n6516
                           , QN => n656);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n9675, CK => CLK, Q => n6515
                           , QN => n659);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n9674, CK => CLK, Q => n6514
                           , QN => n662);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n9673, CK => CLK, Q => n6513
                           , QN => n665);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n9672, CK => CLK, Q => n6512
                           , QN => n668);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n9671, CK => CLK, Q => n6511
                           , QN => n671);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n9670, CK => CLK, Q => n6510
                           , QN => n674);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n9669, CK => CLK, Q => n6509
                           , QN => n677);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n9668, CK => CLK, Q => n6508
                           , QN => n680);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n9667, CK => CLK, Q => n6507,
                           QN => n683);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n9666, CK => CLK, Q => n6506,
                           QN => n686);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n9665, CK => CLK, Q => n6505,
                           QN => n689);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n9664, CK => CLK, Q => n6504,
                           QN => n692);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n9663, CK => CLK, Q => n6503,
                           QN => n695);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n9662, CK => CLK, Q => n6502,
                           QN => n698);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n9661, CK => CLK, Q => n6501,
                           QN => n701);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n9660, CK => CLK, Q => n6500,
                           QN => n704);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n9659, CK => CLK, Q => n6499,
                           QN => n707);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n9658, CK => CLK, Q => n6498,
                           QN => n710);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n9657, CK => CLK, Q => 
                           n6497, QN => n193);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n9656, CK => CLK, Q => 
                           n6496, QN => n196);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n9655, CK => CLK, Q => 
                           n6495, QN => n199);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n9654, CK => CLK, Q => 
                           n6494, QN => n202);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n9653, CK => CLK, Q => 
                           n6493, QN => n205);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n9652, CK => CLK, Q => 
                           n6492, QN => n208);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n9651, CK => CLK, Q => 
                           n6491, QN => n211);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n9650, CK => CLK, Q => 
                           n6490, QN => n214);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n9649, CK => CLK, Q => 
                           n6489, QN => n217);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n9648, CK => CLK, Q => 
                           n6488, QN => n220);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n9647, CK => CLK, Q => 
                           n6487, QN => n223);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n9646, CK => CLK, Q => 
                           n6486, QN => n226);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n9645, CK => CLK, Q => 
                           n6485, QN => n229);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n9644, CK => CLK, Q => 
                           n6484, QN => n232);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n9643, CK => CLK, Q => 
                           n6483, QN => n235);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n9642, CK => CLK, Q => 
                           n6482, QN => n238);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n9641, CK => CLK, Q => 
                           n6481, QN => n241);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n9640, CK => CLK, Q => 
                           n6480, QN => n244);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n9639, CK => CLK, Q => 
                           n6479, QN => n247);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n9638, CK => CLK, Q => 
                           n6478, QN => n250);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n9637, CK => CLK, Q => 
                           n6477, QN => n253);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n9636, CK => CLK, Q => 
                           n6476, QN => n256);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n9635, CK => CLK, Q => n6475
                           , QN => n259);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n9634, CK => CLK, Q => n6474
                           , QN => n262);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n9633, CK => CLK, Q => n6473
                           , QN => n265);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n9632, CK => CLK, Q => n6472
                           , QN => n268);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n9631, CK => CLK, Q => n6471
                           , QN => n271);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n9630, CK => CLK, Q => n6470
                           , QN => n274);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n9629, CK => CLK, Q => n6469
                           , QN => n277);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n9628, CK => CLK, Q => n6468
                           , QN => n280);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n9627, CK => CLK, Q => n6467
                           , QN => n283);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n9626, CK => CLK, Q => n6466
                           , QN => n286);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n9625, CK => CLK, Q => n713
                           , QN => n5694);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n9624, CK => CLK, Q => n716
                           , QN => n5684);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n9623, CK => CLK, Q => n719
                           , QN => n5674);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n9622, CK => CLK, Q => n722
                           , QN => n5664);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n9621, CK => CLK, Q => n725
                           , QN => n5654);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n9620, CK => CLK, Q => n728
                           , QN => n5644);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n9619, CK => CLK, Q => n731
                           , QN => n5634);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n9618, CK => CLK, Q => n734
                           , QN => n5624);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n9617, CK => CLK, Q => n737
                           , QN => n5614);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n9616, CK => CLK, Q => n740
                           , QN => n5604);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n9615, CK => CLK, Q => n743
                           , QN => n5594);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n9614, CK => CLK, Q => n746
                           , QN => n5584);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n9613, CK => CLK, Q => n749
                           , QN => n5574);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n9612, CK => CLK, Q => n752
                           , QN => n5564);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n9611, CK => CLK, Q => n755
                           , QN => n5554);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n9610, CK => CLK, Q => n758
                           , QN => n5544);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n9609, CK => CLK, Q => n761
                           , QN => n5534);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n9608, CK => CLK, Q => n764
                           , QN => n5524);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n9607, CK => CLK, Q => n767
                           , QN => n5514);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n9606, CK => CLK, Q => n770
                           , QN => n5504);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n9605, CK => CLK, Q => n773
                           , QN => n5494);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n9604, CK => CLK, Q => n776
                           , QN => n5484);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n9603, CK => CLK, Q => n779,
                           QN => n5474);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n9602, CK => CLK, Q => n782,
                           QN => n5464);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n9601, CK => CLK, Q => n785,
                           QN => n5454);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n9600, CK => CLK, Q => n788,
                           QN => n5444);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n9599, CK => CLK, Q => n791,
                           QN => n5434);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n9598, CK => CLK, Q => n794,
                           QN => n5424);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n9597, CK => CLK, Q => n797,
                           QN => n5414);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n9596, CK => CLK, Q => n800,
                           QN => n5404);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n9595, CK => CLK, Q => n803,
                           QN => n5394);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n9594, CK => CLK, Q => n806,
                           QN => n5384);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n9593, CK => CLK, Q => n289
                           , QN => n5695);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n9592, CK => CLK, Q => n292
                           , QN => n5685);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n9591, CK => CLK, Q => n295
                           , QN => n5675);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n9590, CK => CLK, Q => n298
                           , QN => n5665);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n9589, CK => CLK, Q => n301
                           , QN => n5655);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n9588, CK => CLK, Q => n304
                           , QN => n5645);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n9587, CK => CLK, Q => n307
                           , QN => n5635);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n9586, CK => CLK, Q => n310
                           , QN => n5625);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n9585, CK => CLK, Q => n313
                           , QN => n5615);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n9584, CK => CLK, Q => n316
                           , QN => n5605);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n9583, CK => CLK, Q => n319
                           , QN => n5595);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n9582, CK => CLK, Q => n322
                           , QN => n5585);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n9581, CK => CLK, Q => n325
                           , QN => n5575);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n9580, CK => CLK, Q => n328
                           , QN => n5565);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n9579, CK => CLK, Q => n331
                           , QN => n5555);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n9578, CK => CLK, Q => n334
                           , QN => n5545);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n9577, CK => CLK, Q => n337
                           , QN => n5535);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n9576, CK => CLK, Q => n340
                           , QN => n5525);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n9575, CK => CLK, Q => n343
                           , QN => n5515);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n9574, CK => CLK, Q => n346
                           , QN => n5505);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n9573, CK => CLK, Q => n349
                           , QN => n5495);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n9572, CK => CLK, Q => n352
                           , QN => n5485);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n9571, CK => CLK, Q => n355,
                           QN => n5475);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n9570, CK => CLK, Q => n358,
                           QN => n5465);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n9569, CK => CLK, Q => n361,
                           QN => n5455);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n9568, CK => CLK, Q => n364,
                           QN => n5445);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n9567, CK => CLK, Q => n367,
                           QN => n5435);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n9566, CK => CLK, Q => n370,
                           QN => n5425);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n9565, CK => CLK, Q => n373,
                           QN => n5415);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n9564, CK => CLK, Q => n376,
                           QN => n5405);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n9563, CK => CLK, Q => n379,
                           QN => n5395);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n9562, CK => CLK, Q => n382,
                           QN => n5385);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n9561, CK => CLK, Q => 
                           n6465, QN => n841);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n9560, CK => CLK, Q => 
                           n6464, QN => n842);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n9559, CK => CLK, Q => 
                           n6463, QN => n843);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n9558, CK => CLK, Q => 
                           n6462, QN => n844);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n9557, CK => CLK, Q => 
                           n6461, QN => n845);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n9556, CK => CLK, Q => 
                           n6460, QN => n846);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n9555, CK => CLK, Q => 
                           n6459, QN => n847);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n9554, CK => CLK, Q => 
                           n6458, QN => n848);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n9553, CK => CLK, Q => 
                           n6457, QN => n849);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n9552, CK => CLK, Q => 
                           n6456, QN => n850);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n9551, CK => CLK, Q => 
                           n6455, QN => n851);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n9550, CK => CLK, Q => 
                           n6454, QN => n852);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n9549, CK => CLK, Q => 
                           n6453, QN => n853);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n9548, CK => CLK, Q => 
                           n6452, QN => n854);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n9547, CK => CLK, Q => 
                           n6451, QN => n855);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n9546, CK => CLK, Q => 
                           n6450, QN => n856);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n9545, CK => CLK, Q => 
                           n6449, QN => n857);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n9544, CK => CLK, Q => 
                           n6448, QN => n858);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n9543, CK => CLK, Q => 
                           n6447, QN => n859);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n9542, CK => CLK, Q => 
                           n6446, QN => n860);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n9541, CK => CLK, Q => 
                           n6445, QN => n861);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n9540, CK => CLK, Q => 
                           n6444, QN => n862);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n9539, CK => CLK, Q => n6443
                           , QN => n863);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n9538, CK => CLK, Q => n6442
                           , QN => n864);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n9537, CK => CLK, Q => n6441
                           , QN => n865);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n9536, CK => CLK, Q => n6440
                           , QN => n866);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n9535, CK => CLK, Q => n6439
                           , QN => n867);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n9534, CK => CLK, Q => n6438
                           , QN => n868);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n9533, CK => CLK, Q => n6437
                           , QN => n869);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n9532, CK => CLK, Q => n6436
                           , QN => n870);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n9531, CK => CLK, Q => n6435
                           , QN => n871);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n9530, CK => CLK, Q => n6434
                           , QN => n872);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n9529, CK => CLK, Q => 
                           n6433, QN => n1193);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n9528, CK => CLK, Q => 
                           n6432, QN => n1194);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n9527, CK => CLK, Q => 
                           n6431, QN => n1195);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n9526, CK => CLK, Q => 
                           n6430, QN => n1196);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n9525, CK => CLK, Q => 
                           n6429, QN => n1197);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n9524, CK => CLK, Q => 
                           n6428, QN => n1198);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n9523, CK => CLK, Q => 
                           n6427, QN => n1199);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n9522, CK => CLK, Q => 
                           n6426, QN => n1200);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n9521, CK => CLK, Q => 
                           n6425, QN => n1201);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n9520, CK => CLK, Q => 
                           n6424, QN => n1202);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n9519, CK => CLK, Q => 
                           n6423, QN => n1203);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n9518, CK => CLK, Q => 
                           n6422, QN => n1204);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n9517, CK => CLK, Q => 
                           n6421, QN => n1205);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n9516, CK => CLK, Q => 
                           n6420, QN => n1206);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n9515, CK => CLK, Q => 
                           n6419, QN => n1207);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n9514, CK => CLK, Q => 
                           n6418, QN => n1208);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n9513, CK => CLK, Q => 
                           n6417, QN => n1209);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n9512, CK => CLK, Q => 
                           n6416, QN => n1210);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n9511, CK => CLK, Q => 
                           n6415, QN => n1211);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n9510, CK => CLK, Q => 
                           n6414, QN => n1212);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n9509, CK => CLK, Q => 
                           n6413, QN => n1213);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n9508, CK => CLK, Q => 
                           n6412, QN => n1214);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n9507, CK => CLK, Q => n6411
                           , QN => n1215);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n9506, CK => CLK, Q => n6410
                           , QN => n1216);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n9505, CK => CLK, Q => n6409
                           , QN => n1217);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n9504, CK => CLK, Q => n6408
                           , QN => n1218);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n9503, CK => CLK, Q => n6407
                           , QN => n1219);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n9502, CK => CLK, Q => n6406
                           , QN => n1220);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n9501, CK => CLK, Q => n6405
                           , QN => n1221);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n9500, CK => CLK, Q => n6404
                           , QN => n1222);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n9499, CK => CLK, Q => n6403
                           , QN => n1223);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n9498, CK => CLK, Q => n6402
                           , QN => n1224);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n9497, CK => CLK, Q => 
                           n_1098, QN => n5281);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n9496, CK => CLK, Q => 
                           n_1099, QN => n5280);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n9495, CK => CLK, Q => 
                           n_1100, QN => n5279);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n9494, CK => CLK, Q => 
                           n_1101, QN => n5278);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n9493, CK => CLK, Q => 
                           n_1102, QN => n5277);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n9492, CK => CLK, Q => 
                           n_1103, QN => n5276);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n9491, CK => CLK, Q => 
                           n_1104, QN => n5275);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n9490, CK => CLK, Q => 
                           n_1105, QN => n5274);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n9489, CK => CLK, Q => 
                           n_1106, QN => n5273);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n9488, CK => CLK, Q => 
                           n_1107, QN => n5272);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n9487, CK => CLK, Q => 
                           n_1108, QN => n5271);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n9486, CK => CLK, Q => 
                           n_1109, QN => n5270);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n9485, CK => CLK, Q => 
                           n_1110, QN => n5269);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n9484, CK => CLK, Q => 
                           n_1111, QN => n5268);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n9483, CK => CLK, Q => 
                           n_1112, QN => n5267);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n9482, CK => CLK, Q => 
                           n_1113, QN => n5266);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n9481, CK => CLK, Q => 
                           n_1114, QN => n5265);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n9480, CK => CLK, Q => 
                           n_1115, QN => n5264);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n9479, CK => CLK, Q => 
                           n_1116, QN => n5263);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n9478, CK => CLK, Q => 
                           n_1117, QN => n5262);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n9477, CK => CLK, Q => 
                           n_1118, QN => n5261);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n9476, CK => CLK, Q => 
                           n_1119, QN => n5260);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n9475, CK => CLK, Q => 
                           n_1120, QN => n5259);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n9474, CK => CLK, Q => 
                           n_1121, QN => n5258);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n9473, CK => CLK, Q => 
                           n_1122, QN => n5257);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n9472, CK => CLK, Q => 
                           n_1123, QN => n5256);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n9471, CK => CLK, Q => 
                           n_1124, QN => n5255);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n9470, CK => CLK, Q => 
                           n_1125, QN => n5254);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n9469, CK => CLK, Q => 
                           n_1126, QN => n5253);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n9468, CK => CLK, Q => 
                           n_1127, QN => n5252);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n9467, CK => CLK, Q => 
                           n_1128, QN => n5251);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n9466, CK => CLK, Q => 
                           n_1129, QN => n5250);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n9465, CK => CLK, Q => 
                           n_1130, QN => n5249);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n9464, CK => CLK, Q => 
                           n_1131, QN => n5248);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n9463, CK => CLK, Q => 
                           n_1132, QN => n5247);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n9462, CK => CLK, Q => 
                           n_1133, QN => n5246);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n9461, CK => CLK, Q => 
                           n_1134, QN => n5245);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n9460, CK => CLK, Q => 
                           n_1135, QN => n5244);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n9459, CK => CLK, Q => 
                           n_1136, QN => n5243);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n9458, CK => CLK, Q => 
                           n_1137, QN => n5242);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n9457, CK => CLK, Q => 
                           n_1138, QN => n5241);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n9456, CK => CLK, Q => 
                           n_1139, QN => n5240);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n9455, CK => CLK, Q => 
                           n_1140, QN => n5239);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n9454, CK => CLK, Q => 
                           n_1141, QN => n5238);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n9453, CK => CLK, Q => 
                           n_1142, QN => n5237);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n9452, CK => CLK, Q => 
                           n_1143, QN => n5236);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n9451, CK => CLK, Q => 
                           n_1144, QN => n5235);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n9450, CK => CLK, Q => 
                           n_1145, QN => n5234);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n9449, CK => CLK, Q => 
                           n_1146, QN => n5233);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n9448, CK => CLK, Q => 
                           n_1147, QN => n5232);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n9447, CK => CLK, Q => 
                           n_1148, QN => n5231);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n9446, CK => CLK, Q => 
                           n_1149, QN => n5230);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n9445, CK => CLK, Q => 
                           n_1150, QN => n5229);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n9444, CK => CLK, Q => 
                           n_1151, QN => n5228);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n9443, CK => CLK, Q => 
                           n_1152, QN => n5227);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n9442, CK => CLK, Q => 
                           n_1153, QN => n5226);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n9441, CK => CLK, Q => 
                           n_1154, QN => n5225);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n9440, CK => CLK, Q => 
                           n_1155, QN => n5224);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n9439, CK => CLK, Q => 
                           n_1156, QN => n5223);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n9438, CK => CLK, Q => 
                           n_1157, QN => n5222);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n9437, CK => CLK, Q => 
                           n_1158, QN => n5221);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n9436, CK => CLK, Q => 
                           n_1159, QN => n5220);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n9435, CK => CLK, Q => 
                           n_1160, QN => n5219);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n9434, CK => CLK, Q => 
                           n_1161, QN => n5218);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n9433, CK => CLK, Q => 
                           n_1162, QN => n5217);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n9432, CK => CLK, Q => 
                           n_1163, QN => n5216);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n9431, CK => CLK, Q => 
                           n_1164, QN => n5215);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n9430, CK => CLK, Q => 
                           n_1165, QN => n5214);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n9429, CK => CLK, Q => 
                           n_1166, QN => n5213);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n9428, CK => CLK, Q => 
                           n_1167, QN => n5212);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n9427, CK => CLK, Q => 
                           n_1168, QN => n5211);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n9426, CK => CLK, Q => 
                           n_1169, QN => n5210);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n9425, CK => CLK, Q => 
                           n_1170, QN => n5209);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n9424, CK => CLK, Q => 
                           n_1171, QN => n5208);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n9423, CK => CLK, Q => 
                           n_1172, QN => n5207);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n9422, CK => CLK, Q => 
                           n_1173, QN => n5206);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n9421, CK => CLK, Q => 
                           n_1174, QN => n5205);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n9420, CK => CLK, Q => 
                           n_1175, QN => n5204);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n9419, CK => CLK, Q => 
                           n_1176, QN => n5203);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n9418, CK => CLK, Q => 
                           n_1177, QN => n5202);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n9417, CK => CLK, Q => 
                           n_1178, QN => n5201);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n9416, CK => CLK, Q => 
                           n_1179, QN => n5200);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n9415, CK => CLK, Q => 
                           n_1180, QN => n5199);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n9414, CK => CLK, Q => 
                           n_1181, QN => n5198);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n9413, CK => CLK, Q => 
                           n_1182, QN => n5197);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n9412, CK => CLK, Q => 
                           n_1183, QN => n5196);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n9411, CK => CLK, Q => 
                           n_1184, QN => n5195);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n9410, CK => CLK, Q => 
                           n_1185, QN => n5194);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n9409, CK => CLK, Q => 
                           n_1186, QN => n5193);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n9408, CK => CLK, Q => 
                           n_1187, QN => n5192);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n9407, CK => CLK, Q => 
                           n_1188, QN => n5191);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n9406, CK => CLK, Q => 
                           n_1189, QN => n5190);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n9405, CK => CLK, Q => 
                           n_1190, QN => n5189);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n9404, CK => CLK, Q => 
                           n_1191, QN => n5188);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n9403, CK => CLK, Q => 
                           n_1192, QN => n5187);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n9402, CK => CLK, Q => 
                           n_1193, QN => n5186);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n9401, CK => CLK, Q => 
                           n_1194, QN => n457);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n9400, CK => CLK, Q => 
                           n_1195, QN => n459);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n9399, CK => CLK, Q => 
                           n_1196, QN => n461);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n9398, CK => CLK, Q => 
                           n_1197, QN => n463);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n9397, CK => CLK, Q => 
                           n_1198, QN => n465);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n9396, CK => CLK, Q => 
                           n_1199, QN => n467);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n9395, CK => CLK, Q => 
                           n_1200, QN => n469);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n9394, CK => CLK, Q => 
                           n_1201, QN => n471);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n9393, CK => CLK, Q => 
                           n_1202, QN => n473);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n9392, CK => CLK, Q => 
                           n_1203, QN => n475);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n9391, CK => CLK, Q => 
                           n_1204, QN => n477);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n9390, CK => CLK, Q => 
                           n_1205, QN => n479);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n9389, CK => CLK, Q => 
                           n_1206, QN => n481);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n9388, CK => CLK, Q => 
                           n_1207, QN => n483);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n9387, CK => CLK, Q => 
                           n_1208, QN => n485);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n9386, CK => CLK, Q => 
                           n_1209, QN => n487);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n9385, CK => CLK, Q => 
                           n_1210, QN => n489);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n9384, CK => CLK, Q => 
                           n_1211, QN => n491);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n9383, CK => CLK, Q => 
                           n_1212, QN => n493);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n9382, CK => CLK, Q => 
                           n_1213, QN => n495);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n9381, CK => CLK, Q => 
                           n_1214, QN => n497);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n9380, CK => CLK, Q => 
                           n_1215, QN => n499);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n9379, CK => CLK, Q => 
                           n_1216, QN => n501);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n9378, CK => CLK, Q => 
                           n_1217, QN => n503);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n9377, CK => CLK, Q => 
                           n_1218, QN => n505);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n9376, CK => CLK, Q => 
                           n_1219, QN => n507);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n9375, CK => CLK, Q => 
                           n_1220, QN => n509);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n9374, CK => CLK, Q => 
                           n_1221, QN => n511);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n9373, CK => CLK, Q => 
                           n_1222, QN => n513);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n9372, CK => CLK, Q => 
                           n_1223, QN => n515);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n9371, CK => CLK, Q => 
                           n_1224, QN => n517);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n9370, CK => CLK, Q => 
                           n_1225, QN => n519);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n9369, CK => CLK, Q => 
                           n_1226, QN => n1);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n9368, CK => CLK, Q => 
                           n_1227, QN => n3);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n9367, CK => CLK, Q => 
                           n_1228, QN => n5);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n9366, CK => CLK, Q => 
                           n_1229, QN => n7);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n9365, CK => CLK, Q => 
                           n_1230, QN => n9);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n9364, CK => CLK, Q => 
                           n_1231, QN => n11);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n9363, CK => CLK, Q => 
                           n_1232, QN => n13);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n9362, CK => CLK, Q => 
                           n_1233, QN => n15);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n9361, CK => CLK, Q => 
                           n_1234, QN => n17);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n9360, CK => CLK, Q => 
                           n_1235, QN => n19);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n9359, CK => CLK, Q => 
                           n_1236, QN => n21);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n9358, CK => CLK, Q => 
                           n_1237, QN => n23);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n9357, CK => CLK, Q => 
                           n_1238, QN => n25);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n9356, CK => CLK, Q => 
                           n_1239, QN => n27);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n9355, CK => CLK, Q => 
                           n_1240, QN => n29);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n9354, CK => CLK, Q => 
                           n_1241, QN => n31);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n9353, CK => CLK, Q => 
                           n_1242, QN => n33);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n9352, CK => CLK, Q => 
                           n_1243, QN => n35);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n9351, CK => CLK, Q => 
                           n_1244, QN => n37);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n9350, CK => CLK, Q => 
                           n_1245, QN => n39);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n9349, CK => CLK, Q => 
                           n_1246, QN => n41);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n9348, CK => CLK, Q => 
                           n_1247, QN => n43);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n9347, CK => CLK, Q => 
                           n_1248, QN => n45);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n9346, CK => CLK, Q => 
                           n_1249, QN => n47);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n9345, CK => CLK, Q => 
                           n_1250, QN => n49);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n9344, CK => CLK, Q => 
                           n_1251, QN => n51);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n9343, CK => CLK, Q => 
                           n_1252, QN => n53);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n9342, CK => CLK, Q => 
                           n_1253, QN => n55);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n9341, CK => CLK, Q => 
                           n_1254, QN => n57);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n9340, CK => CLK, Q => 
                           n_1255, QN => n59);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n9339, CK => CLK, Q => 
                           n_1256, QN => n61);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n9338, CK => CLK, Q => 
                           n_1257, QN => n63);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n9337, CK => CLK, Q => n553
                           , QN => n5824);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n9336, CK => CLK, Q => n555
                           , QN => n5820);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n9335, CK => CLK, Q => n557
                           , QN => n5816);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n9334, CK => CLK, Q => n559
                           , QN => n5812);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n9333, CK => CLK, Q => n561
                           , QN => n5808);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n9332, CK => CLK, Q => n563
                           , QN => n5804);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n9331, CK => CLK, Q => n565
                           , QN => n5800);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n9330, CK => CLK, Q => n567
                           , QN => n5796);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n9329, CK => CLK, Q => n569
                           , QN => n5792);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n9328, CK => CLK, Q => n571
                           , QN => n5788);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n9327, CK => CLK, Q => n573
                           , QN => n5784);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n9326, CK => CLK, Q => n575
                           , QN => n5780);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n9325, CK => CLK, Q => n577
                           , QN => n5776);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n9324, CK => CLK, Q => n579
                           , QN => n5772);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n9323, CK => CLK, Q => n581
                           , QN => n5768);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n9322, CK => CLK, Q => n583
                           , QN => n5764);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n9321, CK => CLK, Q => n585
                           , QN => n5760);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n9320, CK => CLK, Q => n587
                           , QN => n5756);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n9319, CK => CLK, Q => n589
                           , QN => n5752);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n9318, CK => CLK, Q => n591
                           , QN => n5748);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n9317, CK => CLK, Q => n593
                           , QN => n5744);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n9316, CK => CLK, Q => n595
                           , QN => n5740);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n9315, CK => CLK, Q => n597,
                           QN => n5736);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n9314, CK => CLK, Q => n599,
                           QN => n5732);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n9313, CK => CLK, Q => n601,
                           QN => n5728);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n9312, CK => CLK, Q => n603,
                           QN => n5724);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n9311, CK => CLK, Q => n605,
                           QN => n5720);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n9310, CK => CLK, Q => n607,
                           QN => n5716);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n9309, CK => CLK, Q => n609,
                           QN => n5712);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n9308, CK => CLK, Q => n611,
                           QN => n5708);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n9307, CK => CLK, Q => n613,
                           QN => n5704);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n9306, CK => CLK, Q => n615,
                           QN => n5700);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n9305, CK => CLK, Q => n97,
                           QN => n5825);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n9304, CK => CLK, Q => n99,
                           QN => n5821);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n9303, CK => CLK, Q => n101
                           , QN => n5817);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n9302, CK => CLK, Q => n103
                           , QN => n5813);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n9301, CK => CLK, Q => n105
                           , QN => n5809);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n9300, CK => CLK, Q => n107
                           , QN => n5805);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n9299, CK => CLK, Q => n109
                           , QN => n5801);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n9298, CK => CLK, Q => n111
                           , QN => n5797);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n9297, CK => CLK, Q => n113
                           , QN => n5793);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n9296, CK => CLK, Q => n115
                           , QN => n5789);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n9295, CK => CLK, Q => n117
                           , QN => n5785);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n9294, CK => CLK, Q => n119
                           , QN => n5781);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n9293, CK => CLK, Q => n121
                           , QN => n5777);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n9292, CK => CLK, Q => n123
                           , QN => n5773);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n9291, CK => CLK, Q => n125
                           , QN => n5769);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n9290, CK => CLK, Q => n127
                           , QN => n5765);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n9289, CK => CLK, Q => n129
                           , QN => n5761);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n9288, CK => CLK, Q => n131
                           , QN => n5757);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n9287, CK => CLK, Q => n133
                           , QN => n5753);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n9286, CK => CLK, Q => n135
                           , QN => n5749);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n9285, CK => CLK, Q => n137
                           , QN => n5745);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n9284, CK => CLK, Q => n139
                           , QN => n5741);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n9283, CK => CLK, Q => n141,
                           QN => n5737);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n9282, CK => CLK, Q => n143,
                           QN => n5733);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n9281, CK => CLK, Q => n145,
                           QN => n5729);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n9280, CK => CLK, Q => n147,
                           QN => n5725);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n9279, CK => CLK, Q => n149,
                           QN => n5721);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n9278, CK => CLK, Q => n151,
                           QN => n5717);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n9277, CK => CLK, Q => n153,
                           QN => n5713);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n9276, CK => CLK, Q => n155,
                           QN => n5709);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n9275, CK => CLK, Q => n157,
                           QN => n5705);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n9274, CK => CLK, Q => n159,
                           QN => n5701);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n9273, CK => CLK, Q => 
                           n6401, QN => n873);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n9272, CK => CLK, Q => 
                           n6400, QN => n874);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n9271, CK => CLK, Q => 
                           n6399, QN => n875);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n9270, CK => CLK, Q => 
                           n6398, QN => n876);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n9269, CK => CLK, Q => 
                           n6397, QN => n877);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n9268, CK => CLK, Q => 
                           n6396, QN => n878);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n9267, CK => CLK, Q => 
                           n6395, QN => n879);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n9266, CK => CLK, Q => 
                           n6394, QN => n880);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n9265, CK => CLK, Q => 
                           n6393, QN => n881);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n9264, CK => CLK, Q => 
                           n6392, QN => n882);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n9263, CK => CLK, Q => 
                           n6391, QN => n883);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n9262, CK => CLK, Q => 
                           n6390, QN => n884);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n9261, CK => CLK, Q => 
                           n6389, QN => n885);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n9260, CK => CLK, Q => 
                           n6388, QN => n886);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n9259, CK => CLK, Q => 
                           n6387, QN => n887);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n9258, CK => CLK, Q => 
                           n6386, QN => n888);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n9257, CK => CLK, Q => 
                           n6385, QN => n889);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n9256, CK => CLK, Q => 
                           n6384, QN => n890);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n9255, CK => CLK, Q => 
                           n6383, QN => n891);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n9254, CK => CLK, Q => 
                           n6382, QN => n892);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n9253, CK => CLK, Q => 
                           n6381, QN => n893);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n9252, CK => CLK, Q => 
                           n6380, QN => n894);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n9251, CK => CLK, Q => n6379
                           , QN => n895);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n9250, CK => CLK, Q => n6378
                           , QN => n896);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n9249, CK => CLK, Q => n6377
                           , QN => n897);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n9248, CK => CLK, Q => n6376
                           , QN => n898);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n9247, CK => CLK, Q => n6375
                           , QN => n899);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n9246, CK => CLK, Q => n6374
                           , QN => n900);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n9245, CK => CLK, Q => n6373
                           , QN => n901);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n9244, CK => CLK, Q => n6372
                           , QN => n902);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n9243, CK => CLK, Q => n6371
                           , QN => n903);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n9242, CK => CLK, Q => n6370
                           , QN => n904);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n9241, CK => CLK, Q => 
                           n6369, QN => n1225);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n9240, CK => CLK, Q => 
                           n6368, QN => n1226);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n9239, CK => CLK, Q => 
                           n6367, QN => n1227);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n9238, CK => CLK, Q => 
                           n6366, QN => n1228);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n9237, CK => CLK, Q => 
                           n6365, QN => n1229);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n9236, CK => CLK, Q => 
                           n6364, QN => n1230);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n9235, CK => CLK, Q => 
                           n6363, QN => n1231);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n9234, CK => CLK, Q => 
                           n6362, QN => n1232);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n9233, CK => CLK, Q => 
                           n6361, QN => n1233);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n9232, CK => CLK, Q => 
                           n6360, QN => n1234);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n9231, CK => CLK, Q => 
                           n6359, QN => n1235);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n9230, CK => CLK, Q => 
                           n6358, QN => n1236);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n9229, CK => CLK, Q => 
                           n6357, QN => n1237);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n9228, CK => CLK, Q => 
                           n6356, QN => n1238);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n9227, CK => CLK, Q => 
                           n6355, QN => n1239);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n9226, CK => CLK, Q => 
                           n6354, QN => n1240);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n9225, CK => CLK, Q => 
                           n6353, QN => n1241);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n9224, CK => CLK, Q => 
                           n6352, QN => n1242);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n9223, CK => CLK, Q => 
                           n6351, QN => n1243);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n9222, CK => CLK, Q => 
                           n6350, QN => n1244);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n9221, CK => CLK, Q => 
                           n6349, QN => n1245);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n9220, CK => CLK, Q => 
                           n6348, QN => n1246);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n9219, CK => CLK, Q => n6347
                           , QN => n1247);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n9218, CK => CLK, Q => n6346
                           , QN => n1248);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n9217, CK => CLK, Q => n6345
                           , QN => n1249);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n9216, CK => CLK, Q => n6344
                           , QN => n1250);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n9215, CK => CLK, Q => n6343
                           , QN => n1251);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n9214, CK => CLK, Q => n6342
                           , QN => n1252);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n9213, CK => CLK, Q => n6341
                           , QN => n1253);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n9212, CK => CLK, Q => n6340
                           , QN => n1254);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n9211, CK => CLK, Q => n6339
                           , QN => n1255);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n9210, CK => CLK, Q => n6338
                           , QN => n1256);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n9209, CK => CLK, Q => 
                           n_1258, QN => n5185);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n9208, CK => CLK, Q => 
                           n_1259, QN => n5184);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n9207, CK => CLK, Q => 
                           n_1260, QN => n5183);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n9206, CK => CLK, Q => 
                           n_1261, QN => n5182);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n9205, CK => CLK, Q => 
                           n_1262, QN => n5181);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n9204, CK => CLK, Q => 
                           n_1263, QN => n5180);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n9203, CK => CLK, Q => 
                           n_1264, QN => n5179);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n9202, CK => CLK, Q => 
                           n_1265, QN => n5178);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n9201, CK => CLK, Q => 
                           n_1266, QN => n5177);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n9200, CK => CLK, Q => 
                           n_1267, QN => n5176);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n9199, CK => CLK, Q => 
                           n_1268, QN => n5175);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n9198, CK => CLK, Q => 
                           n_1269, QN => n5174);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n9197, CK => CLK, Q => 
                           n_1270, QN => n5173);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n9196, CK => CLK, Q => 
                           n_1271, QN => n5172);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n9195, CK => CLK, Q => 
                           n_1272, QN => n5171);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n9194, CK => CLK, Q => 
                           n_1273, QN => n5170);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n9193, CK => CLK, Q => 
                           n_1274, QN => n5169);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n9192, CK => CLK, Q => 
                           n_1275, QN => n5168);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n9191, CK => CLK, Q => 
                           n_1276, QN => n5167);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n9190, CK => CLK, Q => 
                           n_1277, QN => n5166);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n9189, CK => CLK, Q => 
                           n_1278, QN => n5165);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n9188, CK => CLK, Q => 
                           n_1279, QN => n5164);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n9187, CK => CLK, Q => 
                           n_1280, QN => n5163);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n9186, CK => CLK, Q => 
                           n_1281, QN => n5162);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n9185, CK => CLK, Q => 
                           n_1282, QN => n5161);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n9184, CK => CLK, Q => 
                           n_1283, QN => n5160);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n9183, CK => CLK, Q => 
                           n_1284, QN => n5159);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n9182, CK => CLK, Q => 
                           n_1285, QN => n5158);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n9181, CK => CLK, Q => 
                           n_1286, QN => n5157);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n9180, CK => CLK, Q => 
                           n_1287, QN => n5156);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n9179, CK => CLK, Q => 
                           n_1288, QN => n5155);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n9178, CK => CLK, Q => 
                           n_1289, QN => n5154);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n9177, CK => CLK, Q => 
                           n_1290, QN => n5153);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n9176, CK => CLK, Q => 
                           n_1291, QN => n5152);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n9175, CK => CLK, Q => 
                           n_1292, QN => n5151);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n9174, CK => CLK, Q => 
                           n_1293, QN => n5150);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n9173, CK => CLK, Q => 
                           n_1294, QN => n5149);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n9172, CK => CLK, Q => 
                           n_1295, QN => n5148);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n9171, CK => CLK, Q => 
                           n_1296, QN => n5147);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n9170, CK => CLK, Q => 
                           n_1297, QN => n5146);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n9169, CK => CLK, Q => 
                           n_1298, QN => n5145);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n9168, CK => CLK, Q => 
                           n_1299, QN => n5144);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n9167, CK => CLK, Q => 
                           n_1300, QN => n5143);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n9166, CK => CLK, Q => 
                           n_1301, QN => n5142);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n9165, CK => CLK, Q => 
                           n_1302, QN => n5141);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n9164, CK => CLK, Q => 
                           n_1303, QN => n5140);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n9163, CK => CLK, Q => 
                           n_1304, QN => n5139);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n9162, CK => CLK, Q => 
                           n_1305, QN => n5138);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n9161, CK => CLK, Q => 
                           n_1306, QN => n5137);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n9160, CK => CLK, Q => 
                           n_1307, QN => n5136);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n9159, CK => CLK, Q => 
                           n_1308, QN => n5135);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n9158, CK => CLK, Q => 
                           n_1309, QN => n5134);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n9157, CK => CLK, Q => 
                           n_1310, QN => n5133);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n9156, CK => CLK, Q => 
                           n_1311, QN => n5132);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n9155, CK => CLK, Q => 
                           n_1312, QN => n5131);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n9154, CK => CLK, Q => 
                           n_1313, QN => n5130);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n9153, CK => CLK, Q => 
                           n_1314, QN => n5129);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n9152, CK => CLK, Q => 
                           n_1315, QN => n5128);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n9151, CK => CLK, Q => 
                           n_1316, QN => n5127);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n9150, CK => CLK, Q => 
                           n_1317, QN => n5126);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n9149, CK => CLK, Q => 
                           n_1318, QN => n5125);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n9148, CK => CLK, Q => 
                           n_1319, QN => n5124);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n9147, CK => CLK, Q => 
                           n_1320, QN => n5123);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n9146, CK => CLK, Q => 
                           n_1321, QN => n5122);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n9145, CK => CLK, Q => 
                           n_1322, QN => n5121);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n9144, CK => CLK, Q => 
                           n_1323, QN => n5120);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n9143, CK => CLK, Q => 
                           n_1324, QN => n5119);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n9142, CK => CLK, Q => 
                           n_1325, QN => n5118);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n9141, CK => CLK, Q => 
                           n_1326, QN => n5117);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n9140, CK => CLK, Q => 
                           n_1327, QN => n5116);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n9139, CK => CLK, Q => 
                           n_1328, QN => n5115);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n9138, CK => CLK, Q => 
                           n_1329, QN => n5114);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n9137, CK => CLK, Q => 
                           n_1330, QN => n5113);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n9136, CK => CLK, Q => 
                           n_1331, QN => n5112);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n9135, CK => CLK, Q => 
                           n_1332, QN => n5111);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n9134, CK => CLK, Q => 
                           n_1333, QN => n5110);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n9133, CK => CLK, Q => 
                           n_1334, QN => n5109);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n9132, CK => CLK, Q => 
                           n_1335, QN => n5108);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n9131, CK => CLK, Q => 
                           n_1336, QN => n5107);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n9130, CK => CLK, Q => 
                           n_1337, QN => n5106);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n9129, CK => CLK, Q => 
                           n_1338, QN => n5105);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n9128, CK => CLK, Q => 
                           n_1339, QN => n5104);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n9127, CK => CLK, Q => 
                           n_1340, QN => n5103);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n9126, CK => CLK, Q => 
                           n_1341, QN => n5102);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n9125, CK => CLK, Q => 
                           n_1342, QN => n5101);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n9124, CK => CLK, Q => 
                           n_1343, QN => n5100);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n9123, CK => CLK, Q => 
                           n_1344, QN => n5099);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n9122, CK => CLK, Q => 
                           n_1345, QN => n5098);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n9121, CK => CLK, Q => 
                           n_1346, QN => n5097);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n9120, CK => CLK, Q => 
                           n_1347, QN => n5096);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n9119, CK => CLK, Q => 
                           n_1348, QN => n5095);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n9118, CK => CLK, Q => 
                           n_1349, QN => n5094);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n9117, CK => CLK, Q => 
                           n_1350, QN => n5093);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n9116, CK => CLK, Q => 
                           n_1351, QN => n5092);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n9115, CK => CLK, Q => 
                           n_1352, QN => n5091);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n9114, CK => CLK, Q => 
                           n_1353, QN => n5090);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n9113, CK => CLK, Q => 
                           n_1354, QN => n65);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n9112, CK => CLK, Q => 
                           n_1355, QN => n66);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n9111, CK => CLK, Q => 
                           n_1356, QN => n67);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n9110, CK => CLK, Q => 
                           n_1357, QN => n68);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n9109, CK => CLK, Q => 
                           n_1358, QN => n69);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n9108, CK => CLK, Q => 
                           n_1359, QN => n70);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n9107, CK => CLK, Q => 
                           n_1360, QN => n71);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n9106, CK => CLK, Q => 
                           n_1361, QN => n72);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n9105, CK => CLK, Q => 
                           n_1362, QN => n73);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n9104, CK => CLK, Q => 
                           n_1363, QN => n74);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n9103, CK => CLK, Q => 
                           n_1364, QN => n75);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n9102, CK => CLK, Q => 
                           n_1365, QN => n76);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n9101, CK => CLK, Q => 
                           n_1366, QN => n77);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n9100, CK => CLK, Q => 
                           n_1367, QN => n78);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n9099, CK => CLK, Q => 
                           n_1368, QN => n79);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n9098, CK => CLK, Q => 
                           n_1369, QN => n80);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n9097, CK => CLK, Q => 
                           n_1370, QN => n81);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n9096, CK => CLK, Q => 
                           n_1371, QN => n82);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n9095, CK => CLK, Q => 
                           n_1372, QN => n83);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n9094, CK => CLK, Q => 
                           n_1373, QN => n84);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n9093, CK => CLK, Q => 
                           n_1374, QN => n85);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n9092, CK => CLK, Q => 
                           n_1375, QN => n86);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n9091, CK => CLK, Q => 
                           n_1376, QN => n87);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n9090, CK => CLK, Q => 
                           n_1377, QN => n88);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n9089, CK => CLK, Q => 
                           n_1378, QN => n89);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n9088, CK => CLK, Q => 
                           n_1379, QN => n90);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n9087, CK => CLK, Q => 
                           n_1380, QN => n91);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n9086, CK => CLK, Q => 
                           n_1381, QN => n92);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n9085, CK => CLK, Q => 
                           n_1382, QN => n93);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n9084, CK => CLK, Q => 
                           n_1383, QN => n94);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n9083, CK => CLK, Q => 
                           n_1384, QN => n95);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n9082, CK => CLK, Q => 
                           n_1385, QN => n96);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n9081, CK => CLK, Q => 
                           n_1386, QN => n425);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n9080, CK => CLK, Q => 
                           n_1387, QN => n426);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n9079, CK => CLK, Q => 
                           n_1388, QN => n427);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n9078, CK => CLK, Q => 
                           n_1389, QN => n428);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n9077, CK => CLK, Q => 
                           n_1390, QN => n429);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n9076, CK => CLK, Q => 
                           n_1391, QN => n430);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n9075, CK => CLK, Q => 
                           n_1392, QN => n431);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n9074, CK => CLK, Q => 
                           n_1393, QN => n432);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n9073, CK => CLK, Q => 
                           n_1394, QN => n433);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n9072, CK => CLK, Q => 
                           n_1395, QN => n434);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n9071, CK => CLK, Q => 
                           n_1396, QN => n435);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n9070, CK => CLK, Q => 
                           n_1397, QN => n436);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n9069, CK => CLK, Q => 
                           n_1398, QN => n437);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n9068, CK => CLK, Q => 
                           n_1399, QN => n438);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n9067, CK => CLK, Q => 
                           n_1400, QN => n439);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n9066, CK => CLK, Q => 
                           n_1401, QN => n440);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n9065, CK => CLK, Q => 
                           n_1402, QN => n441);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n9064, CK => CLK, Q => 
                           n_1403, QN => n442);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n9063, CK => CLK, Q => 
                           n_1404, QN => n443);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n9062, CK => CLK, Q => 
                           n_1405, QN => n444);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n9061, CK => CLK, Q => 
                           n_1406, QN => n445);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n9060, CK => CLK, Q => 
                           n_1407, QN => n446);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n9059, CK => CLK, Q => 
                           n_1408, QN => n447);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n9058, CK => CLK, Q => 
                           n_1409, QN => n448);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n9057, CK => CLK, Q => 
                           n_1410, QN => n449);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n9056, CK => CLK, Q => 
                           n_1411, QN => n450);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n9055, CK => CLK, Q => 
                           n_1412, QN => n451);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n9054, CK => CLK, Q => 
                           n_1413, QN => n452);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n9053, CK => CLK, Q => 
                           n_1414, QN => n453);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n9052, CK => CLK, Q => 
                           n_1415, QN => n454);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n9051, CK => CLK, Q => 
                           n_1416, QN => n455);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n9050, CK => CLK, Q => 
                           n_1417, QN => n456);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n9049, CK => CLK, Q => n521
                           , QN => n5692);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n9048, CK => CLK, Q => n522
                           , QN => n5682);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n9047, CK => CLK, Q => n523
                           , QN => n5672);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n9046, CK => CLK, Q => n524
                           , QN => n5662);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n9045, CK => CLK, Q => n525
                           , QN => n5652);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n9044, CK => CLK, Q => n526
                           , QN => n5642);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n9043, CK => CLK, Q => n527
                           , QN => n5632);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n9042, CK => CLK, Q => n528
                           , QN => n5622);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n9041, CK => CLK, Q => n529
                           , QN => n5612);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n9040, CK => CLK, Q => n530
                           , QN => n5602);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n9039, CK => CLK, Q => n531
                           , QN => n5592);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n9038, CK => CLK, Q => n532
                           , QN => n5582);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n9037, CK => CLK, Q => n533
                           , QN => n5572);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n9036, CK => CLK, Q => n534
                           , QN => n5562);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n9035, CK => CLK, Q => n535
                           , QN => n5552);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n9034, CK => CLK, Q => n536
                           , QN => n5542);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n9033, CK => CLK, Q => n537
                           , QN => n5532);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n9032, CK => CLK, Q => n538
                           , QN => n5522);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n9031, CK => CLK, Q => n539
                           , QN => n5512);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n9030, CK => CLK, Q => n540
                           , QN => n5502);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n9029, CK => CLK, Q => n541
                           , QN => n5492);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n9028, CK => CLK, Q => n542
                           , QN => n5482);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n9027, CK => CLK, Q => n543,
                           QN => n5472);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n9026, CK => CLK, Q => n544,
                           QN => n5462);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n9025, CK => CLK, Q => n545,
                           QN => n5452);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n9024, CK => CLK, Q => n546,
                           QN => n5442);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n9023, CK => CLK, Q => n547,
                           QN => n5432);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n9022, CK => CLK, Q => n548,
                           QN => n5422);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n9021, CK => CLK, Q => n549,
                           QN => n5412);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n9020, CK => CLK, Q => n550,
                           QN => n5402);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n9019, CK => CLK, Q => n551,
                           QN => n5392);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n9018, CK => CLK, Q => n552,
                           QN => n5382);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n9017, CK => CLK, Q => n161
                           , QN => n5693);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n9016, CK => CLK, Q => n162
                           , QN => n5683);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n9015, CK => CLK, Q => n163
                           , QN => n5673);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n9014, CK => CLK, Q => n164
                           , QN => n5663);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n9013, CK => CLK, Q => n165
                           , QN => n5653);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n9012, CK => CLK, Q => n166
                           , QN => n5643);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n9011, CK => CLK, Q => n167
                           , QN => n5633);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n9010, CK => CLK, Q => n168
                           , QN => n5623);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n9009, CK => CLK, Q => n169
                           , QN => n5613);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n9008, CK => CLK, Q => n170
                           , QN => n5603);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n9007, CK => CLK, Q => n171
                           , QN => n5593);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n9006, CK => CLK, Q => n172
                           , QN => n5583);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n9005, CK => CLK, Q => n173
                           , QN => n5573);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n9004, CK => CLK, Q => n174
                           , QN => n5563);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n9003, CK => CLK, Q => n175
                           , QN => n5553);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n9002, CK => CLK, Q => n176
                           , QN => n5543);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n9001, CK => CLK, Q => n177
                           , QN => n5533);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n9000, CK => CLK, Q => n178
                           , QN => n5523);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n8999, CK => CLK, Q => n179
                           , QN => n5513);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n8998, CK => CLK, Q => n180
                           , QN => n5503);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n8997, CK => CLK, Q => n181
                           , QN => n5493);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n8996, CK => CLK, Q => n182
                           , QN => n5483);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n8995, CK => CLK, Q => n183,
                           QN => n5473);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n8994, CK => CLK, Q => n184,
                           QN => n5463);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n8993, CK => CLK, Q => n185,
                           QN => n5453);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n8992, CK => CLK, Q => n186,
                           QN => n5443);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n8991, CK => CLK, Q => n187,
                           QN => n5433);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n8990, CK => CLK, Q => n188,
                           QN => n5423);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n8989, CK => CLK, Q => n189,
                           QN => n5413);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n8988, CK => CLK, Q => n190,
                           QN => n5403);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n8987, CK => CLK, Q => n191,
                           QN => n5393);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n8986, CK => CLK, Q => n192,
                           QN => n5383);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n8985, CK => CLK, Q => 
                           n6337, QN => n905);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n8984, CK => CLK, Q => 
                           n6336, QN => n906);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n8983, CK => CLK, Q => 
                           n6335, QN => n907);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n8982, CK => CLK, Q => 
                           n6334, QN => n908);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n8981, CK => CLK, Q => 
                           n6333, QN => n909);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n8980, CK => CLK, Q => 
                           n6332, QN => n910);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n8979, CK => CLK, Q => 
                           n6331, QN => n911);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n8978, CK => CLK, Q => 
                           n6330, QN => n912);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n8977, CK => CLK, Q => 
                           n6329, QN => n913);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n8976, CK => CLK, Q => 
                           n6328, QN => n914);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n8975, CK => CLK, Q => 
                           n6327, QN => n915);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n8974, CK => CLK, Q => 
                           n6326, QN => n916);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n8973, CK => CLK, Q => 
                           n6325, QN => n917);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n8972, CK => CLK, Q => 
                           n6324, QN => n918);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n8971, CK => CLK, Q => 
                           n6323, QN => n919);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n8970, CK => CLK, Q => 
                           n6322, QN => n920);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n8969, CK => CLK, Q => 
                           n6321, QN => n921);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n8968, CK => CLK, Q => 
                           n6320, QN => n922);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n8967, CK => CLK, Q => 
                           n6319, QN => n923);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n8966, CK => CLK, Q => 
                           n6318, QN => n924);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n8965, CK => CLK, Q => 
                           n6317, QN => n925);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n8964, CK => CLK, Q => 
                           n6316, QN => n926);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n8963, CK => CLK, Q => n6315
                           , QN => n927);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n8962, CK => CLK, Q => n6314
                           , QN => n928);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n8961, CK => CLK, Q => n6313
                           , QN => n929);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n8960, CK => CLK, Q => n6312
                           , QN => n930);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n8959, CK => CLK, Q => n6311
                           , QN => n931);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n8958, CK => CLK, Q => n6310
                           , QN => n932);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n8957, CK => CLK, Q => n6309
                           , QN => n933);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n8956, CK => CLK, Q => n6308
                           , QN => n934);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n8955, CK => CLK, Q => n6307
                           , QN => n935);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n8954, CK => CLK, Q => n6306
                           , QN => n936);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n8953, CK => CLK, Q => 
                           n6305, QN => n1257);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n8952, CK => CLK, Q => 
                           n6304, QN => n1258);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n8951, CK => CLK, Q => 
                           n6303, QN => n1259);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n8950, CK => CLK, Q => 
                           n6302, QN => n1260);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n8949, CK => CLK, Q => 
                           n6301, QN => n1261);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n8948, CK => CLK, Q => 
                           n6300, QN => n1262);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n8947, CK => CLK, Q => 
                           n6299, QN => n1263);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n8946, CK => CLK, Q => 
                           n6298, QN => n1264);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n8945, CK => CLK, Q => 
                           n6297, QN => n1265);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n8944, CK => CLK, Q => 
                           n6296, QN => n1266);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n8943, CK => CLK, Q => 
                           n6295, QN => n1267);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n8942, CK => CLK, Q => 
                           n6294, QN => n1268);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n8941, CK => CLK, Q => 
                           n6293, QN => n1269);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n8940, CK => CLK, Q => 
                           n6292, QN => n1270);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n8939, CK => CLK, Q => 
                           n6291, QN => n1271);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n8938, CK => CLK, Q => 
                           n6290, QN => n1272);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n8937, CK => CLK, Q => 
                           n6289, QN => n1273);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n8936, CK => CLK, Q => 
                           n6288, QN => n1274);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n8935, CK => CLK, Q => 
                           n6287, QN => n1275);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n8934, CK => CLK, Q => 
                           n6286, QN => n1276);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n8933, CK => CLK, Q => 
                           n6285, QN => n1277);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n8932, CK => CLK, Q => 
                           n6284, QN => n1278);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n8931, CK => CLK, Q => n6283
                           , QN => n1279);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n8930, CK => CLK, Q => n6282
                           , QN => n1280);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n8929, CK => CLK, Q => n6281
                           , QN => n1281);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n8928, CK => CLK, Q => n6280
                           , QN => n1282);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n8927, CK => CLK, Q => n6279
                           , QN => n1283);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n8926, CK => CLK, Q => n6278
                           , QN => n1284);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n8925, CK => CLK, Q => n6277
                           , QN => n1285);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n8924, CK => CLK, Q => n6276
                           , QN => n1286);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n8923, CK => CLK, Q => n6275
                           , QN => n1287);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n8922, CK => CLK, Q => n6274
                           , QN => n1288);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n8921, CK => CLK, Q => 
                           n_1418, QN => n5089);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n8920, CK => CLK, Q => 
                           n_1419, QN => n5088);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n8919, CK => CLK, Q => 
                           n_1420, QN => n5087);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n8918, CK => CLK, Q => 
                           n_1421, QN => n5086);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n8917, CK => CLK, Q => 
                           n_1422, QN => n5085);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n8916, CK => CLK, Q => 
                           n_1423, QN => n5084);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n8915, CK => CLK, Q => 
                           n_1424, QN => n5083);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n8914, CK => CLK, Q => 
                           n_1425, QN => n5082);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n8913, CK => CLK, Q => 
                           n_1426, QN => n5081);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n8912, CK => CLK, Q => 
                           n_1427, QN => n5080);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n8911, CK => CLK, Q => 
                           n_1428, QN => n5079);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n8910, CK => CLK, Q => 
                           n_1429, QN => n5078);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n8909, CK => CLK, Q => 
                           n_1430, QN => n5077);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n8908, CK => CLK, Q => 
                           n_1431, QN => n5076);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n8907, CK => CLK, Q => 
                           n_1432, QN => n5075);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n8906, CK => CLK, Q => 
                           n_1433, QN => n5074);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n8905, CK => CLK, Q => 
                           n_1434, QN => n5073);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n8904, CK => CLK, Q => 
                           n_1435, QN => n5072);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n8903, CK => CLK, Q => 
                           n_1436, QN => n5071);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n8902, CK => CLK, Q => 
                           n_1437, QN => n5070);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n8901, CK => CLK, Q => 
                           n_1438, QN => n5069);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n8900, CK => CLK, Q => 
                           n_1439, QN => n5068);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n8899, CK => CLK, Q => 
                           n_1440, QN => n5067);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n8898, CK => CLK, Q => 
                           n_1441, QN => n5066);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n8897, CK => CLK, Q => 
                           n_1442, QN => n5065);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n8896, CK => CLK, Q => 
                           n_1443, QN => n5064);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n8895, CK => CLK, Q => 
                           n_1444, QN => n5063);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n8894, CK => CLK, Q => 
                           n_1445, QN => n5062);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n8893, CK => CLK, Q => 
                           n_1446, QN => n5061);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n8892, CK => CLK, Q => 
                           n_1447, QN => n5060);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n8891, CK => CLK, Q => 
                           n_1448, QN => n5059);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n8890, CK => CLK, Q => 
                           n_1449, QN => n5058);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n8889, CK => CLK, Q => 
                           n_1450, QN => n5057);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n8888, CK => CLK, Q => 
                           n_1451, QN => n5056);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n8887, CK => CLK, Q => 
                           n_1452, QN => n5055);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n8886, CK => CLK, Q => 
                           n_1453, QN => n5054);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n8885, CK => CLK, Q => 
                           n_1454, QN => n5053);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n8884, CK => CLK, Q => 
                           n_1455, QN => n5052);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n8883, CK => CLK, Q => 
                           n_1456, QN => n5051);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n8882, CK => CLK, Q => 
                           n_1457, QN => n5050);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n8881, CK => CLK, Q => 
                           n_1458, QN => n5049);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n8880, CK => CLK, Q => 
                           n_1459, QN => n5048);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n8879, CK => CLK, Q => 
                           n_1460, QN => n5047);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n8878, CK => CLK, Q => 
                           n_1461, QN => n5046);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n8877, CK => CLK, Q => 
                           n_1462, QN => n5045);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n8876, CK => CLK, Q => 
                           n_1463, QN => n5044);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n8875, CK => CLK, Q => 
                           n_1464, QN => n5043);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n8874, CK => CLK, Q => 
                           n_1465, QN => n5042);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n8873, CK => CLK, Q => 
                           n_1466, QN => n5041);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n8872, CK => CLK, Q => 
                           n_1467, QN => n5040);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n8871, CK => CLK, Q => 
                           n_1468, QN => n5039);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n8870, CK => CLK, Q => 
                           n_1469, QN => n5038);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n8869, CK => CLK, Q => 
                           n_1470, QN => n5037);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n8868, CK => CLK, Q => 
                           n_1471, QN => n5036);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n8867, CK => CLK, Q => 
                           n_1472, QN => n5035);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n8866, CK => CLK, Q => 
                           n_1473, QN => n5034);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n8865, CK => CLK, Q => 
                           n_1474, QN => n5033);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n8864, CK => CLK, Q => 
                           n_1475, QN => n5032);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n8863, CK => CLK, Q => 
                           n_1476, QN => n5031);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n8862, CK => CLK, Q => 
                           n_1477, QN => n5030);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n8861, CK => CLK, Q => 
                           n_1478, QN => n5029);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n8860, CK => CLK, Q => 
                           n_1479, QN => n5028);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n8859, CK => CLK, Q => 
                           n_1480, QN => n5027);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n8858, CK => CLK, Q => 
                           n_1481, QN => n5026);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n8857, CK => CLK, Q => 
                           n_1482, QN => n5025);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n8856, CK => CLK, Q => 
                           n_1483, QN => n5024);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n8855, CK => CLK, Q => 
                           n_1484, QN => n5023);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n8854, CK => CLK, Q => 
                           n_1485, QN => n5022);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n8853, CK => CLK, Q => 
                           n_1486, QN => n5021);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n8852, CK => CLK, Q => 
                           n_1487, QN => n5020);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n8851, CK => CLK, Q => 
                           n_1488, QN => n5019);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n8850, CK => CLK, Q => 
                           n_1489, QN => n5018);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n8849, CK => CLK, Q => 
                           n_1490, QN => n5017);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n8848, CK => CLK, Q => 
                           n_1491, QN => n5016);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n8847, CK => CLK, Q => 
                           n_1492, QN => n5015);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n8846, CK => CLK, Q => 
                           n_1493, QN => n5014);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n8845, CK => CLK, Q => 
                           n_1494, QN => n5013);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n8844, CK => CLK, Q => 
                           n_1495, QN => n5012);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n8843, CK => CLK, Q => 
                           n_1496, QN => n5011);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n8842, CK => CLK, Q => 
                           n_1497, QN => n5010);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n8841, CK => CLK, Q => 
                           n_1498, QN => n5009);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n8840, CK => CLK, Q => 
                           n_1499, QN => n5008);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n8839, CK => CLK, Q => 
                           n_1500, QN => n5007);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n8838, CK => CLK, Q => 
                           n_1501, QN => n5006);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n8837, CK => CLK, Q => 
                           n_1502, QN => n5005);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n8836, CK => CLK, Q => 
                           n_1503, QN => n5004);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n8835, CK => CLK, Q => 
                           n_1504, QN => n5003);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n8834, CK => CLK, Q => 
                           n_1505, QN => n5002);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n8833, CK => CLK, Q => 
                           n_1506, QN => n5001);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n8832, CK => CLK, Q => 
                           n_1507, QN => n5000);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n8831, CK => CLK, Q => 
                           n_1508, QN => n4999);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n8830, CK => CLK, Q => 
                           n_1509, QN => n4998);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n8829, CK => CLK, Q => 
                           n_1510, QN => n4997);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n8828, CK => CLK, Q => 
                           n_1511, QN => n4996);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n8827, CK => CLK, Q => 
                           n_1512, QN => n4995);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n8826, CK => CLK, Q => 
                           n_1513, QN => n4994);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n8825, CK => CLK, Q => 
                           n_1514, QN => n458);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n8824, CK => CLK, Q => 
                           n_1515, QN => n460);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n8823, CK => CLK, Q => 
                           n_1516, QN => n462);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n8822, CK => CLK, Q => 
                           n_1517, QN => n464);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n8821, CK => CLK, Q => 
                           n_1518, QN => n466);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n8820, CK => CLK, Q => 
                           n_1519, QN => n468);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n8819, CK => CLK, Q => 
                           n_1520, QN => n470);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n8818, CK => CLK, Q => 
                           n_1521, QN => n472);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n8817, CK => CLK, Q => 
                           n_1522, QN => n474);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n8816, CK => CLK, Q => 
                           n_1523, QN => n476);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n8815, CK => CLK, Q => 
                           n_1524, QN => n478);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n8814, CK => CLK, Q => 
                           n_1525, QN => n480);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n8813, CK => CLK, Q => 
                           n_1526, QN => n482);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n8812, CK => CLK, Q => 
                           n_1527, QN => n484);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n8811, CK => CLK, Q => 
                           n_1528, QN => n486);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n8810, CK => CLK, Q => 
                           n_1529, QN => n488);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n8809, CK => CLK, Q => 
                           n_1530, QN => n490);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n8808, CK => CLK, Q => 
                           n_1531, QN => n492);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n8807, CK => CLK, Q => 
                           n_1532, QN => n494);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n8806, CK => CLK, Q => 
                           n_1533, QN => n496);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n8805, CK => CLK, Q => 
                           n_1534, QN => n498);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n8804, CK => CLK, Q => 
                           n_1535, QN => n500);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n8803, CK => CLK, Q => 
                           n_1536, QN => n502);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n8802, CK => CLK, Q => 
                           n_1537, QN => n504);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n8801, CK => CLK, Q => 
                           n_1538, QN => n506);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n8800, CK => CLK, Q => 
                           n_1539, QN => n508);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n8799, CK => CLK, Q => 
                           n_1540, QN => n510);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n8798, CK => CLK, Q => 
                           n_1541, QN => n512);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n8797, CK => CLK, Q => 
                           n_1542, QN => n514);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n8796, CK => CLK, Q => 
                           n_1543, QN => n516);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n8795, CK => CLK, Q => 
                           n_1544, QN => n518);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n8794, CK => CLK, Q => 
                           n_1545, QN => n520);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n8793, CK => CLK, Q => 
                           n_1546, QN => n2);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n8792, CK => CLK, Q => 
                           n_1547, QN => n4);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n8791, CK => CLK, Q => 
                           n_1548, QN => n6);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n8790, CK => CLK, Q => 
                           n_1549, QN => n8);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n8789, CK => CLK, Q => 
                           n_1550, QN => n10);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n8788, CK => CLK, Q => 
                           n_1551, QN => n12);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n8787, CK => CLK, Q => 
                           n_1552, QN => n14);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n8786, CK => CLK, Q => 
                           n_1553, QN => n16);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n8785, CK => CLK, Q => 
                           n_1554, QN => n18);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n8784, CK => CLK, Q => 
                           n_1555, QN => n20);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n8783, CK => CLK, Q => 
                           n_1556, QN => n22);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n8782, CK => CLK, Q => 
                           n_1557, QN => n24);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n8781, CK => CLK, Q => 
                           n_1558, QN => n26);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n8780, CK => CLK, Q => 
                           n_1559, QN => n28);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n8779, CK => CLK, Q => 
                           n_1560, QN => n30);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n8778, CK => CLK, Q => 
                           n_1561, QN => n32);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n8777, CK => CLK, Q => 
                           n_1562, QN => n34);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n8776, CK => CLK, Q => 
                           n_1563, QN => n36);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n8775, CK => CLK, Q => 
                           n_1564, QN => n38);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n8774, CK => CLK, Q => 
                           n_1565, QN => n40);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n8773, CK => CLK, Q => 
                           n_1566, QN => n42);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n8772, CK => CLK, Q => 
                           n_1567, QN => n44);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n8771, CK => CLK, Q => 
                           n_1568, QN => n46);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n8770, CK => CLK, Q => 
                           n_1569, QN => n48);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n8769, CK => CLK, Q => 
                           n_1570, QN => n50);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n8768, CK => CLK, Q => 
                           n_1571, QN => n52);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n8767, CK => CLK, Q => 
                           n_1572, QN => n54);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n8766, CK => CLK, Q => 
                           n_1573, QN => n56);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n8765, CK => CLK, Q => 
                           n_1574, QN => n58);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n8764, CK => CLK, Q => 
                           n_1575, QN => n60);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n8763, CK => CLK, Q => 
                           n_1576, QN => n62);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n8762, CK => CLK, Q => 
                           n_1577, QN => n64);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n8761, CK => CLK, Q => n554
                           , QN => n5822);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n8760, CK => CLK, Q => n556
                           , QN => n5818);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n8759, CK => CLK, Q => n558
                           , QN => n5814);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n8758, CK => CLK, Q => n560
                           , QN => n5810);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n8757, CK => CLK, Q => n562
                           , QN => n5806);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n8756, CK => CLK, Q => n564
                           , QN => n5802);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n8755, CK => CLK, Q => n566
                           , QN => n5798);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n8754, CK => CLK, Q => n568
                           , QN => n5794);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n8753, CK => CLK, Q => n570
                           , QN => n5790);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n8752, CK => CLK, Q => n572
                           , QN => n5786);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n8751, CK => CLK, Q => n574
                           , QN => n5782);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n8750, CK => CLK, Q => n576
                           , QN => n5778);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n8749, CK => CLK, Q => n578
                           , QN => n5774);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n8748, CK => CLK, Q => n580
                           , QN => n5770);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n8747, CK => CLK, Q => n582
                           , QN => n5766);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n8746, CK => CLK, Q => n584
                           , QN => n5762);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n8745, CK => CLK, Q => n586
                           , QN => n5758);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n8744, CK => CLK, Q => n588
                           , QN => n5754);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n8743, CK => CLK, Q => n590
                           , QN => n5750);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n8742, CK => CLK, Q => n592
                           , QN => n5746);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n8741, CK => CLK, Q => n594
                           , QN => n5742);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n8740, CK => CLK, Q => n596
                           , QN => n5738);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n8739, CK => CLK, Q => n598,
                           QN => n5734);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n8738, CK => CLK, Q => n600,
                           QN => n5730);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n8737, CK => CLK, Q => n602,
                           QN => n5726);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n8736, CK => CLK, Q => n604,
                           QN => n5722);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n8735, CK => CLK, Q => n606,
                           QN => n5718);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n8734, CK => CLK, Q => n608,
                           QN => n5714);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n8733, CK => CLK, Q => n610,
                           QN => n5710);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n8732, CK => CLK, Q => n612,
                           QN => n5706);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n8731, CK => CLK, Q => n614,
                           QN => n5702);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n8730, CK => CLK, Q => n616,
                           QN => n5698);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n8729, CK => CLK, Q => n98,
                           QN => n5823);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n8728, CK => CLK, Q => n100
                           , QN => n5819);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n8727, CK => CLK, Q => n102
                           , QN => n5815);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n8726, CK => CLK, Q => n104
                           , QN => n5811);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n8725, CK => CLK, Q => n106
                           , QN => n5807);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n8724, CK => CLK, Q => n108
                           , QN => n5803);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n8723, CK => CLK, Q => n110
                           , QN => n5799);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n8722, CK => CLK, Q => n112
                           , QN => n5795);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n8721, CK => CLK, Q => n114
                           , QN => n5791);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n8720, CK => CLK, Q => n116
                           , QN => n5787);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n8719, CK => CLK, Q => n118
                           , QN => n5783);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n8718, CK => CLK, Q => n120
                           , QN => n5779);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n8717, CK => CLK, Q => n122
                           , QN => n5775);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n8716, CK => CLK, Q => n124
                           , QN => n5771);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n8715, CK => CLK, Q => n126
                           , QN => n5767);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n8714, CK => CLK, Q => n128
                           , QN => n5763);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n8713, CK => CLK, Q => n130
                           , QN => n5759);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n8712, CK => CLK, Q => n132
                           , QN => n5755);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n8711, CK => CLK, Q => n134
                           , QN => n5751);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n8710, CK => CLK, Q => n136
                           , QN => n5747);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n8709, CK => CLK, Q => n138
                           , QN => n5743);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n8708, CK => CLK, Q => n140
                           , QN => n5739);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n8707, CK => CLK, Q => n142,
                           QN => n5735);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n8706, CK => CLK, Q => n144,
                           QN => n5731);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n8705, CK => CLK, Q => n146,
                           QN => n5727);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n8704, CK => CLK, Q => n148,
                           QN => n5723);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n8703, CK => CLK, Q => n150,
                           QN => n5719);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n8702, CK => CLK, Q => n152,
                           QN => n5715);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n8701, CK => CLK, Q => n154,
                           QN => n5711);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n8700, CK => CLK, Q => n156,
                           QN => n5707);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n8699, CK => CLK, Q => n158,
                           QN => n5703);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n8698, CK => CLK, Q => n160,
                           QN => n5699);
   REGISTERS_reg_40_31_inst : DFF_X1 port map( D => n8697, CK => CLK, Q => 
                           n6273, QN => n937);
   REGISTERS_reg_40_30_inst : DFF_X1 port map( D => n8696, CK => CLK, Q => 
                           n6272, QN => n938);
   REGISTERS_reg_40_29_inst : DFF_X1 port map( D => n8695, CK => CLK, Q => 
                           n6271, QN => n939);
   REGISTERS_reg_40_28_inst : DFF_X1 port map( D => n8694, CK => CLK, Q => 
                           n6270, QN => n940);
   REGISTERS_reg_40_27_inst : DFF_X1 port map( D => n8693, CK => CLK, Q => 
                           n6269, QN => n941);
   REGISTERS_reg_40_26_inst : DFF_X1 port map( D => n8692, CK => CLK, Q => 
                           n6268, QN => n942);
   REGISTERS_reg_40_25_inst : DFF_X1 port map( D => n8691, CK => CLK, Q => 
                           n6267, QN => n943);
   REGISTERS_reg_40_24_inst : DFF_X1 port map( D => n8690, CK => CLK, Q => 
                           n6266, QN => n944);
   REGISTERS_reg_40_23_inst : DFF_X1 port map( D => n8689, CK => CLK, Q => 
                           n6265, QN => n945);
   REGISTERS_reg_40_22_inst : DFF_X1 port map( D => n8688, CK => CLK, Q => 
                           n6264, QN => n946);
   REGISTERS_reg_40_21_inst : DFF_X1 port map( D => n8687, CK => CLK, Q => 
                           n6263, QN => n947);
   REGISTERS_reg_40_20_inst : DFF_X1 port map( D => n8686, CK => CLK, Q => 
                           n6262, QN => n948);
   REGISTERS_reg_40_19_inst : DFF_X1 port map( D => n8685, CK => CLK, Q => 
                           n6261, QN => n949);
   REGISTERS_reg_40_18_inst : DFF_X1 port map( D => n8684, CK => CLK, Q => 
                           n6260, QN => n950);
   REGISTERS_reg_40_17_inst : DFF_X1 port map( D => n8683, CK => CLK, Q => 
                           n6259, QN => n951);
   REGISTERS_reg_40_16_inst : DFF_X1 port map( D => n8682, CK => CLK, Q => 
                           n6258, QN => n952);
   REGISTERS_reg_40_15_inst : DFF_X1 port map( D => n8681, CK => CLK, Q => 
                           n6257, QN => n953);
   REGISTERS_reg_40_14_inst : DFF_X1 port map( D => n8680, CK => CLK, Q => 
                           n6256, QN => n954);
   REGISTERS_reg_40_13_inst : DFF_X1 port map( D => n8679, CK => CLK, Q => 
                           n6255, QN => n955);
   REGISTERS_reg_40_12_inst : DFF_X1 port map( D => n8678, CK => CLK, Q => 
                           n6254, QN => n956);
   REGISTERS_reg_40_11_inst : DFF_X1 port map( D => n8677, CK => CLK, Q => 
                           n6253, QN => n957);
   REGISTERS_reg_40_10_inst : DFF_X1 port map( D => n8676, CK => CLK, Q => 
                           n6252, QN => n958);
   REGISTERS_reg_40_9_inst : DFF_X1 port map( D => n8675, CK => CLK, Q => n6251
                           , QN => n959);
   REGISTERS_reg_40_8_inst : DFF_X1 port map( D => n8674, CK => CLK, Q => n6250
                           , QN => n960);
   REGISTERS_reg_40_7_inst : DFF_X1 port map( D => n8673, CK => CLK, Q => n6249
                           , QN => n961);
   REGISTERS_reg_40_6_inst : DFF_X1 port map( D => n8672, CK => CLK, Q => n6248
                           , QN => n962);
   REGISTERS_reg_40_5_inst : DFF_X1 port map( D => n8671, CK => CLK, Q => n6247
                           , QN => n963);
   REGISTERS_reg_40_4_inst : DFF_X1 port map( D => n8670, CK => CLK, Q => n6246
                           , QN => n964);
   REGISTERS_reg_40_3_inst : DFF_X1 port map( D => n8669, CK => CLK, Q => n6245
                           , QN => n965);
   REGISTERS_reg_40_2_inst : DFF_X1 port map( D => n8668, CK => CLK, Q => n6244
                           , QN => n966);
   REGISTERS_reg_40_1_inst : DFF_X1 port map( D => n8667, CK => CLK, Q => n6243
                           , QN => n967);
   REGISTERS_reg_40_0_inst : DFF_X1 port map( D => n8666, CK => CLK, Q => n6242
                           , QN => n968);
   REGISTERS_reg_41_31_inst : DFF_X1 port map( D => n8665, CK => CLK, Q => 
                           n6241, QN => n1289);
   REGISTERS_reg_41_30_inst : DFF_X1 port map( D => n8664, CK => CLK, Q => 
                           n6240, QN => n1290);
   REGISTERS_reg_41_29_inst : DFF_X1 port map( D => n8663, CK => CLK, Q => 
                           n6239, QN => n1291);
   REGISTERS_reg_41_28_inst : DFF_X1 port map( D => n8662, CK => CLK, Q => 
                           n6238, QN => n1292);
   REGISTERS_reg_41_27_inst : DFF_X1 port map( D => n8661, CK => CLK, Q => 
                           n6237, QN => n1293);
   REGISTERS_reg_41_26_inst : DFF_X1 port map( D => n8660, CK => CLK, Q => 
                           n6236, QN => n1294);
   REGISTERS_reg_41_25_inst : DFF_X1 port map( D => n8659, CK => CLK, Q => 
                           n6235, QN => n1295);
   REGISTERS_reg_41_24_inst : DFF_X1 port map( D => n8658, CK => CLK, Q => 
                           n6234, QN => n1296);
   REGISTERS_reg_41_23_inst : DFF_X1 port map( D => n8657, CK => CLK, Q => 
                           n6233, QN => n1297);
   REGISTERS_reg_41_22_inst : DFF_X1 port map( D => n8656, CK => CLK, Q => 
                           n6232, QN => n1298);
   REGISTERS_reg_41_21_inst : DFF_X1 port map( D => n8655, CK => CLK, Q => 
                           n6231, QN => n1299);
   REGISTERS_reg_41_20_inst : DFF_X1 port map( D => n8654, CK => CLK, Q => 
                           n6230, QN => n1300);
   REGISTERS_reg_41_19_inst : DFF_X1 port map( D => n8653, CK => CLK, Q => 
                           n6229, QN => n1301);
   REGISTERS_reg_41_18_inst : DFF_X1 port map( D => n8652, CK => CLK, Q => 
                           n6228, QN => n1302);
   REGISTERS_reg_41_17_inst : DFF_X1 port map( D => n8651, CK => CLK, Q => 
                           n6227, QN => n1303);
   REGISTERS_reg_41_16_inst : DFF_X1 port map( D => n8650, CK => CLK, Q => 
                           n6226, QN => n1304);
   REGISTERS_reg_41_15_inst : DFF_X1 port map( D => n8649, CK => CLK, Q => 
                           n6225, QN => n1305);
   REGISTERS_reg_41_14_inst : DFF_X1 port map( D => n8648, CK => CLK, Q => 
                           n6224, QN => n1306);
   REGISTERS_reg_41_13_inst : DFF_X1 port map( D => n8647, CK => CLK, Q => 
                           n6223, QN => n1307);
   REGISTERS_reg_41_12_inst : DFF_X1 port map( D => n8646, CK => CLK, Q => 
                           n6222, QN => n1308);
   REGISTERS_reg_41_11_inst : DFF_X1 port map( D => n8645, CK => CLK, Q => 
                           n6221, QN => n1309);
   REGISTERS_reg_41_10_inst : DFF_X1 port map( D => n8644, CK => CLK, Q => 
                           n6220, QN => n1310);
   REGISTERS_reg_41_9_inst : DFF_X1 port map( D => n8643, CK => CLK, Q => n6219
                           , QN => n1311);
   REGISTERS_reg_41_8_inst : DFF_X1 port map( D => n8642, CK => CLK, Q => n6218
                           , QN => n1312);
   REGISTERS_reg_41_7_inst : DFF_X1 port map( D => n8641, CK => CLK, Q => n6217
                           , QN => n1313);
   REGISTERS_reg_41_6_inst : DFF_X1 port map( D => n8640, CK => CLK, Q => n6216
                           , QN => n1314);
   REGISTERS_reg_41_5_inst : DFF_X1 port map( D => n8639, CK => CLK, Q => n6215
                           , QN => n1315);
   REGISTERS_reg_41_4_inst : DFF_X1 port map( D => n8638, CK => CLK, Q => n6214
                           , QN => n1316);
   REGISTERS_reg_41_3_inst : DFF_X1 port map( D => n8637, CK => CLK, Q => n6213
                           , QN => n1317);
   REGISTERS_reg_41_2_inst : DFF_X1 port map( D => n8636, CK => CLK, Q => n6212
                           , QN => n1318);
   REGISTERS_reg_41_1_inst : DFF_X1 port map( D => n8635, CK => CLK, Q => n6211
                           , QN => n1319);
   REGISTERS_reg_41_0_inst : DFF_X1 port map( D => n8634, CK => CLK, Q => n6210
                           , QN => n1320);
   REGISTERS_reg_42_31_inst : DFF_X1 port map( D => n8633, CK => CLK, Q => 
                           n_1578, QN => n4993);
   REGISTERS_reg_42_30_inst : DFF_X1 port map( D => n8632, CK => CLK, Q => 
                           n_1579, QN => n4992);
   REGISTERS_reg_42_29_inst : DFF_X1 port map( D => n8631, CK => CLK, Q => 
                           n_1580, QN => n4991);
   REGISTERS_reg_42_28_inst : DFF_X1 port map( D => n8630, CK => CLK, Q => 
                           n_1581, QN => n4990);
   REGISTERS_reg_42_27_inst : DFF_X1 port map( D => n8629, CK => CLK, Q => 
                           n_1582, QN => n4989);
   REGISTERS_reg_42_26_inst : DFF_X1 port map( D => n8628, CK => CLK, Q => 
                           n_1583, QN => n4988);
   REGISTERS_reg_42_25_inst : DFF_X1 port map( D => n8627, CK => CLK, Q => 
                           n_1584, QN => n4987);
   REGISTERS_reg_42_24_inst : DFF_X1 port map( D => n8626, CK => CLK, Q => 
                           n_1585, QN => n4986);
   REGISTERS_reg_42_23_inst : DFF_X1 port map( D => n8625, CK => CLK, Q => 
                           n_1586, QN => n4985);
   REGISTERS_reg_42_22_inst : DFF_X1 port map( D => n8624, CK => CLK, Q => 
                           n_1587, QN => n4984);
   REGISTERS_reg_42_21_inst : DFF_X1 port map( D => n8623, CK => CLK, Q => 
                           n_1588, QN => n4983);
   REGISTERS_reg_42_20_inst : DFF_X1 port map( D => n8622, CK => CLK, Q => 
                           n_1589, QN => n4982);
   REGISTERS_reg_42_19_inst : DFF_X1 port map( D => n8621, CK => CLK, Q => 
                           n_1590, QN => n4981);
   REGISTERS_reg_42_18_inst : DFF_X1 port map( D => n8620, CK => CLK, Q => 
                           n_1591, QN => n4980);
   REGISTERS_reg_42_17_inst : DFF_X1 port map( D => n8619, CK => CLK, Q => 
                           n_1592, QN => n4979);
   REGISTERS_reg_42_16_inst : DFF_X1 port map( D => n8618, CK => CLK, Q => 
                           n_1593, QN => n4978);
   REGISTERS_reg_42_15_inst : DFF_X1 port map( D => n8617, CK => CLK, Q => 
                           n_1594, QN => n4977);
   REGISTERS_reg_42_14_inst : DFF_X1 port map( D => n8616, CK => CLK, Q => 
                           n_1595, QN => n4976);
   REGISTERS_reg_42_13_inst : DFF_X1 port map( D => n8615, CK => CLK, Q => 
                           n_1596, QN => n4975);
   REGISTERS_reg_42_12_inst : DFF_X1 port map( D => n8614, CK => CLK, Q => 
                           n_1597, QN => n4974);
   REGISTERS_reg_42_11_inst : DFF_X1 port map( D => n8613, CK => CLK, Q => 
                           n_1598, QN => n4973);
   REGISTERS_reg_42_10_inst : DFF_X1 port map( D => n8612, CK => CLK, Q => 
                           n_1599, QN => n4972);
   REGISTERS_reg_42_9_inst : DFF_X1 port map( D => n8611, CK => CLK, Q => 
                           n_1600, QN => n4971);
   REGISTERS_reg_42_8_inst : DFF_X1 port map( D => n8610, CK => CLK, Q => 
                           n_1601, QN => n4970);
   REGISTERS_reg_42_7_inst : DFF_X1 port map( D => n8609, CK => CLK, Q => 
                           n_1602, QN => n4969);
   REGISTERS_reg_42_6_inst : DFF_X1 port map( D => n8608, CK => CLK, Q => 
                           n_1603, QN => n4968);
   REGISTERS_reg_42_5_inst : DFF_X1 port map( D => n8607, CK => CLK, Q => 
                           n_1604, QN => n4967);
   REGISTERS_reg_42_4_inst : DFF_X1 port map( D => n8606, CK => CLK, Q => 
                           n_1605, QN => n4966);
   REGISTERS_reg_42_3_inst : DFF_X1 port map( D => n8605, CK => CLK, Q => 
                           n_1606, QN => n4965);
   REGISTERS_reg_42_2_inst : DFF_X1 port map( D => n8604, CK => CLK, Q => 
                           n_1607, QN => n4964);
   REGISTERS_reg_42_1_inst : DFF_X1 port map( D => n8603, CK => CLK, Q => 
                           n_1608, QN => n4963);
   REGISTERS_reg_42_0_inst : DFF_X1 port map( D => n8602, CK => CLK, Q => 
                           n_1609, QN => n4962);
   REGISTERS_reg_43_31_inst : DFF_X1 port map( D => n8601, CK => CLK, Q => 
                           n_1610, QN => n4961);
   REGISTERS_reg_43_30_inst : DFF_X1 port map( D => n8600, CK => CLK, Q => 
                           n_1611, QN => n4960);
   REGISTERS_reg_43_29_inst : DFF_X1 port map( D => n8599, CK => CLK, Q => 
                           n_1612, QN => n4959);
   REGISTERS_reg_43_28_inst : DFF_X1 port map( D => n8598, CK => CLK, Q => 
                           n_1613, QN => n4958);
   REGISTERS_reg_43_27_inst : DFF_X1 port map( D => n8597, CK => CLK, Q => 
                           n_1614, QN => n4957);
   REGISTERS_reg_43_26_inst : DFF_X1 port map( D => n8596, CK => CLK, Q => 
                           n_1615, QN => n4956);
   REGISTERS_reg_43_25_inst : DFF_X1 port map( D => n8595, CK => CLK, Q => 
                           n_1616, QN => n4955);
   REGISTERS_reg_43_24_inst : DFF_X1 port map( D => n8594, CK => CLK, Q => 
                           n_1617, QN => n4954);
   REGISTERS_reg_43_23_inst : DFF_X1 port map( D => n8593, CK => CLK, Q => 
                           n_1618, QN => n4953);
   REGISTERS_reg_43_22_inst : DFF_X1 port map( D => n8592, CK => CLK, Q => 
                           n_1619, QN => n4952);
   REGISTERS_reg_43_21_inst : DFF_X1 port map( D => n8591, CK => CLK, Q => 
                           n_1620, QN => n4951);
   REGISTERS_reg_43_20_inst : DFF_X1 port map( D => n8590, CK => CLK, Q => 
                           n_1621, QN => n4950);
   REGISTERS_reg_43_19_inst : DFF_X1 port map( D => n8589, CK => CLK, Q => 
                           n_1622, QN => n4949);
   REGISTERS_reg_43_18_inst : DFF_X1 port map( D => n8588, CK => CLK, Q => 
                           n_1623, QN => n4948);
   REGISTERS_reg_43_17_inst : DFF_X1 port map( D => n8587, CK => CLK, Q => 
                           n_1624, QN => n4947);
   REGISTERS_reg_43_16_inst : DFF_X1 port map( D => n8586, CK => CLK, Q => 
                           n_1625, QN => n4946);
   REGISTERS_reg_43_15_inst : DFF_X1 port map( D => n8585, CK => CLK, Q => 
                           n_1626, QN => n4945);
   REGISTERS_reg_43_14_inst : DFF_X1 port map( D => n8584, CK => CLK, Q => 
                           n_1627, QN => n4944);
   REGISTERS_reg_43_13_inst : DFF_X1 port map( D => n8583, CK => CLK, Q => 
                           n_1628, QN => n4943);
   REGISTERS_reg_43_12_inst : DFF_X1 port map( D => n8582, CK => CLK, Q => 
                           n_1629, QN => n4942);
   REGISTERS_reg_43_11_inst : DFF_X1 port map( D => n8581, CK => CLK, Q => 
                           n_1630, QN => n4941);
   REGISTERS_reg_43_10_inst : DFF_X1 port map( D => n8580, CK => CLK, Q => 
                           n_1631, QN => n4940);
   REGISTERS_reg_43_9_inst : DFF_X1 port map( D => n8579, CK => CLK, Q => 
                           n_1632, QN => n4939);
   REGISTERS_reg_43_8_inst : DFF_X1 port map( D => n8578, CK => CLK, Q => 
                           n_1633, QN => n4938);
   REGISTERS_reg_43_7_inst : DFF_X1 port map( D => n8577, CK => CLK, Q => 
                           n_1634, QN => n4937);
   REGISTERS_reg_43_6_inst : DFF_X1 port map( D => n8576, CK => CLK, Q => 
                           n_1635, QN => n4936);
   REGISTERS_reg_43_5_inst : DFF_X1 port map( D => n8575, CK => CLK, Q => 
                           n_1636, QN => n4935);
   REGISTERS_reg_43_4_inst : DFF_X1 port map( D => n8574, CK => CLK, Q => 
                           n_1637, QN => n4934);
   REGISTERS_reg_43_3_inst : DFF_X1 port map( D => n8573, CK => CLK, Q => 
                           n_1638, QN => n4933);
   REGISTERS_reg_43_2_inst : DFF_X1 port map( D => n8572, CK => CLK, Q => 
                           n_1639, QN => n4932);
   REGISTERS_reg_43_1_inst : DFF_X1 port map( D => n8571, CK => CLK, Q => 
                           n_1640, QN => n4931);
   REGISTERS_reg_43_0_inst : DFF_X1 port map( D => n8570, CK => CLK, Q => 
                           n_1641, QN => n4930);
   REGISTERS_reg_44_31_inst : DFF_X1 port map( D => n8569, CK => CLK, Q => 
                           n_1642, QN => n4929);
   REGISTERS_reg_44_30_inst : DFF_X1 port map( D => n8568, CK => CLK, Q => 
                           n_1643, QN => n4928);
   REGISTERS_reg_44_29_inst : DFF_X1 port map( D => n8567, CK => CLK, Q => 
                           n_1644, QN => n4927);
   REGISTERS_reg_44_28_inst : DFF_X1 port map( D => n8566, CK => CLK, Q => 
                           n_1645, QN => n4926);
   REGISTERS_reg_44_27_inst : DFF_X1 port map( D => n8565, CK => CLK, Q => 
                           n_1646, QN => n4925);
   REGISTERS_reg_44_26_inst : DFF_X1 port map( D => n8564, CK => CLK, Q => 
                           n_1647, QN => n4924);
   REGISTERS_reg_44_25_inst : DFF_X1 port map( D => n8563, CK => CLK, Q => 
                           n_1648, QN => n4923);
   REGISTERS_reg_44_24_inst : DFF_X1 port map( D => n8562, CK => CLK, Q => 
                           n_1649, QN => n4922);
   REGISTERS_reg_44_23_inst : DFF_X1 port map( D => n8561, CK => CLK, Q => 
                           n_1650, QN => n4921);
   REGISTERS_reg_44_22_inst : DFF_X1 port map( D => n8560, CK => CLK, Q => 
                           n_1651, QN => n4920);
   REGISTERS_reg_44_21_inst : DFF_X1 port map( D => n8559, CK => CLK, Q => 
                           n_1652, QN => n4919);
   REGISTERS_reg_44_20_inst : DFF_X1 port map( D => n8558, CK => CLK, Q => 
                           n_1653, QN => n4918);
   REGISTERS_reg_44_19_inst : DFF_X1 port map( D => n8557, CK => CLK, Q => 
                           n_1654, QN => n4917);
   REGISTERS_reg_44_18_inst : DFF_X1 port map( D => n8556, CK => CLK, Q => 
                           n_1655, QN => n4916);
   REGISTERS_reg_44_17_inst : DFF_X1 port map( D => n8555, CK => CLK, Q => 
                           n_1656, QN => n4915);
   REGISTERS_reg_44_16_inst : DFF_X1 port map( D => n8554, CK => CLK, Q => 
                           n_1657, QN => n4914);
   REGISTERS_reg_44_15_inst : DFF_X1 port map( D => n8553, CK => CLK, Q => 
                           n_1658, QN => n4913);
   REGISTERS_reg_44_14_inst : DFF_X1 port map( D => n8552, CK => CLK, Q => 
                           n_1659, QN => n4912);
   REGISTERS_reg_44_13_inst : DFF_X1 port map( D => n8551, CK => CLK, Q => 
                           n_1660, QN => n4911);
   REGISTERS_reg_44_12_inst : DFF_X1 port map( D => n8550, CK => CLK, Q => 
                           n_1661, QN => n4910);
   REGISTERS_reg_44_11_inst : DFF_X1 port map( D => n8549, CK => CLK, Q => 
                           n_1662, QN => n4909);
   REGISTERS_reg_44_10_inst : DFF_X1 port map( D => n8548, CK => CLK, Q => 
                           n_1663, QN => n4908);
   REGISTERS_reg_44_9_inst : DFF_X1 port map( D => n8547, CK => CLK, Q => 
                           n_1664, QN => n4907);
   REGISTERS_reg_44_8_inst : DFF_X1 port map( D => n8546, CK => CLK, Q => 
                           n_1665, QN => n4906);
   REGISTERS_reg_44_7_inst : DFF_X1 port map( D => n8545, CK => CLK, Q => 
                           n_1666, QN => n4905);
   REGISTERS_reg_44_6_inst : DFF_X1 port map( D => n8544, CK => CLK, Q => 
                           n_1667, QN => n4904);
   REGISTERS_reg_44_5_inst : DFF_X1 port map( D => n8543, CK => CLK, Q => 
                           n_1668, QN => n4903);
   REGISTERS_reg_44_4_inst : DFF_X1 port map( D => n8542, CK => CLK, Q => 
                           n_1669, QN => n4902);
   REGISTERS_reg_44_3_inst : DFF_X1 port map( D => n8541, CK => CLK, Q => 
                           n_1670, QN => n4901);
   REGISTERS_reg_44_2_inst : DFF_X1 port map( D => n8540, CK => CLK, Q => 
                           n_1671, QN => n4900);
   REGISTERS_reg_44_1_inst : DFF_X1 port map( D => n8539, CK => CLK, Q => 
                           n_1672, QN => n4899);
   REGISTERS_reg_44_0_inst : DFF_X1 port map( D => n8538, CK => CLK, Q => 
                           n_1673, QN => n4898);
   REGISTERS_reg_45_31_inst : DFF_X1 port map( D => n8537, CK => CLK, Q => 
                           n6209, QN => n619);
   REGISTERS_reg_45_30_inst : DFF_X1 port map( D => n8536, CK => CLK, Q => 
                           n6208, QN => n622);
   REGISTERS_reg_45_29_inst : DFF_X1 port map( D => n8535, CK => CLK, Q => 
                           n6207, QN => n625);
   REGISTERS_reg_45_28_inst : DFF_X1 port map( D => n8534, CK => CLK, Q => 
                           n6206, QN => n628);
   REGISTERS_reg_45_27_inst : DFF_X1 port map( D => n8533, CK => CLK, Q => 
                           n6205, QN => n631);
   REGISTERS_reg_45_26_inst : DFF_X1 port map( D => n8532, CK => CLK, Q => 
                           n6204, QN => n634);
   REGISTERS_reg_45_25_inst : DFF_X1 port map( D => n8531, CK => CLK, Q => 
                           n6203, QN => n637);
   REGISTERS_reg_45_24_inst : DFF_X1 port map( D => n8530, CK => CLK, Q => 
                           n6202, QN => n640);
   REGISTERS_reg_45_23_inst : DFF_X1 port map( D => n8529, CK => CLK, Q => 
                           n6201, QN => n643);
   REGISTERS_reg_45_22_inst : DFF_X1 port map( D => n8528, CK => CLK, Q => 
                           n6200, QN => n646);
   REGISTERS_reg_45_21_inst : DFF_X1 port map( D => n8527, CK => CLK, Q => 
                           n6199, QN => n649);
   REGISTERS_reg_45_20_inst : DFF_X1 port map( D => n8526, CK => CLK, Q => 
                           n6198, QN => n652);
   REGISTERS_reg_45_19_inst : DFF_X1 port map( D => n8525, CK => CLK, Q => 
                           n6197, QN => n655);
   REGISTERS_reg_45_18_inst : DFF_X1 port map( D => n8524, CK => CLK, Q => 
                           n6196, QN => n658);
   REGISTERS_reg_45_17_inst : DFF_X1 port map( D => n8523, CK => CLK, Q => 
                           n6195, QN => n661);
   REGISTERS_reg_45_16_inst : DFF_X1 port map( D => n8522, CK => CLK, Q => 
                           n6194, QN => n664);
   REGISTERS_reg_45_15_inst : DFF_X1 port map( D => n8521, CK => CLK, Q => 
                           n6193, QN => n667);
   REGISTERS_reg_45_14_inst : DFF_X1 port map( D => n8520, CK => CLK, Q => 
                           n6192, QN => n670);
   REGISTERS_reg_45_13_inst : DFF_X1 port map( D => n8519, CK => CLK, Q => 
                           n6191, QN => n673);
   REGISTERS_reg_45_12_inst : DFF_X1 port map( D => n8518, CK => CLK, Q => 
                           n6190, QN => n676);
   REGISTERS_reg_45_11_inst : DFF_X1 port map( D => n8517, CK => CLK, Q => 
                           n6189, QN => n679);
   REGISTERS_reg_45_10_inst : DFF_X1 port map( D => n8516, CK => CLK, Q => 
                           n6188, QN => n682);
   REGISTERS_reg_45_9_inst : DFF_X1 port map( D => n8515, CK => CLK, Q => n6187
                           , QN => n685);
   REGISTERS_reg_45_8_inst : DFF_X1 port map( D => n8514, CK => CLK, Q => n6186
                           , QN => n688);
   REGISTERS_reg_45_7_inst : DFF_X1 port map( D => n8513, CK => CLK, Q => n6185
                           , QN => n691);
   REGISTERS_reg_45_6_inst : DFF_X1 port map( D => n8512, CK => CLK, Q => n6184
                           , QN => n694);
   REGISTERS_reg_45_5_inst : DFF_X1 port map( D => n8511, CK => CLK, Q => n6183
                           , QN => n697);
   REGISTERS_reg_45_4_inst : DFF_X1 port map( D => n8510, CK => CLK, Q => n6182
                           , QN => n700);
   REGISTERS_reg_45_3_inst : DFF_X1 port map( D => n8509, CK => CLK, Q => n6181
                           , QN => n703);
   REGISTERS_reg_45_2_inst : DFF_X1 port map( D => n8508, CK => CLK, Q => n6180
                           , QN => n706);
   REGISTERS_reg_45_1_inst : DFF_X1 port map( D => n8507, CK => CLK, Q => n6179
                           , QN => n709);
   REGISTERS_reg_45_0_inst : DFF_X1 port map( D => n8506, CK => CLK, Q => n6178
                           , QN => n712);
   REGISTERS_reg_46_31_inst : DFF_X1 port map( D => n8505, CK => CLK, Q => 
                           n6177, QN => n195);
   REGISTERS_reg_46_30_inst : DFF_X1 port map( D => n8504, CK => CLK, Q => 
                           n6176, QN => n198);
   REGISTERS_reg_46_29_inst : DFF_X1 port map( D => n8503, CK => CLK, Q => 
                           n6175, QN => n201);
   REGISTERS_reg_46_28_inst : DFF_X1 port map( D => n8502, CK => CLK, Q => 
                           n6174, QN => n204);
   REGISTERS_reg_46_27_inst : DFF_X1 port map( D => n8501, CK => CLK, Q => 
                           n6173, QN => n207);
   REGISTERS_reg_46_26_inst : DFF_X1 port map( D => n8500, CK => CLK, Q => 
                           n6172, QN => n210);
   REGISTERS_reg_46_25_inst : DFF_X1 port map( D => n8499, CK => CLK, Q => 
                           n6171, QN => n213);
   REGISTERS_reg_46_24_inst : DFF_X1 port map( D => n8498, CK => CLK, Q => 
                           n6170, QN => n216);
   REGISTERS_reg_46_23_inst : DFF_X1 port map( D => n8497, CK => CLK, Q => 
                           n6169, QN => n219);
   REGISTERS_reg_46_22_inst : DFF_X1 port map( D => n8496, CK => CLK, Q => 
                           n6168, QN => n222);
   REGISTERS_reg_46_21_inst : DFF_X1 port map( D => n8495, CK => CLK, Q => 
                           n6167, QN => n225);
   REGISTERS_reg_46_20_inst : DFF_X1 port map( D => n8494, CK => CLK, Q => 
                           n6166, QN => n228);
   REGISTERS_reg_46_19_inst : DFF_X1 port map( D => n8493, CK => CLK, Q => 
                           n6165, QN => n231);
   REGISTERS_reg_46_18_inst : DFF_X1 port map( D => n8492, CK => CLK, Q => 
                           n6164, QN => n234);
   REGISTERS_reg_46_17_inst : DFF_X1 port map( D => n8491, CK => CLK, Q => 
                           n6163, QN => n237);
   REGISTERS_reg_46_16_inst : DFF_X1 port map( D => n8490, CK => CLK, Q => 
                           n6162, QN => n240);
   REGISTERS_reg_46_15_inst : DFF_X1 port map( D => n8489, CK => CLK, Q => 
                           n6161, QN => n243);
   REGISTERS_reg_46_14_inst : DFF_X1 port map( D => n8488, CK => CLK, Q => 
                           n6160, QN => n246);
   REGISTERS_reg_46_13_inst : DFF_X1 port map( D => n8487, CK => CLK, Q => 
                           n6159, QN => n249);
   REGISTERS_reg_46_12_inst : DFF_X1 port map( D => n8486, CK => CLK, Q => 
                           n6158, QN => n252);
   REGISTERS_reg_46_11_inst : DFF_X1 port map( D => n8485, CK => CLK, Q => 
                           n6157, QN => n255);
   REGISTERS_reg_46_10_inst : DFF_X1 port map( D => n8484, CK => CLK, Q => 
                           n6156, QN => n258);
   REGISTERS_reg_46_9_inst : DFF_X1 port map( D => n8483, CK => CLK, Q => n6155
                           , QN => n261);
   REGISTERS_reg_46_8_inst : DFF_X1 port map( D => n8482, CK => CLK, Q => n6154
                           , QN => n264);
   REGISTERS_reg_46_7_inst : DFF_X1 port map( D => n8481, CK => CLK, Q => n6153
                           , QN => n267);
   REGISTERS_reg_46_6_inst : DFF_X1 port map( D => n8480, CK => CLK, Q => n6152
                           , QN => n270);
   REGISTERS_reg_46_5_inst : DFF_X1 port map( D => n8479, CK => CLK, Q => n6151
                           , QN => n273);
   REGISTERS_reg_46_4_inst : DFF_X1 port map( D => n8478, CK => CLK, Q => n6150
                           , QN => n276);
   REGISTERS_reg_46_3_inst : DFF_X1 port map( D => n8477, CK => CLK, Q => n6149
                           , QN => n279);
   REGISTERS_reg_46_2_inst : DFF_X1 port map( D => n8476, CK => CLK, Q => n6148
                           , QN => n282);
   REGISTERS_reg_46_1_inst : DFF_X1 port map( D => n8475, CK => CLK, Q => n6147
                           , QN => n285);
   REGISTERS_reg_46_0_inst : DFF_X1 port map( D => n8474, CK => CLK, Q => n6146
                           , QN => n288);
   REGISTERS_reg_47_31_inst : DFF_X1 port map( D => n8473, CK => CLK, Q => n715
                           , QN => n5690);
   REGISTERS_reg_47_30_inst : DFF_X1 port map( D => n8472, CK => CLK, Q => n718
                           , QN => n5680);
   REGISTERS_reg_47_29_inst : DFF_X1 port map( D => n8471, CK => CLK, Q => n721
                           , QN => n5670);
   REGISTERS_reg_47_28_inst : DFF_X1 port map( D => n8470, CK => CLK, Q => n724
                           , QN => n5660);
   REGISTERS_reg_47_27_inst : DFF_X1 port map( D => n8469, CK => CLK, Q => n727
                           , QN => n5650);
   REGISTERS_reg_47_26_inst : DFF_X1 port map( D => n8468, CK => CLK, Q => n730
                           , QN => n5640);
   REGISTERS_reg_47_25_inst : DFF_X1 port map( D => n8467, CK => CLK, Q => n733
                           , QN => n5630);
   REGISTERS_reg_47_24_inst : DFF_X1 port map( D => n8466, CK => CLK, Q => n736
                           , QN => n5620);
   REGISTERS_reg_47_23_inst : DFF_X1 port map( D => n8465, CK => CLK, Q => n739
                           , QN => n5610);
   REGISTERS_reg_47_22_inst : DFF_X1 port map( D => n8464, CK => CLK, Q => n742
                           , QN => n5600);
   REGISTERS_reg_47_21_inst : DFF_X1 port map( D => n8463, CK => CLK, Q => n745
                           , QN => n5590);
   REGISTERS_reg_47_20_inst : DFF_X1 port map( D => n8462, CK => CLK, Q => n748
                           , QN => n5580);
   REGISTERS_reg_47_19_inst : DFF_X1 port map( D => n8461, CK => CLK, Q => n751
                           , QN => n5570);
   REGISTERS_reg_47_18_inst : DFF_X1 port map( D => n8460, CK => CLK, Q => n754
                           , QN => n5560);
   REGISTERS_reg_47_17_inst : DFF_X1 port map( D => n8459, CK => CLK, Q => n757
                           , QN => n5550);
   REGISTERS_reg_47_16_inst : DFF_X1 port map( D => n8458, CK => CLK, Q => n760
                           , QN => n5540);
   REGISTERS_reg_47_15_inst : DFF_X1 port map( D => n8457, CK => CLK, Q => n763
                           , QN => n5530);
   REGISTERS_reg_47_14_inst : DFF_X1 port map( D => n8456, CK => CLK, Q => n766
                           , QN => n5520);
   REGISTERS_reg_47_13_inst : DFF_X1 port map( D => n8455, CK => CLK, Q => n769
                           , QN => n5510);
   REGISTERS_reg_47_12_inst : DFF_X1 port map( D => n8454, CK => CLK, Q => n772
                           , QN => n5500);
   REGISTERS_reg_47_11_inst : DFF_X1 port map( D => n8453, CK => CLK, Q => n775
                           , QN => n5490);
   REGISTERS_reg_47_10_inst : DFF_X1 port map( D => n8452, CK => CLK, Q => n778
                           , QN => n5480);
   REGISTERS_reg_47_9_inst : DFF_X1 port map( D => n8451, CK => CLK, Q => n781,
                           QN => n5470);
   REGISTERS_reg_47_8_inst : DFF_X1 port map( D => n8450, CK => CLK, Q => n784,
                           QN => n5460);
   REGISTERS_reg_47_7_inst : DFF_X1 port map( D => n8449, CK => CLK, Q => n787,
                           QN => n5450);
   REGISTERS_reg_47_6_inst : DFF_X1 port map( D => n8448, CK => CLK, Q => n790,
                           QN => n5440);
   REGISTERS_reg_47_5_inst : DFF_X1 port map( D => n8447, CK => CLK, Q => n793,
                           QN => n5430);
   REGISTERS_reg_47_4_inst : DFF_X1 port map( D => n8446, CK => CLK, Q => n796,
                           QN => n5420);
   REGISTERS_reg_47_3_inst : DFF_X1 port map( D => n8445, CK => CLK, Q => n799,
                           QN => n5410);
   REGISTERS_reg_47_2_inst : DFF_X1 port map( D => n8444, CK => CLK, Q => n802,
                           QN => n5400);
   REGISTERS_reg_47_1_inst : DFF_X1 port map( D => n8443, CK => CLK, Q => n805,
                           QN => n5390);
   REGISTERS_reg_47_0_inst : DFF_X1 port map( D => n8442, CK => CLK, Q => n808,
                           QN => n5380);
   REGISTERS_reg_48_31_inst : DFF_X1 port map( D => n8441, CK => CLK, Q => n291
                           , QN => n5691);
   REGISTERS_reg_48_30_inst : DFF_X1 port map( D => n8440, CK => CLK, Q => n294
                           , QN => n5681);
   REGISTERS_reg_48_29_inst : DFF_X1 port map( D => n8439, CK => CLK, Q => n297
                           , QN => n5671);
   REGISTERS_reg_48_28_inst : DFF_X1 port map( D => n8438, CK => CLK, Q => n300
                           , QN => n5661);
   REGISTERS_reg_48_27_inst : DFF_X1 port map( D => n8437, CK => CLK, Q => n303
                           , QN => n5651);
   REGISTERS_reg_48_26_inst : DFF_X1 port map( D => n8436, CK => CLK, Q => n306
                           , QN => n5641);
   REGISTERS_reg_48_25_inst : DFF_X1 port map( D => n8435, CK => CLK, Q => n309
                           , QN => n5631);
   REGISTERS_reg_48_24_inst : DFF_X1 port map( D => n8434, CK => CLK, Q => n312
                           , QN => n5621);
   REGISTERS_reg_48_23_inst : DFF_X1 port map( D => n8433, CK => CLK, Q => n315
                           , QN => n5611);
   REGISTERS_reg_48_22_inst : DFF_X1 port map( D => n8432, CK => CLK, Q => n318
                           , QN => n5601);
   REGISTERS_reg_48_21_inst : DFF_X1 port map( D => n8431, CK => CLK, Q => n321
                           , QN => n5591);
   REGISTERS_reg_48_20_inst : DFF_X1 port map( D => n8430, CK => CLK, Q => n324
                           , QN => n5581);
   REGISTERS_reg_48_19_inst : DFF_X1 port map( D => n8429, CK => CLK, Q => n327
                           , QN => n5571);
   REGISTERS_reg_48_18_inst : DFF_X1 port map( D => n8428, CK => CLK, Q => n330
                           , QN => n5561);
   REGISTERS_reg_48_17_inst : DFF_X1 port map( D => n8427, CK => CLK, Q => n333
                           , QN => n5551);
   REGISTERS_reg_48_16_inst : DFF_X1 port map( D => n8426, CK => CLK, Q => n336
                           , QN => n5541);
   REGISTERS_reg_48_15_inst : DFF_X1 port map( D => n8425, CK => CLK, Q => n339
                           , QN => n5531);
   REGISTERS_reg_48_14_inst : DFF_X1 port map( D => n8424, CK => CLK, Q => n342
                           , QN => n5521);
   REGISTERS_reg_48_13_inst : DFF_X1 port map( D => n8423, CK => CLK, Q => n345
                           , QN => n5511);
   REGISTERS_reg_48_12_inst : DFF_X1 port map( D => n8422, CK => CLK, Q => n348
                           , QN => n5501);
   REGISTERS_reg_48_11_inst : DFF_X1 port map( D => n8421, CK => CLK, Q => n351
                           , QN => n5491);
   REGISTERS_reg_48_10_inst : DFF_X1 port map( D => n8420, CK => CLK, Q => n354
                           , QN => n5481);
   REGISTERS_reg_48_9_inst : DFF_X1 port map( D => n8419, CK => CLK, Q => n357,
                           QN => n5471);
   REGISTERS_reg_48_8_inst : DFF_X1 port map( D => n8418, CK => CLK, Q => n360,
                           QN => n5461);
   REGISTERS_reg_48_7_inst : DFF_X1 port map( D => n8417, CK => CLK, Q => n363,
                           QN => n5451);
   REGISTERS_reg_48_6_inst : DFF_X1 port map( D => n8416, CK => CLK, Q => n366,
                           QN => n5441);
   REGISTERS_reg_48_5_inst : DFF_X1 port map( D => n8415, CK => CLK, Q => n369,
                           QN => n5431);
   REGISTERS_reg_48_4_inst : DFF_X1 port map( D => n8414, CK => CLK, Q => n372,
                           QN => n5421);
   REGISTERS_reg_48_3_inst : DFF_X1 port map( D => n8413, CK => CLK, Q => n375,
                           QN => n5411);
   REGISTERS_reg_48_2_inst : DFF_X1 port map( D => n8412, CK => CLK, Q => n378,
                           QN => n5401);
   REGISTERS_reg_48_1_inst : DFF_X1 port map( D => n8411, CK => CLK, Q => n381,
                           QN => n5391);
   REGISTERS_reg_48_0_inst : DFF_X1 port map( D => n8410, CK => CLK, Q => n384,
                           QN => n5381);
   REGISTERS_reg_49_31_inst : DFF_X1 port map( D => n8409, CK => CLK, Q => 
                           n6145, QN => n969);
   REGISTERS_reg_49_30_inst : DFF_X1 port map( D => n8408, CK => CLK, Q => 
                           n6144, QN => n970);
   REGISTERS_reg_49_29_inst : DFF_X1 port map( D => n8407, CK => CLK, Q => 
                           n6143, QN => n971);
   REGISTERS_reg_49_28_inst : DFF_X1 port map( D => n8406, CK => CLK, Q => 
                           n6142, QN => n972);
   REGISTERS_reg_49_27_inst : DFF_X1 port map( D => n8405, CK => CLK, Q => 
                           n6141, QN => n973);
   REGISTERS_reg_49_26_inst : DFF_X1 port map( D => n8404, CK => CLK, Q => 
                           n6140, QN => n974);
   REGISTERS_reg_49_25_inst : DFF_X1 port map( D => n8403, CK => CLK, Q => 
                           n6139, QN => n975);
   REGISTERS_reg_49_24_inst : DFF_X1 port map( D => n8402, CK => CLK, Q => 
                           n6138, QN => n976);
   REGISTERS_reg_49_23_inst : DFF_X1 port map( D => n8401, CK => CLK, Q => 
                           n6137, QN => n977);
   REGISTERS_reg_49_22_inst : DFF_X1 port map( D => n8400, CK => CLK, Q => 
                           n6136, QN => n978);
   REGISTERS_reg_49_21_inst : DFF_X1 port map( D => n8399, CK => CLK, Q => 
                           n6135, QN => n979);
   REGISTERS_reg_49_20_inst : DFF_X1 port map( D => n8398, CK => CLK, Q => 
                           n6134, QN => n980);
   REGISTERS_reg_49_19_inst : DFF_X1 port map( D => n8397, CK => CLK, Q => 
                           n6133, QN => n981);
   REGISTERS_reg_49_18_inst : DFF_X1 port map( D => n8396, CK => CLK, Q => 
                           n6132, QN => n982);
   REGISTERS_reg_49_17_inst : DFF_X1 port map( D => n8395, CK => CLK, Q => 
                           n6131, QN => n983);
   REGISTERS_reg_49_16_inst : DFF_X1 port map( D => n8394, CK => CLK, Q => 
                           n6130, QN => n984);
   REGISTERS_reg_49_15_inst : DFF_X1 port map( D => n8393, CK => CLK, Q => 
                           n6129, QN => n985);
   REGISTERS_reg_49_14_inst : DFF_X1 port map( D => n8392, CK => CLK, Q => 
                           n6128, QN => n986);
   REGISTERS_reg_49_13_inst : DFF_X1 port map( D => n8391, CK => CLK, Q => 
                           n6127, QN => n987);
   REGISTERS_reg_49_12_inst : DFF_X1 port map( D => n8390, CK => CLK, Q => 
                           n6126, QN => n988);
   REGISTERS_reg_49_11_inst : DFF_X1 port map( D => n8389, CK => CLK, Q => 
                           n6125, QN => n989);
   REGISTERS_reg_49_10_inst : DFF_X1 port map( D => n8388, CK => CLK, Q => 
                           n6124, QN => n990);
   REGISTERS_reg_49_9_inst : DFF_X1 port map( D => n8387, CK => CLK, Q => n6123
                           , QN => n991);
   REGISTERS_reg_49_8_inst : DFF_X1 port map( D => n8386, CK => CLK, Q => n6122
                           , QN => n992);
   REGISTERS_reg_49_7_inst : DFF_X1 port map( D => n8385, CK => CLK, Q => n6121
                           , QN => n993);
   REGISTERS_reg_49_6_inst : DFF_X1 port map( D => n8384, CK => CLK, Q => n6120
                           , QN => n994);
   REGISTERS_reg_49_5_inst : DFF_X1 port map( D => n8383, CK => CLK, Q => n6119
                           , QN => n995);
   REGISTERS_reg_49_4_inst : DFF_X1 port map( D => n8382, CK => CLK, Q => n6118
                           , QN => n996);
   REGISTERS_reg_49_3_inst : DFF_X1 port map( D => n8381, CK => CLK, Q => n6117
                           , QN => n997);
   REGISTERS_reg_49_2_inst : DFF_X1 port map( D => n8380, CK => CLK, Q => n6116
                           , QN => n998);
   REGISTERS_reg_49_1_inst : DFF_X1 port map( D => n8379, CK => CLK, Q => n6115
                           , QN => n999);
   REGISTERS_reg_49_0_inst : DFF_X1 port map( D => n8378, CK => CLK, Q => n6114
                           , QN => n1000);
   REGISTERS_reg_50_31_inst : DFF_X1 port map( D => n8377, CK => CLK, Q => 
                           n6113, QN => n1321);
   REGISTERS_reg_50_30_inst : DFF_X1 port map( D => n8376, CK => CLK, Q => 
                           n6112, QN => n1322);
   REGISTERS_reg_50_29_inst : DFF_X1 port map( D => n8375, CK => CLK, Q => 
                           n6111, QN => n1323);
   REGISTERS_reg_50_28_inst : DFF_X1 port map( D => n8374, CK => CLK, Q => 
                           n6110, QN => n1324);
   REGISTERS_reg_50_27_inst : DFF_X1 port map( D => n8373, CK => CLK, Q => 
                           n6109, QN => n1325);
   REGISTERS_reg_50_26_inst : DFF_X1 port map( D => n8372, CK => CLK, Q => 
                           n6108, QN => n1326);
   REGISTERS_reg_50_25_inst : DFF_X1 port map( D => n8371, CK => CLK, Q => 
                           n6107, QN => n1327);
   REGISTERS_reg_50_24_inst : DFF_X1 port map( D => n8370, CK => CLK, Q => 
                           n6106, QN => n1328);
   REGISTERS_reg_50_23_inst : DFF_X1 port map( D => n8369, CK => CLK, Q => 
                           n6105, QN => n1329);
   REGISTERS_reg_50_22_inst : DFF_X1 port map( D => n8368, CK => CLK, Q => 
                           n6104, QN => n1330);
   REGISTERS_reg_50_21_inst : DFF_X1 port map( D => n8367, CK => CLK, Q => 
                           n6103, QN => n1331);
   REGISTERS_reg_50_20_inst : DFF_X1 port map( D => n8366, CK => CLK, Q => 
                           n6102, QN => n1332);
   REGISTERS_reg_50_19_inst : DFF_X1 port map( D => n8365, CK => CLK, Q => 
                           n6101, QN => n1333);
   REGISTERS_reg_50_18_inst : DFF_X1 port map( D => n8364, CK => CLK, Q => 
                           n6100, QN => n1334);
   REGISTERS_reg_50_17_inst : DFF_X1 port map( D => n8363, CK => CLK, Q => 
                           n6099, QN => n1335);
   REGISTERS_reg_50_16_inst : DFF_X1 port map( D => n8362, CK => CLK, Q => 
                           n6098, QN => n1336);
   REGISTERS_reg_50_15_inst : DFF_X1 port map( D => n8361, CK => CLK, Q => 
                           n6097, QN => n1337);
   REGISTERS_reg_50_14_inst : DFF_X1 port map( D => n8360, CK => CLK, Q => 
                           n6096, QN => n1338);
   REGISTERS_reg_50_13_inst : DFF_X1 port map( D => n8359, CK => CLK, Q => 
                           n6095, QN => n1339);
   REGISTERS_reg_50_12_inst : DFF_X1 port map( D => n8358, CK => CLK, Q => 
                           n6094, QN => n1340);
   REGISTERS_reg_50_11_inst : DFF_X1 port map( D => n8357, CK => CLK, Q => 
                           n6093, QN => n1341);
   REGISTERS_reg_50_10_inst : DFF_X1 port map( D => n8356, CK => CLK, Q => 
                           n6092, QN => n1342);
   REGISTERS_reg_50_9_inst : DFF_X1 port map( D => n8355, CK => CLK, Q => n6091
                           , QN => n1343);
   REGISTERS_reg_50_8_inst : DFF_X1 port map( D => n8354, CK => CLK, Q => n6090
                           , QN => n1344);
   REGISTERS_reg_50_7_inst : DFF_X1 port map( D => n8353, CK => CLK, Q => n6089
                           , QN => n1345);
   REGISTERS_reg_50_6_inst : DFF_X1 port map( D => n8352, CK => CLK, Q => n6088
                           , QN => n1346);
   REGISTERS_reg_50_5_inst : DFF_X1 port map( D => n8351, CK => CLK, Q => n6087
                           , QN => n1347);
   REGISTERS_reg_50_4_inst : DFF_X1 port map( D => n8350, CK => CLK, Q => n6086
                           , QN => n1348);
   REGISTERS_reg_50_3_inst : DFF_X1 port map( D => n8349, CK => CLK, Q => n6085
                           , QN => n1349);
   REGISTERS_reg_50_2_inst : DFF_X1 port map( D => n8348, CK => CLK, Q => n6084
                           , QN => n1350);
   REGISTERS_reg_50_1_inst : DFF_X1 port map( D => n8347, CK => CLK, Q => n6083
                           , QN => n1351);
   REGISTERS_reg_50_0_inst : DFF_X1 port map( D => n8346, CK => CLK, Q => n6082
                           , QN => n1352);
   REGISTERS_reg_51_31_inst : DFF_X1 port map( D => n8345, CK => CLK, Q => 
                           n_1674, QN => n4897);
   REGISTERS_reg_51_30_inst : DFF_X1 port map( D => n8344, CK => CLK, Q => 
                           n_1675, QN => n4896);
   REGISTERS_reg_51_29_inst : DFF_X1 port map( D => n8343, CK => CLK, Q => 
                           n_1676, QN => n4895);
   REGISTERS_reg_51_28_inst : DFF_X1 port map( D => n8342, CK => CLK, Q => 
                           n_1677, QN => n4894);
   REGISTERS_reg_51_27_inst : DFF_X1 port map( D => n8341, CK => CLK, Q => 
                           n_1678, QN => n4893);
   REGISTERS_reg_51_26_inst : DFF_X1 port map( D => n8340, CK => CLK, Q => 
                           n_1679, QN => n4892);
   REGISTERS_reg_51_25_inst : DFF_X1 port map( D => n8339, CK => CLK, Q => 
                           n_1680, QN => n4891);
   REGISTERS_reg_51_24_inst : DFF_X1 port map( D => n8338, CK => CLK, Q => 
                           n_1681, QN => n4890);
   REGISTERS_reg_51_23_inst : DFF_X1 port map( D => n8337, CK => CLK, Q => 
                           n_1682, QN => n4889);
   REGISTERS_reg_51_22_inst : DFF_X1 port map( D => n8336, CK => CLK, Q => 
                           n_1683, QN => n4888);
   REGISTERS_reg_51_21_inst : DFF_X1 port map( D => n8335, CK => CLK, Q => 
                           n_1684, QN => n4887);
   REGISTERS_reg_51_20_inst : DFF_X1 port map( D => n8334, CK => CLK, Q => 
                           n_1685, QN => n4886);
   REGISTERS_reg_51_19_inst : DFF_X1 port map( D => n8333, CK => CLK, Q => 
                           n_1686, QN => n4885);
   REGISTERS_reg_51_18_inst : DFF_X1 port map( D => n8332, CK => CLK, Q => 
                           n_1687, QN => n4884);
   REGISTERS_reg_51_17_inst : DFF_X1 port map( D => n8331, CK => CLK, Q => 
                           n_1688, QN => n4883);
   REGISTERS_reg_51_16_inst : DFF_X1 port map( D => n8330, CK => CLK, Q => 
                           n_1689, QN => n4882);
   REGISTERS_reg_51_15_inst : DFF_X1 port map( D => n8329, CK => CLK, Q => 
                           n_1690, QN => n4881);
   REGISTERS_reg_51_14_inst : DFF_X1 port map( D => n8328, CK => CLK, Q => 
                           n_1691, QN => n4880);
   REGISTERS_reg_51_13_inst : DFF_X1 port map( D => n8327, CK => CLK, Q => 
                           n_1692, QN => n4879);
   REGISTERS_reg_51_12_inst : DFF_X1 port map( D => n8326, CK => CLK, Q => 
                           n_1693, QN => n4878);
   REGISTERS_reg_51_11_inst : DFF_X1 port map( D => n8325, CK => CLK, Q => 
                           n_1694, QN => n4877);
   REGISTERS_reg_51_10_inst : DFF_X1 port map( D => n8324, CK => CLK, Q => 
                           n_1695, QN => n4876);
   REGISTERS_reg_51_9_inst : DFF_X1 port map( D => n8323, CK => CLK, Q => 
                           n_1696, QN => n4875);
   REGISTERS_reg_51_8_inst : DFF_X1 port map( D => n8322, CK => CLK, Q => 
                           n_1697, QN => n4874);
   REGISTERS_reg_51_7_inst : DFF_X1 port map( D => n8321, CK => CLK, Q => 
                           n_1698, QN => n4873);
   REGISTERS_reg_51_6_inst : DFF_X1 port map( D => n8320, CK => CLK, Q => 
                           n_1699, QN => n4872);
   REGISTERS_reg_51_5_inst : DFF_X1 port map( D => n8319, CK => CLK, Q => 
                           n_1700, QN => n4871);
   REGISTERS_reg_51_4_inst : DFF_X1 port map( D => n8318, CK => CLK, Q => 
                           n_1701, QN => n4870);
   REGISTERS_reg_51_3_inst : DFF_X1 port map( D => n8317, CK => CLK, Q => 
                           n_1702, QN => n4869);
   REGISTERS_reg_51_2_inst : DFF_X1 port map( D => n8316, CK => CLK, Q => 
                           n_1703, QN => n4868);
   REGISTERS_reg_51_1_inst : DFF_X1 port map( D => n8315, CK => CLK, Q => 
                           n_1704, QN => n4867);
   REGISTERS_reg_51_0_inst : DFF_X1 port map( D => n8314, CK => CLK, Q => 
                           n_1705, QN => n4866);
   REGISTERS_reg_52_31_inst : DFF_X1 port map( D => n8313, CK => CLK, Q => 
                           n_1706, QN => n4865);
   REGISTERS_reg_52_30_inst : DFF_X1 port map( D => n8312, CK => CLK, Q => 
                           n_1707, QN => n4864);
   REGISTERS_reg_52_29_inst : DFF_X1 port map( D => n8311, CK => CLK, Q => 
                           n_1708, QN => n4863);
   REGISTERS_reg_52_28_inst : DFF_X1 port map( D => n8310, CK => CLK, Q => 
                           n_1709, QN => n4862);
   REGISTERS_reg_52_27_inst : DFF_X1 port map( D => n8309, CK => CLK, Q => 
                           n_1710, QN => n4861);
   REGISTERS_reg_52_26_inst : DFF_X1 port map( D => n8308, CK => CLK, Q => 
                           n_1711, QN => n4860);
   REGISTERS_reg_52_25_inst : DFF_X1 port map( D => n8307, CK => CLK, Q => 
                           n_1712, QN => n4859);
   REGISTERS_reg_52_24_inst : DFF_X1 port map( D => n8306, CK => CLK, Q => 
                           n_1713, QN => n4858);
   REGISTERS_reg_52_23_inst : DFF_X1 port map( D => n8305, CK => CLK, Q => 
                           n_1714, QN => n4857);
   REGISTERS_reg_52_22_inst : DFF_X1 port map( D => n8304, CK => CLK, Q => 
                           n_1715, QN => n4856);
   REGISTERS_reg_52_21_inst : DFF_X1 port map( D => n8303, CK => CLK, Q => 
                           n_1716, QN => n4855);
   REGISTERS_reg_52_20_inst : DFF_X1 port map( D => n8302, CK => CLK, Q => 
                           n_1717, QN => n4854);
   REGISTERS_reg_52_19_inst : DFF_X1 port map( D => n8301, CK => CLK, Q => 
                           n_1718, QN => n4853);
   REGISTERS_reg_52_18_inst : DFF_X1 port map( D => n8300, CK => CLK, Q => 
                           n_1719, QN => n4852);
   REGISTERS_reg_52_17_inst : DFF_X1 port map( D => n8299, CK => CLK, Q => 
                           n_1720, QN => n4851);
   REGISTERS_reg_52_16_inst : DFF_X1 port map( D => n8298, CK => CLK, Q => 
                           n_1721, QN => n4850);
   REGISTERS_reg_52_15_inst : DFF_X1 port map( D => n8297, CK => CLK, Q => 
                           n_1722, QN => n4849);
   REGISTERS_reg_52_14_inst : DFF_X1 port map( D => n8296, CK => CLK, Q => 
                           n_1723, QN => n4848);
   REGISTERS_reg_52_13_inst : DFF_X1 port map( D => n8295, CK => CLK, Q => 
                           n_1724, QN => n4847);
   REGISTERS_reg_52_12_inst : DFF_X1 port map( D => n8294, CK => CLK, Q => 
                           n_1725, QN => n4846);
   REGISTERS_reg_52_11_inst : DFF_X1 port map( D => n8293, CK => CLK, Q => 
                           n_1726, QN => n4845);
   REGISTERS_reg_52_10_inst : DFF_X1 port map( D => n8292, CK => CLK, Q => 
                           n_1727, QN => n4844);
   REGISTERS_reg_52_9_inst : DFF_X1 port map( D => n8291, CK => CLK, Q => 
                           n_1728, QN => n4843);
   REGISTERS_reg_52_8_inst : DFF_X1 port map( D => n8290, CK => CLK, Q => 
                           n_1729, QN => n4842);
   REGISTERS_reg_52_7_inst : DFF_X1 port map( D => n8289, CK => CLK, Q => 
                           n_1730, QN => n4841);
   REGISTERS_reg_52_6_inst : DFF_X1 port map( D => n8288, CK => CLK, Q => 
                           n_1731, QN => n4840);
   REGISTERS_reg_52_5_inst : DFF_X1 port map( D => n8287, CK => CLK, Q => 
                           n_1732, QN => n4839);
   REGISTERS_reg_52_4_inst : DFF_X1 port map( D => n8286, CK => CLK, Q => 
                           n_1733, QN => n4838);
   REGISTERS_reg_52_3_inst : DFF_X1 port map( D => n8285, CK => CLK, Q => 
                           n_1734, QN => n4837);
   REGISTERS_reg_52_2_inst : DFF_X1 port map( D => n8284, CK => CLK, Q => 
                           n_1735, QN => n4836);
   REGISTERS_reg_52_1_inst : DFF_X1 port map( D => n8283, CK => CLK, Q => 
                           n_1736, QN => n4835);
   REGISTERS_reg_52_0_inst : DFF_X1 port map( D => n8282, CK => CLK, Q => 
                           n_1737, QN => n4834);
   REGISTERS_reg_53_31_inst : DFF_X1 port map( D => n8281, CK => CLK, Q => 
                           n_1738, QN => n4833);
   REGISTERS_reg_53_30_inst : DFF_X1 port map( D => n8280, CK => CLK, Q => 
                           n_1739, QN => n4832);
   REGISTERS_reg_53_29_inst : DFF_X1 port map( D => n8279, CK => CLK, Q => 
                           n_1740, QN => n4831);
   REGISTERS_reg_53_28_inst : DFF_X1 port map( D => n8278, CK => CLK, Q => 
                           n_1741, QN => n4830);
   REGISTERS_reg_53_27_inst : DFF_X1 port map( D => n8277, CK => CLK, Q => 
                           n_1742, QN => n4829);
   REGISTERS_reg_53_26_inst : DFF_X1 port map( D => n8276, CK => CLK, Q => 
                           n_1743, QN => n4828);
   REGISTERS_reg_53_25_inst : DFF_X1 port map( D => n8275, CK => CLK, Q => 
                           n_1744, QN => n4827);
   REGISTERS_reg_53_24_inst : DFF_X1 port map( D => n8274, CK => CLK, Q => 
                           n_1745, QN => n4826);
   REGISTERS_reg_53_23_inst : DFF_X1 port map( D => n8273, CK => CLK, Q => 
                           n_1746, QN => n4825);
   REGISTERS_reg_53_22_inst : DFF_X1 port map( D => n8272, CK => CLK, Q => 
                           n_1747, QN => n4824);
   REGISTERS_reg_53_21_inst : DFF_X1 port map( D => n8271, CK => CLK, Q => 
                           n_1748, QN => n4823);
   REGISTERS_reg_53_20_inst : DFF_X1 port map( D => n8270, CK => CLK, Q => 
                           n_1749, QN => n4822);
   REGISTERS_reg_53_19_inst : DFF_X1 port map( D => n8269, CK => CLK, Q => 
                           n_1750, QN => n4821);
   REGISTERS_reg_53_18_inst : DFF_X1 port map( D => n8268, CK => CLK, Q => 
                           n_1751, QN => n4820);
   REGISTERS_reg_53_17_inst : DFF_X1 port map( D => n8267, CK => CLK, Q => 
                           n_1752, QN => n4819);
   REGISTERS_reg_53_16_inst : DFF_X1 port map( D => n8266, CK => CLK, Q => 
                           n_1753, QN => n4818);
   REGISTERS_reg_53_15_inst : DFF_X1 port map( D => n8265, CK => CLK, Q => 
                           n_1754, QN => n4817);
   REGISTERS_reg_53_14_inst : DFF_X1 port map( D => n8264, CK => CLK, Q => 
                           n_1755, QN => n4816);
   REGISTERS_reg_53_13_inst : DFF_X1 port map( D => n8263, CK => CLK, Q => 
                           n_1756, QN => n4815);
   REGISTERS_reg_53_12_inst : DFF_X1 port map( D => n8262, CK => CLK, Q => 
                           n_1757, QN => n4814);
   REGISTERS_reg_53_11_inst : DFF_X1 port map( D => n8261, CK => CLK, Q => 
                           n_1758, QN => n4813);
   REGISTERS_reg_53_10_inst : DFF_X1 port map( D => n8260, CK => CLK, Q => 
                           n_1759, QN => n4812);
   REGISTERS_reg_53_9_inst : DFF_X1 port map( D => n8259, CK => CLK, Q => 
                           n_1760, QN => n4811);
   REGISTERS_reg_53_8_inst : DFF_X1 port map( D => n8258, CK => CLK, Q => 
                           n_1761, QN => n4810);
   REGISTERS_reg_53_7_inst : DFF_X1 port map( D => n8257, CK => CLK, Q => 
                           n_1762, QN => n4809);
   REGISTERS_reg_53_6_inst : DFF_X1 port map( D => n8256, CK => CLK, Q => 
                           n_1763, QN => n4808);
   REGISTERS_reg_53_5_inst : DFF_X1 port map( D => n8255, CK => CLK, Q => 
                           n_1764, QN => n4807);
   REGISTERS_reg_53_4_inst : DFF_X1 port map( D => n8254, CK => CLK, Q => 
                           n_1765, QN => n4806);
   REGISTERS_reg_53_3_inst : DFF_X1 port map( D => n8253, CK => CLK, Q => 
                           n_1766, QN => n4805);
   REGISTERS_reg_53_2_inst : DFF_X1 port map( D => n8252, CK => CLK, Q => 
                           n_1767, QN => n4804);
   REGISTERS_reg_53_1_inst : DFF_X1 port map( D => n8251, CK => CLK, Q => 
                           n_1768, QN => n4803);
   REGISTERS_reg_53_0_inst : DFF_X1 port map( D => n8250, CK => CLK, Q => 
                           n_1769, QN => n4802);
   REGISTERS_reg_54_31_inst : DFF_X1 port map( D => n8249, CK => CLK, Q => 
                           n_1770, QN => n5688);
   REGISTERS_reg_54_30_inst : DFF_X1 port map( D => n8248, CK => CLK, Q => 
                           n_1771, QN => n5678);
   REGISTERS_reg_54_29_inst : DFF_X1 port map( D => n8247, CK => CLK, Q => 
                           n_1772, QN => n5668);
   REGISTERS_reg_54_28_inst : DFF_X1 port map( D => n8246, CK => CLK, Q => 
                           n_1773, QN => n5658);
   REGISTERS_reg_54_27_inst : DFF_X1 port map( D => n8245, CK => CLK, Q => 
                           n_1774, QN => n5648);
   REGISTERS_reg_54_26_inst : DFF_X1 port map( D => n8244, CK => CLK, Q => 
                           n_1775, QN => n5638);
   REGISTERS_reg_54_25_inst : DFF_X1 port map( D => n8243, CK => CLK, Q => 
                           n_1776, QN => n5628);
   REGISTERS_reg_54_24_inst : DFF_X1 port map( D => n8242, CK => CLK, Q => 
                           n_1777, QN => n5618);
   REGISTERS_reg_54_23_inst : DFF_X1 port map( D => n8241, CK => CLK, Q => 
                           n_1778, QN => n5608);
   REGISTERS_reg_54_22_inst : DFF_X1 port map( D => n8240, CK => CLK, Q => 
                           n_1779, QN => n5598);
   REGISTERS_reg_54_21_inst : DFF_X1 port map( D => n8239, CK => CLK, Q => 
                           n_1780, QN => n5588);
   REGISTERS_reg_54_20_inst : DFF_X1 port map( D => n8238, CK => CLK, Q => 
                           n_1781, QN => n5578);
   REGISTERS_reg_54_19_inst : DFF_X1 port map( D => n8237, CK => CLK, Q => 
                           n_1782, QN => n5568);
   REGISTERS_reg_54_18_inst : DFF_X1 port map( D => n8236, CK => CLK, Q => 
                           n_1783, QN => n5558);
   REGISTERS_reg_54_17_inst : DFF_X1 port map( D => n8235, CK => CLK, Q => 
                           n_1784, QN => n5548);
   REGISTERS_reg_54_16_inst : DFF_X1 port map( D => n8234, CK => CLK, Q => 
                           n_1785, QN => n5538);
   REGISTERS_reg_54_15_inst : DFF_X1 port map( D => n8233, CK => CLK, Q => 
                           n_1786, QN => n5528);
   REGISTERS_reg_54_14_inst : DFF_X1 port map( D => n8232, CK => CLK, Q => 
                           n_1787, QN => n5518);
   REGISTERS_reg_54_13_inst : DFF_X1 port map( D => n8231, CK => CLK, Q => 
                           n_1788, QN => n5508);
   REGISTERS_reg_54_12_inst : DFF_X1 port map( D => n8230, CK => CLK, Q => 
                           n_1789, QN => n5498);
   REGISTERS_reg_54_11_inst : DFF_X1 port map( D => n8229, CK => CLK, Q => 
                           n_1790, QN => n5488);
   REGISTERS_reg_54_10_inst : DFF_X1 port map( D => n8228, CK => CLK, Q => 
                           n_1791, QN => n5478);
   REGISTERS_reg_54_9_inst : DFF_X1 port map( D => n8227, CK => CLK, Q => 
                           n_1792, QN => n5468);
   REGISTERS_reg_54_8_inst : DFF_X1 port map( D => n8226, CK => CLK, Q => 
                           n_1793, QN => n5458);
   REGISTERS_reg_54_7_inst : DFF_X1 port map( D => n8225, CK => CLK, Q => 
                           n_1794, QN => n5448);
   REGISTERS_reg_54_6_inst : DFF_X1 port map( D => n8224, CK => CLK, Q => 
                           n_1795, QN => n5438);
   REGISTERS_reg_54_5_inst : DFF_X1 port map( D => n8223, CK => CLK, Q => 
                           n_1796, QN => n5428);
   REGISTERS_reg_54_4_inst : DFF_X1 port map( D => n8222, CK => CLK, Q => 
                           n_1797, QN => n5418);
   REGISTERS_reg_54_3_inst : DFF_X1 port map( D => n8221, CK => CLK, Q => 
                           n_1798, QN => n5408);
   REGISTERS_reg_54_2_inst : DFF_X1 port map( D => n8220, CK => CLK, Q => 
                           n_1799, QN => n5398);
   REGISTERS_reg_54_1_inst : DFF_X1 port map( D => n8219, CK => CLK, Q => 
                           n_1800, QN => n5388);
   REGISTERS_reg_54_0_inst : DFF_X1 port map( D => n8218, CK => CLK, Q => 
                           n_1801, QN => n5378);
   REGISTERS_reg_55_31_inst : DFF_X1 port map( D => n8217, CK => CLK, Q => 
                           n_1802, QN => n5689);
   REGISTERS_reg_55_30_inst : DFF_X1 port map( D => n8216, CK => CLK, Q => 
                           n_1803, QN => n5679);
   REGISTERS_reg_55_29_inst : DFF_X1 port map( D => n8215, CK => CLK, Q => 
                           n_1804, QN => n5669);
   REGISTERS_reg_55_28_inst : DFF_X1 port map( D => n8214, CK => CLK, Q => 
                           n_1805, QN => n5659);
   REGISTERS_reg_55_27_inst : DFF_X1 port map( D => n8213, CK => CLK, Q => 
                           n_1806, QN => n5649);
   REGISTERS_reg_55_26_inst : DFF_X1 port map( D => n8212, CK => CLK, Q => 
                           n_1807, QN => n5639);
   REGISTERS_reg_55_25_inst : DFF_X1 port map( D => n8211, CK => CLK, Q => 
                           n_1808, QN => n5629);
   REGISTERS_reg_55_24_inst : DFF_X1 port map( D => n8210, CK => CLK, Q => 
                           n_1809, QN => n5619);
   REGISTERS_reg_55_23_inst : DFF_X1 port map( D => n8209, CK => CLK, Q => 
                           n_1810, QN => n5609);
   REGISTERS_reg_55_22_inst : DFF_X1 port map( D => n8208, CK => CLK, Q => 
                           n_1811, QN => n5599);
   REGISTERS_reg_55_21_inst : DFF_X1 port map( D => n8207, CK => CLK, Q => 
                           n_1812, QN => n5589);
   REGISTERS_reg_55_20_inst : DFF_X1 port map( D => n8206, CK => CLK, Q => 
                           n_1813, QN => n5579);
   REGISTERS_reg_55_19_inst : DFF_X1 port map( D => n8205, CK => CLK, Q => 
                           n_1814, QN => n5569);
   REGISTERS_reg_55_18_inst : DFF_X1 port map( D => n8204, CK => CLK, Q => 
                           n_1815, QN => n5559);
   REGISTERS_reg_55_17_inst : DFF_X1 port map( D => n8203, CK => CLK, Q => 
                           n_1816, QN => n5549);
   REGISTERS_reg_55_16_inst : DFF_X1 port map( D => n8202, CK => CLK, Q => 
                           n_1817, QN => n5539);
   REGISTERS_reg_55_15_inst : DFF_X1 port map( D => n8201, CK => CLK, Q => 
                           n_1818, QN => n5529);
   REGISTERS_reg_55_14_inst : DFF_X1 port map( D => n8200, CK => CLK, Q => 
                           n_1819, QN => n5519);
   REGISTERS_reg_55_13_inst : DFF_X1 port map( D => n8199, CK => CLK, Q => 
                           n_1820, QN => n5509);
   REGISTERS_reg_55_12_inst : DFF_X1 port map( D => n8198, CK => CLK, Q => 
                           n_1821, QN => n5499);
   REGISTERS_reg_55_11_inst : DFF_X1 port map( D => n8197, CK => CLK, Q => 
                           n_1822, QN => n5489);
   REGISTERS_reg_55_10_inst : DFF_X1 port map( D => n8196, CK => CLK, Q => 
                           n_1823, QN => n5479);
   REGISTERS_reg_55_9_inst : DFF_X1 port map( D => n8195, CK => CLK, Q => 
                           n_1824, QN => n5469);
   REGISTERS_reg_55_8_inst : DFF_X1 port map( D => n8194, CK => CLK, Q => 
                           n_1825, QN => n5459);
   REGISTERS_reg_55_7_inst : DFF_X1 port map( D => n8193, CK => CLK, Q => 
                           n_1826, QN => n5449);
   REGISTERS_reg_55_6_inst : DFF_X1 port map( D => n8192, CK => CLK, Q => 
                           n_1827, QN => n5439);
   REGISTERS_reg_55_5_inst : DFF_X1 port map( D => n8191, CK => CLK, Q => 
                           n_1828, QN => n5429);
   REGISTERS_reg_55_4_inst : DFF_X1 port map( D => n8190, CK => CLK, Q => 
                           n_1829, QN => n5419);
   REGISTERS_reg_55_3_inst : DFF_X1 port map( D => n8189, CK => CLK, Q => 
                           n_1830, QN => n5409);
   REGISTERS_reg_55_2_inst : DFF_X1 port map( D => n8188, CK => CLK, Q => 
                           n_1831, QN => n5399);
   REGISTERS_reg_55_1_inst : DFF_X1 port map( D => n8187, CK => CLK, Q => 
                           n_1832, QN => n5389);
   REGISTERS_reg_55_0_inst : DFF_X1 port map( D => n8186, CK => CLK, Q => 
                           n_1833, QN => n5379);
   REGISTERS_reg_56_31_inst : DFF_X1 port map( D => n8185, CK => CLK, Q => 
                           n6081, QN => n1097);
   REGISTERS_reg_56_30_inst : DFF_X1 port map( D => n8184, CK => CLK, Q => 
                           n6080, QN => n1098);
   REGISTERS_reg_56_29_inst : DFF_X1 port map( D => n8183, CK => CLK, Q => 
                           n6079, QN => n1099);
   REGISTERS_reg_56_28_inst : DFF_X1 port map( D => n8182, CK => CLK, Q => 
                           n6078, QN => n1100);
   REGISTERS_reg_56_27_inst : DFF_X1 port map( D => n8181, CK => CLK, Q => 
                           n6077, QN => n1101);
   REGISTERS_reg_56_26_inst : DFF_X1 port map( D => n8180, CK => CLK, Q => 
                           n6076, QN => n1102);
   REGISTERS_reg_56_25_inst : DFF_X1 port map( D => n8179, CK => CLK, Q => 
                           n6075, QN => n1103);
   REGISTERS_reg_56_24_inst : DFF_X1 port map( D => n8178, CK => CLK, Q => 
                           n6074, QN => n1104);
   REGISTERS_reg_56_23_inst : DFF_X1 port map( D => n8177, CK => CLK, Q => 
                           n6073, QN => n1105);
   REGISTERS_reg_56_22_inst : DFF_X1 port map( D => n8176, CK => CLK, Q => 
                           n6072, QN => n1106);
   REGISTERS_reg_56_21_inst : DFF_X1 port map( D => n8175, CK => CLK, Q => 
                           n6071, QN => n1107);
   REGISTERS_reg_56_20_inst : DFF_X1 port map( D => n8174, CK => CLK, Q => 
                           n6070, QN => n1108);
   REGISTERS_reg_56_19_inst : DFF_X1 port map( D => n8173, CK => CLK, Q => 
                           n6069, QN => n1109);
   REGISTERS_reg_56_18_inst : DFF_X1 port map( D => n8172, CK => CLK, Q => 
                           n6068, QN => n1110);
   REGISTERS_reg_56_17_inst : DFF_X1 port map( D => n8171, CK => CLK, Q => 
                           n6067, QN => n1111);
   REGISTERS_reg_56_16_inst : DFF_X1 port map( D => n8170, CK => CLK, Q => 
                           n6066, QN => n1112);
   REGISTERS_reg_56_15_inst : DFF_X1 port map( D => n8169, CK => CLK, Q => 
                           n6065, QN => n1113);
   REGISTERS_reg_56_14_inst : DFF_X1 port map( D => n8168, CK => CLK, Q => 
                           n6064, QN => n1114);
   REGISTERS_reg_56_13_inst : DFF_X1 port map( D => n8167, CK => CLK, Q => 
                           n6063, QN => n1115);
   REGISTERS_reg_56_12_inst : DFF_X1 port map( D => n8166, CK => CLK, Q => 
                           n6062, QN => n1116);
   REGISTERS_reg_56_11_inst : DFF_X1 port map( D => n8165, CK => CLK, Q => 
                           n6061, QN => n1117);
   REGISTERS_reg_56_10_inst : DFF_X1 port map( D => n8164, CK => CLK, Q => 
                           n6060, QN => n1118);
   REGISTERS_reg_56_9_inst : DFF_X1 port map( D => n8163, CK => CLK, Q => n6059
                           , QN => n1119);
   REGISTERS_reg_56_8_inst : DFF_X1 port map( D => n8162, CK => CLK, Q => n6058
                           , QN => n1120);
   REGISTERS_reg_56_7_inst : DFF_X1 port map( D => n8161, CK => CLK, Q => n6057
                           , QN => n1121);
   REGISTERS_reg_56_6_inst : DFF_X1 port map( D => n8160, CK => CLK, Q => n6056
                           , QN => n1122);
   REGISTERS_reg_56_5_inst : DFF_X1 port map( D => n8159, CK => CLK, Q => n6055
                           , QN => n1123);
   REGISTERS_reg_56_4_inst : DFF_X1 port map( D => n8158, CK => CLK, Q => n6054
                           , QN => n1124);
   REGISTERS_reg_56_3_inst : DFF_X1 port map( D => n8157, CK => CLK, Q => n6053
                           , QN => n1125);
   REGISTERS_reg_56_2_inst : DFF_X1 port map( D => n8156, CK => CLK, Q => n6052
                           , QN => n1126);
   REGISTERS_reg_56_1_inst : DFF_X1 port map( D => n8155, CK => CLK, Q => n6051
                           , QN => n1127);
   REGISTERS_reg_56_0_inst : DFF_X1 port map( D => n8154, CK => CLK, Q => n6050
                           , QN => n1128);
   REGISTERS_reg_57_31_inst : DFF_X1 port map( D => n8153, CK => CLK, Q => 
                           n6049, QN => n1129);
   REGISTERS_reg_57_30_inst : DFF_X1 port map( D => n8152, CK => CLK, Q => 
                           n6048, QN => n1130);
   REGISTERS_reg_57_29_inst : DFF_X1 port map( D => n8151, CK => CLK, Q => 
                           n6047, QN => n1131);
   REGISTERS_reg_57_28_inst : DFF_X1 port map( D => n8150, CK => CLK, Q => 
                           n6046, QN => n1132);
   REGISTERS_reg_57_27_inst : DFF_X1 port map( D => n8149, CK => CLK, Q => 
                           n6045, QN => n1133);
   REGISTERS_reg_57_26_inst : DFF_X1 port map( D => n8148, CK => CLK, Q => 
                           n6044, QN => n1134);
   REGISTERS_reg_57_25_inst : DFF_X1 port map( D => n8147, CK => CLK, Q => 
                           n6043, QN => n1135);
   REGISTERS_reg_57_24_inst : DFF_X1 port map( D => n8146, CK => CLK, Q => 
                           n6042, QN => n1136);
   REGISTERS_reg_57_23_inst : DFF_X1 port map( D => n8145, CK => CLK, Q => 
                           n6041, QN => n1137);
   REGISTERS_reg_57_22_inst : DFF_X1 port map( D => n8144, CK => CLK, Q => 
                           n6040, QN => n1138);
   REGISTERS_reg_57_21_inst : DFF_X1 port map( D => n8143, CK => CLK, Q => 
                           n6039, QN => n1139);
   REGISTERS_reg_57_20_inst : DFF_X1 port map( D => n8142, CK => CLK, Q => 
                           n6038, QN => n1140);
   REGISTERS_reg_57_19_inst : DFF_X1 port map( D => n8141, CK => CLK, Q => 
                           n6037, QN => n1141);
   REGISTERS_reg_57_18_inst : DFF_X1 port map( D => n8140, CK => CLK, Q => 
                           n6036, QN => n1142);
   REGISTERS_reg_57_17_inst : DFF_X1 port map( D => n8139, CK => CLK, Q => 
                           n6035, QN => n1143);
   REGISTERS_reg_57_16_inst : DFF_X1 port map( D => n8138, CK => CLK, Q => 
                           n6034, QN => n1144);
   REGISTERS_reg_57_15_inst : DFF_X1 port map( D => n8137, CK => CLK, Q => 
                           n6033, QN => n1145);
   REGISTERS_reg_57_14_inst : DFF_X1 port map( D => n8136, CK => CLK, Q => 
                           n6032, QN => n1146);
   REGISTERS_reg_57_13_inst : DFF_X1 port map( D => n8135, CK => CLK, Q => 
                           n6031, QN => n1147);
   REGISTERS_reg_57_12_inst : DFF_X1 port map( D => n8134, CK => CLK, Q => 
                           n6030, QN => n1148);
   REGISTERS_reg_57_11_inst : DFF_X1 port map( D => n8133, CK => CLK, Q => 
                           n6029, QN => n1149);
   REGISTERS_reg_57_10_inst : DFF_X1 port map( D => n8132, CK => CLK, Q => 
                           n6028, QN => n1150);
   REGISTERS_reg_57_9_inst : DFF_X1 port map( D => n8131, CK => CLK, Q => n6027
                           , QN => n1151);
   REGISTERS_reg_57_8_inst : DFF_X1 port map( D => n8130, CK => CLK, Q => n6026
                           , QN => n1152);
   REGISTERS_reg_57_7_inst : DFF_X1 port map( D => n8129, CK => CLK, Q => n6025
                           , QN => n1153);
   REGISTERS_reg_57_6_inst : DFF_X1 port map( D => n8128, CK => CLK, Q => n6024
                           , QN => n1154);
   REGISTERS_reg_57_5_inst : DFF_X1 port map( D => n8127, CK => CLK, Q => n6023
                           , QN => n1155);
   REGISTERS_reg_57_4_inst : DFF_X1 port map( D => n8126, CK => CLK, Q => n6022
                           , QN => n1156);
   REGISTERS_reg_57_3_inst : DFF_X1 port map( D => n8125, CK => CLK, Q => n6021
                           , QN => n1157);
   REGISTERS_reg_57_2_inst : DFF_X1 port map( D => n8124, CK => CLK, Q => n6020
                           , QN => n1158);
   REGISTERS_reg_57_1_inst : DFF_X1 port map( D => n8123, CK => CLK, Q => n6019
                           , QN => n1159);
   REGISTERS_reg_57_0_inst : DFF_X1 port map( D => n8122, CK => CLK, Q => n6018
                           , QN => n1160);
   REGISTERS_reg_58_31_inst : DFF_X1 port map( D => n8121, CK => CLK, Q => 
                           n6017, QN => n1001);
   REGISTERS_reg_58_30_inst : DFF_X1 port map( D => n8120, CK => CLK, Q => 
                           n6016, QN => n1002);
   REGISTERS_reg_58_29_inst : DFF_X1 port map( D => n8119, CK => CLK, Q => 
                           n6015, QN => n1003);
   REGISTERS_reg_58_28_inst : DFF_X1 port map( D => n8118, CK => CLK, Q => 
                           n6014, QN => n1004);
   REGISTERS_reg_58_27_inst : DFF_X1 port map( D => n8117, CK => CLK, Q => 
                           n6013, QN => n1005);
   REGISTERS_reg_58_26_inst : DFF_X1 port map( D => n8116, CK => CLK, Q => 
                           n6012, QN => n1006);
   REGISTERS_reg_58_25_inst : DFF_X1 port map( D => n8115, CK => CLK, Q => 
                           n6011, QN => n1007);
   REGISTERS_reg_58_24_inst : DFF_X1 port map( D => n8114, CK => CLK, Q => 
                           n6010, QN => n1008);
   REGISTERS_reg_58_23_inst : DFF_X1 port map( D => n8113, CK => CLK, Q => 
                           n6009, QN => n1009);
   REGISTERS_reg_58_22_inst : DFF_X1 port map( D => n8112, CK => CLK, Q => 
                           n6008, QN => n1010);
   REGISTERS_reg_58_21_inst : DFF_X1 port map( D => n8111, CK => CLK, Q => 
                           n6007, QN => n1011);
   REGISTERS_reg_58_20_inst : DFF_X1 port map( D => n8110, CK => CLK, Q => 
                           n6006, QN => n1012);
   REGISTERS_reg_58_19_inst : DFF_X1 port map( D => n8109, CK => CLK, Q => 
                           n6005, QN => n1013);
   REGISTERS_reg_58_18_inst : DFF_X1 port map( D => n8108, CK => CLK, Q => 
                           n6004, QN => n1014);
   REGISTERS_reg_58_17_inst : DFF_X1 port map( D => n8107, CK => CLK, Q => 
                           n6003, QN => n1015);
   REGISTERS_reg_58_16_inst : DFF_X1 port map( D => n8106, CK => CLK, Q => 
                           n6002, QN => n1016);
   REGISTERS_reg_58_15_inst : DFF_X1 port map( D => n8105, CK => CLK, Q => 
                           n6001, QN => n1017);
   REGISTERS_reg_58_14_inst : DFF_X1 port map( D => n8104, CK => CLK, Q => 
                           n6000, QN => n1018);
   REGISTERS_reg_58_13_inst : DFF_X1 port map( D => n8103, CK => CLK, Q => 
                           n5999, QN => n1019);
   REGISTERS_reg_58_12_inst : DFF_X1 port map( D => n8102, CK => CLK, Q => 
                           n5998, QN => n1020);
   REGISTERS_reg_58_11_inst : DFF_X1 port map( D => n8101, CK => CLK, Q => 
                           n5997, QN => n1021);
   REGISTERS_reg_58_10_inst : DFF_X1 port map( D => n8100, CK => CLK, Q => 
                           n5996, QN => n1022);
   REGISTERS_reg_58_9_inst : DFF_X1 port map( D => n8099, CK => CLK, Q => n5995
                           , QN => n1023);
   REGISTERS_reg_58_8_inst : DFF_X1 port map( D => n8098, CK => CLK, Q => n5994
                           , QN => n1024);
   REGISTERS_reg_58_7_inst : DFF_X1 port map( D => n8097, CK => CLK, Q => n5993
                           , QN => n1025);
   REGISTERS_reg_58_6_inst : DFF_X1 port map( D => n8096, CK => CLK, Q => n5992
                           , QN => n1026);
   REGISTERS_reg_58_5_inst : DFF_X1 port map( D => n8095, CK => CLK, Q => n5991
                           , QN => n1027);
   REGISTERS_reg_58_4_inst : DFF_X1 port map( D => n8094, CK => CLK, Q => n5990
                           , QN => n1028);
   REGISTERS_reg_58_3_inst : DFF_X1 port map( D => n8093, CK => CLK, Q => n5989
                           , QN => n1029);
   REGISTERS_reg_58_2_inst : DFF_X1 port map( D => n8092, CK => CLK, Q => n5988
                           , QN => n1030);
   REGISTERS_reg_58_1_inst : DFF_X1 port map( D => n8091, CK => CLK, Q => n5987
                           , QN => n1031);
   REGISTERS_reg_58_0_inst : DFF_X1 port map( D => n8090, CK => CLK, Q => n5986
                           , QN => n1032);
   REGISTERS_reg_59_31_inst : DFF_X1 port map( D => n8089, CK => CLK, Q => 
                           n5985, QN => n1353);
   REGISTERS_reg_59_30_inst : DFF_X1 port map( D => n8088, CK => CLK, Q => 
                           n5984, QN => n1354);
   REGISTERS_reg_59_29_inst : DFF_X1 port map( D => n8087, CK => CLK, Q => 
                           n5983, QN => n1355);
   REGISTERS_reg_59_28_inst : DFF_X1 port map( D => n8086, CK => CLK, Q => 
                           n5982, QN => n1356);
   REGISTERS_reg_59_27_inst : DFF_X1 port map( D => n8085, CK => CLK, Q => 
                           n5981, QN => n1357);
   REGISTERS_reg_59_26_inst : DFF_X1 port map( D => n8084, CK => CLK, Q => 
                           n5980, QN => n1358);
   REGISTERS_reg_59_25_inst : DFF_X1 port map( D => n8083, CK => CLK, Q => 
                           n5979, QN => n1359);
   REGISTERS_reg_59_24_inst : DFF_X1 port map( D => n8082, CK => CLK, Q => 
                           n5978, QN => n1360);
   REGISTERS_reg_59_23_inst : DFF_X1 port map( D => n8081, CK => CLK, Q => 
                           n5977, QN => n1361);
   REGISTERS_reg_59_22_inst : DFF_X1 port map( D => n8080, CK => CLK, Q => 
                           n5976, QN => n1362);
   REGISTERS_reg_59_21_inst : DFF_X1 port map( D => n8079, CK => CLK, Q => 
                           n5975, QN => n1363);
   REGISTERS_reg_59_20_inst : DFF_X1 port map( D => n8078, CK => CLK, Q => 
                           n5974, QN => n1364);
   REGISTERS_reg_59_19_inst : DFF_X1 port map( D => n8077, CK => CLK, Q => 
                           n5973, QN => n1365);
   REGISTERS_reg_59_18_inst : DFF_X1 port map( D => n8076, CK => CLK, Q => 
                           n5972, QN => n1366);
   REGISTERS_reg_59_17_inst : DFF_X1 port map( D => n8075, CK => CLK, Q => 
                           n5971, QN => n1367);
   REGISTERS_reg_59_16_inst : DFF_X1 port map( D => n8074, CK => CLK, Q => 
                           n5970, QN => n1368);
   REGISTERS_reg_59_15_inst : DFF_X1 port map( D => n8073, CK => CLK, Q => 
                           n5969, QN => n1369);
   REGISTERS_reg_59_14_inst : DFF_X1 port map( D => n8072, CK => CLK, Q => 
                           n5968, QN => n1370);
   REGISTERS_reg_59_13_inst : DFF_X1 port map( D => n8071, CK => CLK, Q => 
                           n5967, QN => n1371);
   REGISTERS_reg_59_12_inst : DFF_X1 port map( D => n8070, CK => CLK, Q => 
                           n5966, QN => n1372);
   REGISTERS_reg_59_11_inst : DFF_X1 port map( D => n8069, CK => CLK, Q => 
                           n5965, QN => n1373);
   REGISTERS_reg_59_10_inst : DFF_X1 port map( D => n8068, CK => CLK, Q => 
                           n5964, QN => n1374);
   REGISTERS_reg_59_9_inst : DFF_X1 port map( D => n8067, CK => CLK, Q => n5963
                           , QN => n1375);
   REGISTERS_reg_59_8_inst : DFF_X1 port map( D => n8066, CK => CLK, Q => n5962
                           , QN => n1376);
   REGISTERS_reg_59_7_inst : DFF_X1 port map( D => n8065, CK => CLK, Q => n5961
                           , QN => n1377);
   REGISTERS_reg_59_6_inst : DFF_X1 port map( D => n8064, CK => CLK, Q => n5960
                           , QN => n1378);
   REGISTERS_reg_59_5_inst : DFF_X1 port map( D => n8063, CK => CLK, Q => n5959
                           , QN => n1379);
   REGISTERS_reg_59_4_inst : DFF_X1 port map( D => n8062, CK => CLK, Q => n5958
                           , QN => n1380);
   REGISTERS_reg_59_3_inst : DFF_X1 port map( D => n8061, CK => CLK, Q => n5957
                           , QN => n1381);
   REGISTERS_reg_59_2_inst : DFF_X1 port map( D => n8060, CK => CLK, Q => n5956
                           , QN => n1382);
   REGISTERS_reg_59_1_inst : DFF_X1 port map( D => n8059, CK => CLK, Q => n5955
                           , QN => n1383);
   REGISTERS_reg_59_0_inst : DFF_X1 port map( D => n8058, CK => CLK, Q => n5954
                           , QN => n1384);
   REGISTERS_reg_60_31_inst : DFF_X1 port map( D => n8057, CK => CLK, Q => 
                           n_1834, QN => n4801);
   REGISTERS_reg_60_30_inst : DFF_X1 port map( D => n8056, CK => CLK, Q => 
                           n_1835, QN => n4800);
   REGISTERS_reg_60_29_inst : DFF_X1 port map( D => n8055, CK => CLK, Q => 
                           n_1836, QN => n4799);
   REGISTERS_reg_60_28_inst : DFF_X1 port map( D => n8054, CK => CLK, Q => 
                           n_1837, QN => n4798);
   REGISTERS_reg_60_27_inst : DFF_X1 port map( D => n8053, CK => CLK, Q => 
                           n_1838, QN => n4797);
   REGISTERS_reg_60_26_inst : DFF_X1 port map( D => n8052, CK => CLK, Q => 
                           n_1839, QN => n4796);
   REGISTERS_reg_60_25_inst : DFF_X1 port map( D => n8051, CK => CLK, Q => 
                           n_1840, QN => n4795);
   REGISTERS_reg_60_24_inst : DFF_X1 port map( D => n8050, CK => CLK, Q => 
                           n_1841, QN => n4794);
   REGISTERS_reg_60_23_inst : DFF_X1 port map( D => n8049, CK => CLK, Q => 
                           n_1842, QN => n4793);
   REGISTERS_reg_60_22_inst : DFF_X1 port map( D => n8048, CK => CLK, Q => 
                           n_1843, QN => n4792);
   REGISTERS_reg_60_21_inst : DFF_X1 port map( D => n8047, CK => CLK, Q => 
                           n_1844, QN => n4791);
   REGISTERS_reg_60_20_inst : DFF_X1 port map( D => n8046, CK => CLK, Q => 
                           n_1845, QN => n4790);
   REGISTERS_reg_60_19_inst : DFF_X1 port map( D => n8045, CK => CLK, Q => 
                           n_1846, QN => n4789);
   REGISTERS_reg_60_18_inst : DFF_X1 port map( D => n8044, CK => CLK, Q => 
                           n_1847, QN => n4788);
   REGISTERS_reg_60_17_inst : DFF_X1 port map( D => n8043, CK => CLK, Q => 
                           n_1848, QN => n4787);
   REGISTERS_reg_60_16_inst : DFF_X1 port map( D => n8042, CK => CLK, Q => 
                           n_1849, QN => n4786);
   REGISTERS_reg_60_15_inst : DFF_X1 port map( D => n8041, CK => CLK, Q => 
                           n_1850, QN => n4785);
   REGISTERS_reg_60_14_inst : DFF_X1 port map( D => n8040, CK => CLK, Q => 
                           n_1851, QN => n4784);
   REGISTERS_reg_60_13_inst : DFF_X1 port map( D => n8039, CK => CLK, Q => 
                           n_1852, QN => n4783);
   REGISTERS_reg_60_12_inst : DFF_X1 port map( D => n8038, CK => CLK, Q => 
                           n_1853, QN => n4782);
   REGISTERS_reg_60_11_inst : DFF_X1 port map( D => n8037, CK => CLK, Q => 
                           n_1854, QN => n4781);
   REGISTERS_reg_60_10_inst : DFF_X1 port map( D => n8036, CK => CLK, Q => 
                           n_1855, QN => n4780);
   REGISTERS_reg_60_9_inst : DFF_X1 port map( D => n8035, CK => CLK, Q => 
                           n_1856, QN => n4779);
   REGISTERS_reg_60_8_inst : DFF_X1 port map( D => n8034, CK => CLK, Q => 
                           n_1857, QN => n4778);
   REGISTERS_reg_60_7_inst : DFF_X1 port map( D => n8033, CK => CLK, Q => 
                           n_1858, QN => n4777);
   REGISTERS_reg_60_6_inst : DFF_X1 port map( D => n8032, CK => CLK, Q => 
                           n_1859, QN => n4776);
   REGISTERS_reg_60_5_inst : DFF_X1 port map( D => n8031, CK => CLK, Q => 
                           n_1860, QN => n4775);
   REGISTERS_reg_60_4_inst : DFF_X1 port map( D => n8030, CK => CLK, Q => 
                           n_1861, QN => n4774);
   REGISTERS_reg_60_3_inst : DFF_X1 port map( D => n8029, CK => CLK, Q => 
                           n_1862, QN => n4773);
   REGISTERS_reg_60_2_inst : DFF_X1 port map( D => n8028, CK => CLK, Q => 
                           n_1863, QN => n4772);
   REGISTERS_reg_60_1_inst : DFF_X1 port map( D => n8027, CK => CLK, Q => 
                           n_1864, QN => n4771);
   REGISTERS_reg_60_0_inst : DFF_X1 port map( D => n8026, CK => CLK, Q => 
                           n_1865, QN => n4770);
   REGISTERS_reg_61_31_inst : DFF_X1 port map( D => n8025, CK => CLK, Q => 
                           n_1866, QN => n4769);
   REGISTERS_reg_61_30_inst : DFF_X1 port map( D => n8024, CK => CLK, Q => 
                           n_1867, QN => n4768);
   REGISTERS_reg_61_29_inst : DFF_X1 port map( D => n8023, CK => CLK, Q => 
                           n_1868, QN => n4767);
   REGISTERS_reg_61_28_inst : DFF_X1 port map( D => n8022, CK => CLK, Q => 
                           n_1869, QN => n4766);
   REGISTERS_reg_61_27_inst : DFF_X1 port map( D => n8021, CK => CLK, Q => 
                           n_1870, QN => n4765);
   REGISTERS_reg_61_26_inst : DFF_X1 port map( D => n8020, CK => CLK, Q => 
                           n_1871, QN => n4764);
   REGISTERS_reg_61_25_inst : DFF_X1 port map( D => n8019, CK => CLK, Q => 
                           n_1872, QN => n4763);
   REGISTERS_reg_61_24_inst : DFF_X1 port map( D => n8018, CK => CLK, Q => 
                           n_1873, QN => n4762);
   REGISTERS_reg_61_23_inst : DFF_X1 port map( D => n8017, CK => CLK, Q => 
                           n_1874, QN => n4761);
   REGISTERS_reg_61_22_inst : DFF_X1 port map( D => n8016, CK => CLK, Q => 
                           n_1875, QN => n4760);
   REGISTERS_reg_61_21_inst : DFF_X1 port map( D => n8015, CK => CLK, Q => 
                           n_1876, QN => n4759);
   REGISTERS_reg_61_20_inst : DFF_X1 port map( D => n8014, CK => CLK, Q => 
                           n_1877, QN => n4758);
   REGISTERS_reg_61_19_inst : DFF_X1 port map( D => n8013, CK => CLK, Q => 
                           n_1878, QN => n4757);
   REGISTERS_reg_61_18_inst : DFF_X1 port map( D => n8012, CK => CLK, Q => 
                           n_1879, QN => n4756);
   REGISTERS_reg_61_17_inst : DFF_X1 port map( D => n8011, CK => CLK, Q => 
                           n_1880, QN => n4755);
   REGISTERS_reg_61_16_inst : DFF_X1 port map( D => n8010, CK => CLK, Q => 
                           n_1881, QN => n4754);
   REGISTERS_reg_61_15_inst : DFF_X1 port map( D => n8009, CK => CLK, Q => 
                           n_1882, QN => n4753);
   REGISTERS_reg_61_14_inst : DFF_X1 port map( D => n8008, CK => CLK, Q => 
                           n_1883, QN => n4752);
   REGISTERS_reg_61_13_inst : DFF_X1 port map( D => n8007, CK => CLK, Q => 
                           n_1884, QN => n4751);
   REGISTERS_reg_61_12_inst : DFF_X1 port map( D => n8006, CK => CLK, Q => 
                           n_1885, QN => n4750);
   REGISTERS_reg_61_11_inst : DFF_X1 port map( D => n8005, CK => CLK, Q => 
                           n_1886, QN => n4749);
   REGISTERS_reg_61_10_inst : DFF_X1 port map( D => n8004, CK => CLK, Q => 
                           n_1887, QN => n4748);
   REGISTERS_reg_61_9_inst : DFF_X1 port map( D => n8003, CK => CLK, Q => 
                           n_1888, QN => n4747);
   REGISTERS_reg_61_8_inst : DFF_X1 port map( D => n8002, CK => CLK, Q => 
                           n_1889, QN => n4746);
   REGISTERS_reg_61_7_inst : DFF_X1 port map( D => n8001, CK => CLK, Q => 
                           n_1890, QN => n4745);
   REGISTERS_reg_61_6_inst : DFF_X1 port map( D => n8000, CK => CLK, Q => 
                           n_1891, QN => n4744);
   REGISTERS_reg_61_5_inst : DFF_X1 port map( D => n7999, CK => CLK, Q => 
                           n_1892, QN => n4743);
   REGISTERS_reg_61_4_inst : DFF_X1 port map( D => n7998, CK => CLK, Q => 
                           n_1893, QN => n4742);
   REGISTERS_reg_61_3_inst : DFF_X1 port map( D => n7997, CK => CLK, Q => 
                           n_1894, QN => n4741);
   REGISTERS_reg_61_2_inst : DFF_X1 port map( D => n7996, CK => CLK, Q => 
                           n_1895, QN => n4740);
   REGISTERS_reg_61_1_inst : DFF_X1 port map( D => n7995, CK => CLK, Q => 
                           n_1896, QN => n4739);
   REGISTERS_reg_61_0_inst : DFF_X1 port map( D => n7994, CK => CLK, Q => 
                           n_1897, QN => n4738);
   REGISTERS_reg_62_31_inst : DFF_X1 port map( D => n7993, CK => CLK, Q => 
                           n_1898, QN => n4737);
   REGISTERS_reg_62_30_inst : DFF_X1 port map( D => n7992, CK => CLK, Q => 
                           n_1899, QN => n4736);
   REGISTERS_reg_62_29_inst : DFF_X1 port map( D => n7991, CK => CLK, Q => 
                           n_1900, QN => n4735);
   REGISTERS_reg_62_28_inst : DFF_X1 port map( D => n7990, CK => CLK, Q => 
                           n_1901, QN => n4734);
   REGISTERS_reg_62_27_inst : DFF_X1 port map( D => n7989, CK => CLK, Q => 
                           n_1902, QN => n4733);
   REGISTERS_reg_62_26_inst : DFF_X1 port map( D => n7988, CK => CLK, Q => 
                           n_1903, QN => n4732);
   REGISTERS_reg_62_25_inst : DFF_X1 port map( D => n7987, CK => CLK, Q => 
                           n_1904, QN => n4731);
   REGISTERS_reg_62_24_inst : DFF_X1 port map( D => n7986, CK => CLK, Q => 
                           n_1905, QN => n4730);
   REGISTERS_reg_62_23_inst : DFF_X1 port map( D => n7985, CK => CLK, Q => 
                           n_1906, QN => n4729);
   REGISTERS_reg_62_22_inst : DFF_X1 port map( D => n7984, CK => CLK, Q => 
                           n_1907, QN => n4728);
   REGISTERS_reg_62_21_inst : DFF_X1 port map( D => n7983, CK => CLK, Q => 
                           n_1908, QN => n4727);
   REGISTERS_reg_62_20_inst : DFF_X1 port map( D => n7982, CK => CLK, Q => 
                           n_1909, QN => n4726);
   REGISTERS_reg_62_19_inst : DFF_X1 port map( D => n7981, CK => CLK, Q => 
                           n_1910, QN => n4725);
   REGISTERS_reg_62_18_inst : DFF_X1 port map( D => n7980, CK => CLK, Q => 
                           n_1911, QN => n4724);
   REGISTERS_reg_62_17_inst : DFF_X1 port map( D => n7979, CK => CLK, Q => 
                           n_1912, QN => n4723);
   REGISTERS_reg_62_16_inst : DFF_X1 port map( D => n7978, CK => CLK, Q => 
                           n_1913, QN => n4722);
   REGISTERS_reg_62_15_inst : DFF_X1 port map( D => n7977, CK => CLK, Q => 
                           n_1914, QN => n4721);
   REGISTERS_reg_62_14_inst : DFF_X1 port map( D => n7976, CK => CLK, Q => 
                           n_1915, QN => n4720);
   REGISTERS_reg_62_13_inst : DFF_X1 port map( D => n7975, CK => CLK, Q => 
                           n_1916, QN => n4719);
   REGISTERS_reg_62_12_inst : DFF_X1 port map( D => n7974, CK => CLK, Q => 
                           n_1917, QN => n4718);
   REGISTERS_reg_62_11_inst : DFF_X1 port map( D => n7973, CK => CLK, Q => 
                           n_1918, QN => n4717);
   REGISTERS_reg_62_10_inst : DFF_X1 port map( D => n7972, CK => CLK, Q => 
                           n_1919, QN => n4716);
   REGISTERS_reg_62_9_inst : DFF_X1 port map( D => n7971, CK => CLK, Q => 
                           n_1920, QN => n4715);
   REGISTERS_reg_62_8_inst : DFF_X1 port map( D => n7970, CK => CLK, Q => 
                           n_1921, QN => n4714);
   REGISTERS_reg_62_7_inst : DFF_X1 port map( D => n7969, CK => CLK, Q => 
                           n_1922, QN => n4713);
   REGISTERS_reg_62_6_inst : DFF_X1 port map( D => n7968, CK => CLK, Q => 
                           n_1923, QN => n4712);
   REGISTERS_reg_62_5_inst : DFF_X1 port map( D => n7967, CK => CLK, Q => 
                           n_1924, QN => n4711);
   REGISTERS_reg_62_4_inst : DFF_X1 port map( D => n7966, CK => CLK, Q => 
                           n_1925, QN => n4710);
   REGISTERS_reg_62_3_inst : DFF_X1 port map( D => n7965, CK => CLK, Q => 
                           n_1926, QN => n4709);
   REGISTERS_reg_62_2_inst : DFF_X1 port map( D => n7964, CK => CLK, Q => 
                           n_1927, QN => n4708);
   REGISTERS_reg_62_1_inst : DFF_X1 port map( D => n7963, CK => CLK, Q => 
                           n_1928, QN => n4707);
   REGISTERS_reg_62_0_inst : DFF_X1 port map( D => n7962, CK => CLK, Q => 
                           n_1929, QN => n4706);
   REGISTERS_reg_63_31_inst : DFF_X1 port map( D => n7961, CK => CLK, Q => 
                           n5953, QN => n1033);
   REGISTERS_reg_63_30_inst : DFF_X1 port map( D => n7960, CK => CLK, Q => 
                           n5952, QN => n1034);
   REGISTERS_reg_63_29_inst : DFF_X1 port map( D => n7959, CK => CLK, Q => 
                           n5951, QN => n1035);
   REGISTERS_reg_63_28_inst : DFF_X1 port map( D => n7958, CK => CLK, Q => 
                           n5950, QN => n1036);
   REGISTERS_reg_63_27_inst : DFF_X1 port map( D => n7957, CK => CLK, Q => 
                           n5949, QN => n1037);
   REGISTERS_reg_63_26_inst : DFF_X1 port map( D => n7956, CK => CLK, Q => 
                           n5948, QN => n1038);
   REGISTERS_reg_63_25_inst : DFF_X1 port map( D => n7955, CK => CLK, Q => 
                           n5947, QN => n1039);
   REGISTERS_reg_63_24_inst : DFF_X1 port map( D => n7954, CK => CLK, Q => 
                           n5946, QN => n1040);
   REGISTERS_reg_63_23_inst : DFF_X1 port map( D => n7953, CK => CLK, Q => 
                           n5945, QN => n1041);
   REGISTERS_reg_63_22_inst : DFF_X1 port map( D => n7952, CK => CLK, Q => 
                           n5944, QN => n1042);
   REGISTERS_reg_63_21_inst : DFF_X1 port map( D => n7951, CK => CLK, Q => 
                           n5943, QN => n1043);
   REGISTERS_reg_63_20_inst : DFF_X1 port map( D => n7950, CK => CLK, Q => 
                           n5942, QN => n1044);
   REGISTERS_reg_63_19_inst : DFF_X1 port map( D => n7949, CK => CLK, Q => 
                           n5941, QN => n1045);
   REGISTERS_reg_63_18_inst : DFF_X1 port map( D => n7948, CK => CLK, Q => 
                           n5940, QN => n1046);
   REGISTERS_reg_63_17_inst : DFF_X1 port map( D => n7947, CK => CLK, Q => 
                           n5939, QN => n1047);
   REGISTERS_reg_63_16_inst : DFF_X1 port map( D => n7946, CK => CLK, Q => 
                           n5938, QN => n1048);
   REGISTERS_reg_63_15_inst : DFF_X1 port map( D => n7945, CK => CLK, Q => 
                           n5937, QN => n1049);
   REGISTERS_reg_63_14_inst : DFF_X1 port map( D => n7944, CK => CLK, Q => 
                           n5936, QN => n1050);
   REGISTERS_reg_63_13_inst : DFF_X1 port map( D => n7943, CK => CLK, Q => 
                           n5935, QN => n1051);
   REGISTERS_reg_63_12_inst : DFF_X1 port map( D => n7942, CK => CLK, Q => 
                           n5934, QN => n1052);
   REGISTERS_reg_63_11_inst : DFF_X1 port map( D => n7941, CK => CLK, Q => 
                           n5933, QN => n1053);
   REGISTERS_reg_63_10_inst : DFF_X1 port map( D => n7940, CK => CLK, Q => 
                           n5932, QN => n1054);
   REGISTERS_reg_63_9_inst : DFF_X1 port map( D => n7939, CK => CLK, Q => n5931
                           , QN => n1055);
   REGISTERS_reg_63_8_inst : DFF_X1 port map( D => n7938, CK => CLK, Q => n5930
                           , QN => n1056);
   REGISTERS_reg_63_7_inst : DFF_X1 port map( D => n7937, CK => CLK, Q => n5929
                           , QN => n1057);
   REGISTERS_reg_63_6_inst : DFF_X1 port map( D => n7936, CK => CLK, Q => n5928
                           , QN => n1058);
   REGISTERS_reg_63_5_inst : DFF_X1 port map( D => n7935, CK => CLK, Q => n5927
                           , QN => n1059);
   REGISTERS_reg_63_4_inst : DFF_X1 port map( D => n7934, CK => CLK, Q => n5926
                           , QN => n1060);
   REGISTERS_reg_63_3_inst : DFF_X1 port map( D => n7933, CK => CLK, Q => n5925
                           , QN => n1061);
   REGISTERS_reg_63_2_inst : DFF_X1 port map( D => n7932, CK => CLK, Q => n5924
                           , QN => n1062);
   REGISTERS_reg_63_1_inst : DFF_X1 port map( D => n7931, CK => CLK, Q => n5923
                           , QN => n1063);
   REGISTERS_reg_63_0_inst : DFF_X1 port map( D => n7930, CK => CLK, Q => n5922
                           , QN => n1064);
   REGISTERS_reg_64_31_inst : DFF_X1 port map( D => n7929, CK => CLK, Q => 
                           n5921, QN => n1385);
   REGISTERS_reg_64_30_inst : DFF_X1 port map( D => n7928, CK => CLK, Q => 
                           n5920, QN => n1386);
   REGISTERS_reg_64_29_inst : DFF_X1 port map( D => n7927, CK => CLK, Q => 
                           n5919, QN => n1387);
   REGISTERS_reg_64_28_inst : DFF_X1 port map( D => n7926, CK => CLK, Q => 
                           n5918, QN => n1388);
   REGISTERS_reg_64_27_inst : DFF_X1 port map( D => n7925, CK => CLK, Q => 
                           n5917, QN => n1389);
   REGISTERS_reg_64_26_inst : DFF_X1 port map( D => n7924, CK => CLK, Q => 
                           n5916, QN => n1390);
   REGISTERS_reg_64_25_inst : DFF_X1 port map( D => n7923, CK => CLK, Q => 
                           n5915, QN => n1391);
   REGISTERS_reg_64_24_inst : DFF_X1 port map( D => n7922, CK => CLK, Q => 
                           n5914, QN => n1392);
   REGISTERS_reg_64_23_inst : DFF_X1 port map( D => n7921, CK => CLK, Q => 
                           n5913, QN => n1393);
   REGISTERS_reg_64_22_inst : DFF_X1 port map( D => n7920, CK => CLK, Q => 
                           n5912, QN => n1394);
   REGISTERS_reg_64_21_inst : DFF_X1 port map( D => n7919, CK => CLK, Q => 
                           n5911, QN => n1395);
   REGISTERS_reg_64_20_inst : DFF_X1 port map( D => n7918, CK => CLK, Q => 
                           n5910, QN => n1396);
   REGISTERS_reg_64_19_inst : DFF_X1 port map( D => n7917, CK => CLK, Q => 
                           n5909, QN => n1397);
   REGISTERS_reg_64_18_inst : DFF_X1 port map( D => n7916, CK => CLK, Q => 
                           n5908, QN => n1398);
   REGISTERS_reg_64_17_inst : DFF_X1 port map( D => n7915, CK => CLK, Q => 
                           n5907, QN => n1399);
   REGISTERS_reg_64_16_inst : DFF_X1 port map( D => n7914, CK => CLK, Q => 
                           n5906, QN => n1400);
   REGISTERS_reg_64_15_inst : DFF_X1 port map( D => n7913, CK => CLK, Q => 
                           n5905, QN => n1401);
   REGISTERS_reg_64_14_inst : DFF_X1 port map( D => n7912, CK => CLK, Q => 
                           n5904, QN => n1402);
   REGISTERS_reg_64_13_inst : DFF_X1 port map( D => n7911, CK => CLK, Q => 
                           n5903, QN => n1403);
   REGISTERS_reg_64_12_inst : DFF_X1 port map( D => n7910, CK => CLK, Q => 
                           n5902, QN => n1404);
   REGISTERS_reg_64_11_inst : DFF_X1 port map( D => n7909, CK => CLK, Q => 
                           n5901, QN => n1405);
   REGISTERS_reg_64_10_inst : DFF_X1 port map( D => n7908, CK => CLK, Q => 
                           n5900, QN => n1406);
   REGISTERS_reg_64_9_inst : DFF_X1 port map( D => n7907, CK => CLK, Q => n5899
                           , QN => n1407);
   REGISTERS_reg_64_8_inst : DFF_X1 port map( D => n7906, CK => CLK, Q => n5898
                           , QN => n1408);
   REGISTERS_reg_64_7_inst : DFF_X1 port map( D => n7905, CK => CLK, Q => n5897
                           , QN => n1409);
   REGISTERS_reg_64_6_inst : DFF_X1 port map( D => n7904, CK => CLK, Q => n5896
                           , QN => n1410);
   REGISTERS_reg_64_5_inst : DFF_X1 port map( D => n7903, CK => CLK, Q => n5895
                           , QN => n1411);
   REGISTERS_reg_64_4_inst : DFF_X1 port map( D => n7902, CK => CLK, Q => n5894
                           , QN => n1412);
   REGISTERS_reg_64_3_inst : DFF_X1 port map( D => n7901, CK => CLK, Q => n5893
                           , QN => n1413);
   REGISTERS_reg_64_2_inst : DFF_X1 port map( D => n7900, CK => CLK, Q => n5892
                           , QN => n1414);
   REGISTERS_reg_64_1_inst : DFF_X1 port map( D => n7899, CK => CLK, Q => n5891
                           , QN => n1415);
   REGISTERS_reg_64_0_inst : DFF_X1 port map( D => n7898, CK => CLK, Q => n5890
                           , QN => n1416);
   REGISTERS_reg_65_31_inst : DFF_X1 port map( D => n7897, CK => CLK, Q => 
                           n_1930, QN => n4705);
   REGISTERS_reg_65_30_inst : DFF_X1 port map( D => n7896, CK => CLK, Q => 
                           n_1931, QN => n4704);
   REGISTERS_reg_65_29_inst : DFF_X1 port map( D => n7895, CK => CLK, Q => 
                           n_1932, QN => n4703);
   REGISTERS_reg_65_28_inst : DFF_X1 port map( D => n7894, CK => CLK, Q => 
                           n_1933, QN => n4702);
   REGISTERS_reg_65_27_inst : DFF_X1 port map( D => n7893, CK => CLK, Q => 
                           n_1934, QN => n4701);
   REGISTERS_reg_65_26_inst : DFF_X1 port map( D => n7892, CK => CLK, Q => 
                           n_1935, QN => n4700);
   REGISTERS_reg_65_25_inst : DFF_X1 port map( D => n7891, CK => CLK, Q => 
                           n_1936, QN => n4699);
   REGISTERS_reg_65_24_inst : DFF_X1 port map( D => n7890, CK => CLK, Q => 
                           n_1937, QN => n4698);
   REGISTERS_reg_65_23_inst : DFF_X1 port map( D => n7889, CK => CLK, Q => 
                           n_1938, QN => n4697);
   REGISTERS_reg_65_22_inst : DFF_X1 port map( D => n7888, CK => CLK, Q => 
                           n_1939, QN => n4696);
   REGISTERS_reg_65_21_inst : DFF_X1 port map( D => n7887, CK => CLK, Q => 
                           n_1940, QN => n4695);
   REGISTERS_reg_65_20_inst : DFF_X1 port map( D => n7886, CK => CLK, Q => 
                           n_1941, QN => n4694);
   REGISTERS_reg_65_19_inst : DFF_X1 port map( D => n7885, CK => CLK, Q => 
                           n_1942, QN => n4693);
   REGISTERS_reg_65_18_inst : DFF_X1 port map( D => n7884, CK => CLK, Q => 
                           n_1943, QN => n4692);
   REGISTERS_reg_65_17_inst : DFF_X1 port map( D => n7883, CK => CLK, Q => 
                           n_1944, QN => n4691);
   REGISTERS_reg_65_16_inst : DFF_X1 port map( D => n7882, CK => CLK, Q => 
                           n_1945, QN => n4690);
   REGISTERS_reg_65_15_inst : DFF_X1 port map( D => n7881, CK => CLK, Q => 
                           n_1946, QN => n4689);
   REGISTERS_reg_65_14_inst : DFF_X1 port map( D => n7880, CK => CLK, Q => 
                           n_1947, QN => n4688);
   REGISTERS_reg_65_13_inst : DFF_X1 port map( D => n7879, CK => CLK, Q => 
                           n_1948, QN => n4687);
   REGISTERS_reg_65_12_inst : DFF_X1 port map( D => n7878, CK => CLK, Q => 
                           n_1949, QN => n4686);
   REGISTERS_reg_65_11_inst : DFF_X1 port map( D => n7877, CK => CLK, Q => 
                           n_1950, QN => n4685);
   REGISTERS_reg_65_10_inst : DFF_X1 port map( D => n7876, CK => CLK, Q => 
                           n_1951, QN => n4684);
   REGISTERS_reg_65_9_inst : DFF_X1 port map( D => n7875, CK => CLK, Q => 
                           n_1952, QN => n4683);
   REGISTERS_reg_65_8_inst : DFF_X1 port map( D => n7874, CK => CLK, Q => 
                           n_1953, QN => n4682);
   REGISTERS_reg_65_7_inst : DFF_X1 port map( D => n7873, CK => CLK, Q => 
                           n_1954, QN => n4681);
   REGISTERS_reg_65_6_inst : DFF_X1 port map( D => n7872, CK => CLK, Q => 
                           n_1955, QN => n4680);
   REGISTERS_reg_65_5_inst : DFF_X1 port map( D => n7871, CK => CLK, Q => 
                           n_1956, QN => n4679);
   REGISTERS_reg_65_4_inst : DFF_X1 port map( D => n7870, CK => CLK, Q => 
                           n_1957, QN => n4678);
   REGISTERS_reg_65_3_inst : DFF_X1 port map( D => n7869, CK => CLK, Q => 
                           n_1958, QN => n4677);
   REGISTERS_reg_65_2_inst : DFF_X1 port map( D => n7868, CK => CLK, Q => 
                           n_1959, QN => n4676);
   REGISTERS_reg_65_1_inst : DFF_X1 port map( D => n7867, CK => CLK, Q => 
                           n_1960, QN => n4675);
   REGISTERS_reg_65_0_inst : DFF_X1 port map( D => n7866, CK => CLK, Q => 
                           n_1961, QN => n4674);
   REGISTERS_reg_66_31_inst : DFF_X1 port map( D => n7865, CK => CLK, Q => 
                           n_1962, QN => n4673);
   REGISTERS_reg_66_30_inst : DFF_X1 port map( D => n7864, CK => CLK, Q => 
                           n_1963, QN => n4672);
   REGISTERS_reg_66_29_inst : DFF_X1 port map( D => n7863, CK => CLK, Q => 
                           n_1964, QN => n4671);
   REGISTERS_reg_66_28_inst : DFF_X1 port map( D => n7862, CK => CLK, Q => 
                           n_1965, QN => n4670);
   REGISTERS_reg_66_27_inst : DFF_X1 port map( D => n7861, CK => CLK, Q => 
                           n_1966, QN => n4669);
   REGISTERS_reg_66_26_inst : DFF_X1 port map( D => n7860, CK => CLK, Q => 
                           n_1967, QN => n4668);
   REGISTERS_reg_66_25_inst : DFF_X1 port map( D => n7859, CK => CLK, Q => 
                           n_1968, QN => n4667);
   REGISTERS_reg_66_24_inst : DFF_X1 port map( D => n7858, CK => CLK, Q => 
                           n_1969, QN => n4666);
   REGISTERS_reg_66_23_inst : DFF_X1 port map( D => n7857, CK => CLK, Q => 
                           n_1970, QN => n4665);
   REGISTERS_reg_66_22_inst : DFF_X1 port map( D => n7856, CK => CLK, Q => 
                           n_1971, QN => n4664);
   REGISTERS_reg_66_21_inst : DFF_X1 port map( D => n7855, CK => CLK, Q => 
                           n_1972, QN => n4663);
   REGISTERS_reg_66_20_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => 
                           n_1973, QN => n4662);
   REGISTERS_reg_66_19_inst : DFF_X1 port map( D => n7853, CK => CLK, Q => 
                           n_1974, QN => n4661);
   REGISTERS_reg_66_18_inst : DFF_X1 port map( D => n7852, CK => CLK, Q => 
                           n_1975, QN => n4660);
   REGISTERS_reg_66_17_inst : DFF_X1 port map( D => n7851, CK => CLK, Q => 
                           n_1976, QN => n4659);
   REGISTERS_reg_66_16_inst : DFF_X1 port map( D => n7850, CK => CLK, Q => 
                           n_1977, QN => n4658);
   REGISTERS_reg_66_15_inst : DFF_X1 port map( D => n7849, CK => CLK, Q => 
                           n_1978, QN => n4657);
   REGISTERS_reg_66_14_inst : DFF_X1 port map( D => n7848, CK => CLK, Q => 
                           n_1979, QN => n4656);
   REGISTERS_reg_66_13_inst : DFF_X1 port map( D => n7847, CK => CLK, Q => 
                           n_1980, QN => n4655);
   REGISTERS_reg_66_12_inst : DFF_X1 port map( D => n7846, CK => CLK, Q => 
                           n_1981, QN => n4654);
   REGISTERS_reg_66_11_inst : DFF_X1 port map( D => n7845, CK => CLK, Q => 
                           n_1982, QN => n4653);
   REGISTERS_reg_66_10_inst : DFF_X1 port map( D => n7844, CK => CLK, Q => 
                           n_1983, QN => n4652);
   REGISTERS_reg_66_9_inst : DFF_X1 port map( D => n7843, CK => CLK, Q => 
                           n_1984, QN => n4651);
   REGISTERS_reg_66_8_inst : DFF_X1 port map( D => n7842, CK => CLK, Q => 
                           n_1985, QN => n4650);
   REGISTERS_reg_66_7_inst : DFF_X1 port map( D => n7841, CK => CLK, Q => 
                           n_1986, QN => n4649);
   REGISTERS_reg_66_6_inst : DFF_X1 port map( D => n7840, CK => CLK, Q => 
                           n_1987, QN => n4648);
   REGISTERS_reg_66_5_inst : DFF_X1 port map( D => n7839, CK => CLK, Q => 
                           n_1988, QN => n4647);
   REGISTERS_reg_66_4_inst : DFF_X1 port map( D => n7838, CK => CLK, Q => 
                           n_1989, QN => n4646);
   REGISTERS_reg_66_3_inst : DFF_X1 port map( D => n7837, CK => CLK, Q => 
                           n_1990, QN => n4645);
   REGISTERS_reg_66_2_inst : DFF_X1 port map( D => n7836, CK => CLK, Q => 
                           n_1991, QN => n4644);
   REGISTERS_reg_66_1_inst : DFF_X1 port map( D => n7835, CK => CLK, Q => 
                           n_1992, QN => n4643);
   REGISTERS_reg_66_0_inst : DFF_X1 port map( D => n7834, CK => CLK, Q => 
                           n_1993, QN => n4642);
   REGISTERS_reg_67_31_inst : DFF_X1 port map( D => n7833, CK => CLK, Q => 
                           n5889, QN => n1065);
   REGISTERS_reg_67_30_inst : DFF_X1 port map( D => n7832, CK => CLK, Q => 
                           n5888, QN => n1066);
   REGISTERS_reg_67_29_inst : DFF_X1 port map( D => n7831, CK => CLK, Q => 
                           n5887, QN => n1067);
   REGISTERS_reg_67_28_inst : DFF_X1 port map( D => n7830, CK => CLK, Q => 
                           n5886, QN => n1068);
   REGISTERS_reg_67_27_inst : DFF_X1 port map( D => n7829, CK => CLK, Q => 
                           n5885, QN => n1069);
   REGISTERS_reg_67_26_inst : DFF_X1 port map( D => n7828, CK => CLK, Q => 
                           n5884, QN => n1070);
   REGISTERS_reg_67_25_inst : DFF_X1 port map( D => n7827, CK => CLK, Q => 
                           n5883, QN => n1071);
   REGISTERS_reg_67_24_inst : DFF_X1 port map( D => n7826, CK => CLK, Q => 
                           n5882, QN => n1072);
   REGISTERS_reg_67_23_inst : DFF_X1 port map( D => n7825, CK => CLK, Q => 
                           n5881, QN => n1073);
   REGISTERS_reg_67_22_inst : DFF_X1 port map( D => n7824, CK => CLK, Q => 
                           n5880, QN => n1074);
   REGISTERS_reg_67_21_inst : DFF_X1 port map( D => n7823, CK => CLK, Q => 
                           n5879, QN => n1075);
   REGISTERS_reg_67_20_inst : DFF_X1 port map( D => n7822, CK => CLK, Q => 
                           n5878, QN => n1076);
   REGISTERS_reg_67_19_inst : DFF_X1 port map( D => n7821, CK => CLK, Q => 
                           n5877, QN => n1077);
   REGISTERS_reg_67_18_inst : DFF_X1 port map( D => n7820, CK => CLK, Q => 
                           n5876, QN => n1078);
   REGISTERS_reg_67_17_inst : DFF_X1 port map( D => n7819, CK => CLK, Q => 
                           n5875, QN => n1079);
   REGISTERS_reg_67_16_inst : DFF_X1 port map( D => n7818, CK => CLK, Q => 
                           n5874, QN => n1080);
   REGISTERS_reg_67_15_inst : DFF_X1 port map( D => n7817, CK => CLK, Q => 
                           n5873, QN => n1081);
   REGISTERS_reg_67_14_inst : DFF_X1 port map( D => n7816, CK => CLK, Q => 
                           n5872, QN => n1082);
   REGISTERS_reg_67_13_inst : DFF_X1 port map( D => n7815, CK => CLK, Q => 
                           n5871, QN => n1083);
   REGISTERS_reg_67_12_inst : DFF_X1 port map( D => n7814, CK => CLK, Q => 
                           n5870, QN => n1084);
   REGISTERS_reg_67_11_inst : DFF_X1 port map( D => n7813, CK => CLK, Q => 
                           n5869, QN => n1085);
   REGISTERS_reg_67_10_inst : DFF_X1 port map( D => n7812, CK => CLK, Q => 
                           n5868, QN => n1086);
   REGISTERS_reg_67_9_inst : DFF_X1 port map( D => n7811, CK => CLK, Q => n5867
                           , QN => n1087);
   REGISTERS_reg_67_8_inst : DFF_X1 port map( D => n7810, CK => CLK, Q => n5866
                           , QN => n1088);
   REGISTERS_reg_67_7_inst : DFF_X1 port map( D => n7809, CK => CLK, Q => n5865
                           , QN => n1089);
   REGISTERS_reg_67_6_inst : DFF_X1 port map( D => n7808, CK => CLK, Q => n5864
                           , QN => n1090);
   REGISTERS_reg_67_5_inst : DFF_X1 port map( D => n7807, CK => CLK, Q => n5863
                           , QN => n1091);
   REGISTERS_reg_67_4_inst : DFF_X1 port map( D => n7806, CK => CLK, Q => n5862
                           , QN => n1092);
   REGISTERS_reg_67_3_inst : DFF_X1 port map( D => n7805, CK => CLK, Q => n5861
                           , QN => n1093);
   REGISTERS_reg_67_2_inst : DFF_X1 port map( D => n7804, CK => CLK, Q => n5860
                           , QN => n1094);
   REGISTERS_reg_67_1_inst : DFF_X1 port map( D => n7803, CK => CLK, Q => n5859
                           , QN => n1095);
   REGISTERS_reg_67_0_inst : DFF_X1 port map( D => n7802, CK => CLK, Q => n5858
                           , QN => n1096);
   REGISTERS_reg_68_31_inst : DFF_X1 port map( D => n7801, CK => CLK, Q => 
                           n5857, QN => n1417);
   REGISTERS_reg_68_30_inst : DFF_X1 port map( D => n7800, CK => CLK, Q => 
                           n5856, QN => n1418);
   REGISTERS_reg_68_29_inst : DFF_X1 port map( D => n7799, CK => CLK, Q => 
                           n5855, QN => n1419);
   REGISTERS_reg_68_28_inst : DFF_X1 port map( D => n7798, CK => CLK, Q => 
                           n5854, QN => n1420);
   REGISTERS_reg_68_27_inst : DFF_X1 port map( D => n7797, CK => CLK, Q => 
                           n5853, QN => n1421);
   REGISTERS_reg_68_26_inst : DFF_X1 port map( D => n7796, CK => CLK, Q => 
                           n5852, QN => n1422);
   REGISTERS_reg_68_25_inst : DFF_X1 port map( D => n7795, CK => CLK, Q => 
                           n5851, QN => n1423);
   REGISTERS_reg_68_24_inst : DFF_X1 port map( D => n7794, CK => CLK, Q => 
                           n5850, QN => n1424);
   REGISTERS_reg_68_23_inst : DFF_X1 port map( D => n7793, CK => CLK, Q => 
                           n5849, QN => n1425);
   REGISTERS_reg_68_22_inst : DFF_X1 port map( D => n7792, CK => CLK, Q => 
                           n5848, QN => n1426);
   REGISTERS_reg_68_21_inst : DFF_X1 port map( D => n7791, CK => CLK, Q => 
                           n5847, QN => n1427);
   REGISTERS_reg_68_20_inst : DFF_X1 port map( D => n7790, CK => CLK, Q => 
                           n5846, QN => n1428);
   REGISTERS_reg_68_19_inst : DFF_X1 port map( D => n7789, CK => CLK, Q => 
                           n5845, QN => n1429);
   REGISTERS_reg_68_18_inst : DFF_X1 port map( D => n7788, CK => CLK, Q => 
                           n5844, QN => n1430);
   REGISTERS_reg_68_17_inst : DFF_X1 port map( D => n7787, CK => CLK, Q => 
                           n5843, QN => n1431);
   REGISTERS_reg_68_16_inst : DFF_X1 port map( D => n7786, CK => CLK, Q => 
                           n5842, QN => n1432);
   REGISTERS_reg_68_15_inst : DFF_X1 port map( D => n7785, CK => CLK, Q => 
                           n5841, QN => n1433);
   REGISTERS_reg_68_14_inst : DFF_X1 port map( D => n7784, CK => CLK, Q => 
                           n5840, QN => n1434);
   REGISTERS_reg_68_13_inst : DFF_X1 port map( D => n7783, CK => CLK, Q => 
                           n5839, QN => n1435);
   REGISTERS_reg_68_12_inst : DFF_X1 port map( D => n7782, CK => CLK, Q => 
                           n5838, QN => n1436);
   REGISTERS_reg_68_11_inst : DFF_X1 port map( D => n7781, CK => CLK, Q => 
                           n5837, QN => n1437);
   REGISTERS_reg_68_10_inst : DFF_X1 port map( D => n7780, CK => CLK, Q => 
                           n5836, QN => n1438);
   REGISTERS_reg_68_9_inst : DFF_X1 port map( D => n7779, CK => CLK, Q => n5835
                           , QN => n1439);
   REGISTERS_reg_68_8_inst : DFF_X1 port map( D => n7778, CK => CLK, Q => n5834
                           , QN => n1440);
   REGISTERS_reg_68_7_inst : DFF_X1 port map( D => n7777, CK => CLK, Q => n5833
                           , QN => n1441);
   REGISTERS_reg_68_6_inst : DFF_X1 port map( D => n7776, CK => CLK, Q => n5832
                           , QN => n1442);
   REGISTERS_reg_68_5_inst : DFF_X1 port map( D => n7775, CK => CLK, Q => n5831
                           , QN => n1443);
   REGISTERS_reg_68_4_inst : DFF_X1 port map( D => n7774, CK => CLK, Q => n5830
                           , QN => n1444);
   REGISTERS_reg_68_3_inst : DFF_X1 port map( D => n7773, CK => CLK, Q => n5829
                           , QN => n1445);
   REGISTERS_reg_68_2_inst : DFF_X1 port map( D => n7772, CK => CLK, Q => n5828
                           , QN => n1446);
   REGISTERS_reg_68_1_inst : DFF_X1 port map( D => n7771, CK => CLK, Q => n5827
                           , QN => n1447);
   REGISTERS_reg_68_0_inst : DFF_X1 port map( D => n7770, CK => CLK, Q => n5826
                           , QN => n1448);
   REGISTERS_reg_69_31_inst : DFF_X1 port map( D => n7769, CK => CLK, Q => 
                           n_1994, QN => n4641);
   REGISTERS_reg_69_30_inst : DFF_X1 port map( D => n7768, CK => CLK, Q => 
                           n_1995, QN => n4640);
   REGISTERS_reg_69_29_inst : DFF_X1 port map( D => n7767, CK => CLK, Q => 
                           n_1996, QN => n4639);
   REGISTERS_reg_69_28_inst : DFF_X1 port map( D => n7766, CK => CLK, Q => 
                           n_1997, QN => n4638);
   REGISTERS_reg_69_27_inst : DFF_X1 port map( D => n7765, CK => CLK, Q => 
                           n_1998, QN => n4637);
   REGISTERS_reg_69_26_inst : DFF_X1 port map( D => n7764, CK => CLK, Q => 
                           n_1999, QN => n4636);
   REGISTERS_reg_69_25_inst : DFF_X1 port map( D => n7763, CK => CLK, Q => 
                           n_2000, QN => n4635);
   REGISTERS_reg_69_24_inst : DFF_X1 port map( D => n7762, CK => CLK, Q => 
                           n_2001, QN => n4634);
   REGISTERS_reg_69_23_inst : DFF_X1 port map( D => n7761, CK => CLK, Q => 
                           n_2002, QN => n4633);
   REGISTERS_reg_69_22_inst : DFF_X1 port map( D => n7760, CK => CLK, Q => 
                           n_2003, QN => n4632);
   REGISTERS_reg_69_21_inst : DFF_X1 port map( D => n7759, CK => CLK, Q => 
                           n_2004, QN => n4631);
   REGISTERS_reg_69_20_inst : DFF_X1 port map( D => n7758, CK => CLK, Q => 
                           n_2005, QN => n4630);
   REGISTERS_reg_69_19_inst : DFF_X1 port map( D => n7757, CK => CLK, Q => 
                           n_2006, QN => n4629);
   REGISTERS_reg_69_18_inst : DFF_X1 port map( D => n7756, CK => CLK, Q => 
                           n_2007, QN => n4628);
   REGISTERS_reg_69_17_inst : DFF_X1 port map( D => n7755, CK => CLK, Q => 
                           n_2008, QN => n4627);
   REGISTERS_reg_69_16_inst : DFF_X1 port map( D => n7754, CK => CLK, Q => 
                           n_2009, QN => n4626);
   REGISTERS_reg_69_15_inst : DFF_X1 port map( D => n7753, CK => CLK, Q => 
                           n_2010, QN => n4625);
   REGISTERS_reg_69_14_inst : DFF_X1 port map( D => n7752, CK => CLK, Q => 
                           n_2011, QN => n4624);
   REGISTERS_reg_69_13_inst : DFF_X1 port map( D => n7751, CK => CLK, Q => 
                           n_2012, QN => n4623);
   REGISTERS_reg_69_12_inst : DFF_X1 port map( D => n7750, CK => CLK, Q => 
                           n_2013, QN => n4622);
   REGISTERS_reg_69_11_inst : DFF_X1 port map( D => n7749, CK => CLK, Q => 
                           n_2014, QN => n4621);
   REGISTERS_reg_69_10_inst : DFF_X1 port map( D => n7748, CK => CLK, Q => 
                           n_2015, QN => n4620);
   REGISTERS_reg_69_9_inst : DFF_X1 port map( D => n7747, CK => CLK, Q => 
                           n_2016, QN => n4619);
   REGISTERS_reg_69_8_inst : DFF_X1 port map( D => n7746, CK => CLK, Q => 
                           n_2017, QN => n4618);
   REGISTERS_reg_69_7_inst : DFF_X1 port map( D => n7745, CK => CLK, Q => 
                           n_2018, QN => n4617);
   REGISTERS_reg_69_6_inst : DFF_X1 port map( D => n7744, CK => CLK, Q => 
                           n_2019, QN => n4616);
   REGISTERS_reg_69_5_inst : DFF_X1 port map( D => n7743, CK => CLK, Q => 
                           n_2020, QN => n4615);
   REGISTERS_reg_69_4_inst : DFF_X1 port map( D => n7742, CK => CLK, Q => 
                           n_2021, QN => n4614);
   REGISTERS_reg_69_3_inst : DFF_X1 port map( D => n7741, CK => CLK, Q => 
                           n_2022, QN => n4613);
   REGISTERS_reg_69_2_inst : DFF_X1 port map( D => n7740, CK => CLK, Q => 
                           n_2023, QN => n4612);
   REGISTERS_reg_69_1_inst : DFF_X1 port map( D => n7739, CK => CLK, Q => 
                           n_2024, QN => n4611);
   REGISTERS_reg_69_0_inst : DFF_X1 port map( D => n7738, CK => CLK, Q => 
                           n_2025, QN => n4610);
   REGISTERS_reg_70_31_inst : DFF_X1 port map( D => n7737, CK => CLK, Q => 
                           n_2026, QN => n4609);
   REGISTERS_reg_70_30_inst : DFF_X1 port map( D => n7736, CK => CLK, Q => 
                           n_2027, QN => n4608);
   REGISTERS_reg_70_29_inst : DFF_X1 port map( D => n7735, CK => CLK, Q => 
                           n_2028, QN => n4607);
   REGISTERS_reg_70_28_inst : DFF_X1 port map( D => n7734, CK => CLK, Q => 
                           n_2029, QN => n4606);
   REGISTERS_reg_70_27_inst : DFF_X1 port map( D => n7733, CK => CLK, Q => 
                           n_2030, QN => n4605);
   REGISTERS_reg_70_26_inst : DFF_X1 port map( D => n7732, CK => CLK, Q => 
                           n_2031, QN => n4604);
   REGISTERS_reg_70_25_inst : DFF_X1 port map( D => n7731, CK => CLK, Q => 
                           n_2032, QN => n4603);
   REGISTERS_reg_70_24_inst : DFF_X1 port map( D => n7730, CK => CLK, Q => 
                           n_2033, QN => n4602);
   REGISTERS_reg_70_23_inst : DFF_X1 port map( D => n7729, CK => CLK, Q => 
                           n_2034, QN => n4601);
   REGISTERS_reg_70_22_inst : DFF_X1 port map( D => n7728, CK => CLK, Q => 
                           n_2035, QN => n4600);
   REGISTERS_reg_70_21_inst : DFF_X1 port map( D => n7727, CK => CLK, Q => 
                           n_2036, QN => n4599);
   REGISTERS_reg_70_20_inst : DFF_X1 port map( D => n7726, CK => CLK, Q => 
                           n_2037, QN => n4598);
   REGISTERS_reg_70_19_inst : DFF_X1 port map( D => n7725, CK => CLK, Q => 
                           n_2038, QN => n4597);
   REGISTERS_reg_70_18_inst : DFF_X1 port map( D => n7724, CK => CLK, Q => 
                           n_2039, QN => n4596);
   REGISTERS_reg_70_17_inst : DFF_X1 port map( D => n7723, CK => CLK, Q => 
                           n_2040, QN => n4595);
   REGISTERS_reg_70_16_inst : DFF_X1 port map( D => n7722, CK => CLK, Q => 
                           n_2041, QN => n4594);
   REGISTERS_reg_70_15_inst : DFF_X1 port map( D => n7721, CK => CLK, Q => 
                           n_2042, QN => n4593);
   REGISTERS_reg_70_14_inst : DFF_X1 port map( D => n7720, CK => CLK, Q => 
                           n_2043, QN => n4592);
   REGISTERS_reg_70_13_inst : DFF_X1 port map( D => n7719, CK => CLK, Q => 
                           n_2044, QN => n4591);
   REGISTERS_reg_70_12_inst : DFF_X1 port map( D => n7718, CK => CLK, Q => 
                           n_2045, QN => n4590);
   REGISTERS_reg_70_11_inst : DFF_X1 port map( D => n7717, CK => CLK, Q => 
                           n_2046, QN => n4589);
   REGISTERS_reg_70_10_inst : DFF_X1 port map( D => n7716, CK => CLK, Q => 
                           n_2047, QN => n4588);
   REGISTERS_reg_70_9_inst : DFF_X1 port map( D => n7715, CK => CLK, Q => 
                           n_2048, QN => n4587);
   REGISTERS_reg_70_8_inst : DFF_X1 port map( D => n7714, CK => CLK, Q => 
                           n_2049, QN => n4586);
   REGISTERS_reg_70_7_inst : DFF_X1 port map( D => n7713, CK => CLK, Q => 
                           n_2050, QN => n4585);
   REGISTERS_reg_70_6_inst : DFF_X1 port map( D => n7712, CK => CLK, Q => 
                           n_2051, QN => n4584);
   REGISTERS_reg_70_5_inst : DFF_X1 port map( D => n7711, CK => CLK, Q => 
                           n_2052, QN => n4583);
   REGISTERS_reg_70_4_inst : DFF_X1 port map( D => n7710, CK => CLK, Q => 
                           n_2053, QN => n4582);
   REGISTERS_reg_70_3_inst : DFF_X1 port map( D => n7709, CK => CLK, Q => 
                           n_2054, QN => n4581);
   REGISTERS_reg_70_2_inst : DFF_X1 port map( D => n7708, CK => CLK, Q => 
                           n_2055, QN => n4580);
   REGISTERS_reg_70_1_inst : DFF_X1 port map( D => n7707, CK => CLK, Q => 
                           n_2056, QN => n4579);
   REGISTERS_reg_70_0_inst : DFF_X1 port map( D => n7706, CK => CLK, Q => 
                           n_2057, QN => n4578);
   REGISTERS_reg_71_31_inst : DFF_X1 port map( D => n7705, CK => CLK, Q => 
                           n_2058, QN => n4577);
   REGISTERS_reg_71_30_inst : DFF_X1 port map( D => n7704, CK => CLK, Q => 
                           n_2059, QN => n4576);
   REGISTERS_reg_71_29_inst : DFF_X1 port map( D => n7703, CK => CLK, Q => 
                           n_2060, QN => n4575);
   REGISTERS_reg_71_28_inst : DFF_X1 port map( D => n7702, CK => CLK, Q => 
                           n_2061, QN => n4574);
   REGISTERS_reg_71_27_inst : DFF_X1 port map( D => n7701, CK => CLK, Q => 
                           n_2062, QN => n4573);
   REGISTERS_reg_71_26_inst : DFF_X1 port map( D => n7700, CK => CLK, Q => 
                           n_2063, QN => n4572);
   REGISTERS_reg_71_25_inst : DFF_X1 port map( D => n7699, CK => CLK, Q => 
                           n_2064, QN => n4571);
   REGISTERS_reg_71_24_inst : DFF_X1 port map( D => n7698, CK => CLK, Q => 
                           n_2065, QN => n4570);
   REGISTERS_reg_71_23_inst : DFF_X1 port map( D => n7697, CK => CLK, Q => 
                           n_2066, QN => n4569);
   REGISTERS_reg_71_22_inst : DFF_X1 port map( D => n7696, CK => CLK, Q => 
                           n_2067, QN => n4568);
   REGISTERS_reg_71_21_inst : DFF_X1 port map( D => n7695, CK => CLK, Q => 
                           n_2068, QN => n4567);
   REGISTERS_reg_71_20_inst : DFF_X1 port map( D => n7694, CK => CLK, Q => 
                           n_2069, QN => n4566);
   REGISTERS_reg_71_19_inst : DFF_X1 port map( D => n7693, CK => CLK, Q => 
                           n_2070, QN => n4565);
   REGISTERS_reg_71_18_inst : DFF_X1 port map( D => n7692, CK => CLK, Q => 
                           n_2071, QN => n4564);
   REGISTERS_reg_71_17_inst : DFF_X1 port map( D => n7691, CK => CLK, Q => 
                           n_2072, QN => n4563);
   REGISTERS_reg_71_16_inst : DFF_X1 port map( D => n7690, CK => CLK, Q => 
                           n_2073, QN => n4562);
   REGISTERS_reg_71_15_inst : DFF_X1 port map( D => n7689, CK => CLK, Q => 
                           n_2074, QN => n4561);
   REGISTERS_reg_71_14_inst : DFF_X1 port map( D => n7688, CK => CLK, Q => 
                           n_2075, QN => n4560);
   REGISTERS_reg_71_13_inst : DFF_X1 port map( D => n7687, CK => CLK, Q => 
                           n_2076, QN => n4559);
   REGISTERS_reg_71_12_inst : DFF_X1 port map( D => n7686, CK => CLK, Q => 
                           n_2077, QN => n4558);
   REGISTERS_reg_71_11_inst : DFF_X1 port map( D => n7685, CK => CLK, Q => 
                           n_2078, QN => n4557);
   REGISTERS_reg_71_10_inst : DFF_X1 port map( D => n7684, CK => CLK, Q => 
                           n_2079, QN => n4556);
   REGISTERS_reg_71_9_inst : DFF_X1 port map( D => n7683, CK => CLK, Q => 
                           n_2080, QN => n4555);
   REGISTERS_reg_71_8_inst : DFF_X1 port map( D => n7682, CK => CLK, Q => 
                           n_2081, QN => n4554);
   REGISTERS_reg_71_7_inst : DFF_X1 port map( D => n7681, CK => CLK, Q => 
                           n_2082, QN => n4553);
   REGISTERS_reg_71_6_inst : DFF_X1 port map( D => n7680, CK => CLK, Q => 
                           n_2083, QN => n4552);
   REGISTERS_reg_71_5_inst : DFF_X1 port map( D => n7679, CK => CLK, Q => 
                           n_2084, QN => n4551);
   REGISTERS_reg_71_4_inst : DFF_X1 port map( D => n7678, CK => CLK, Q => 
                           n_2085, QN => n4550);
   REGISTERS_reg_71_3_inst : DFF_X1 port map( D => n7677, CK => CLK, Q => 
                           n_2086, QN => n4549);
   REGISTERS_reg_71_2_inst : DFF_X1 port map( D => n7676, CK => CLK, Q => 
                           n_2087, QN => n4548);
   REGISTERS_reg_71_1_inst : DFF_X1 port map( D => n7675, CK => CLK, Q => 
                           n_2088, QN => n4547);
   REGISTERS_reg_71_0_inst : DFF_X1 port map( D => n7674, CK => CLK, Q => 
                           n_2089, QN => n4546);
   OUT1_reg_31_inst : DFF_X1 port map( D => n7673, CK => CLK, Q => n6658, QN =>
                           n1449);
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n7672, CK => CLK, Q => 
                           n6659, QN => n1513);
   OUT1_reg_30_inst : DFF_X1 port map( D => n7671, CK => CLK, Q => n6660, QN =>
                           n1450);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n7670, CK => CLK, Q => 
                           n6661, QN => n1514);
   OUT1_reg_29_inst : DFF_X1 port map( D => n7669, CK => CLK, Q => n6662, QN =>
                           n1451);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n7668, CK => CLK, Q => 
                           n6663, QN => n1515);
   OUT1_reg_28_inst : DFF_X1 port map( D => n7667, CK => CLK, Q => n6664, QN =>
                           n1452);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n7666, CK => CLK, Q => 
                           n6665, QN => n1516);
   OUT1_reg_27_inst : DFF_X1 port map( D => n7665, CK => CLK, Q => n6666, QN =>
                           n1453);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n7664, CK => CLK, Q => 
                           n6667, QN => n1517);
   OUT1_reg_26_inst : DFF_X1 port map( D => n7663, CK => CLK, Q => n6668, QN =>
                           n1454);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n7662, CK => CLK, Q => 
                           n6669, QN => n1518);
   OUT1_reg_25_inst : DFF_X1 port map( D => n7661, CK => CLK, Q => n6670, QN =>
                           n1455);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n7660, CK => CLK, Q => 
                           n6671, QN => n1519);
   OUT1_reg_24_inst : DFF_X1 port map( D => n7659, CK => CLK, Q => n6672, QN =>
                           n1456);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n7658, CK => CLK, Q => 
                           n6673, QN => n1520);
   OUT1_reg_23_inst : DFF_X1 port map( D => n7657, CK => CLK, Q => n6674, QN =>
                           n1457);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n7656, CK => CLK, Q => 
                           n6675, QN => n1521);
   OUT1_reg_22_inst : DFF_X1 port map( D => n7655, CK => CLK, Q => n6676, QN =>
                           n1458);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n7654, CK => CLK, Q => 
                           n6677, QN => n1522);
   OUT1_reg_21_inst : DFF_X1 port map( D => n7653, CK => CLK, Q => n6678, QN =>
                           n1459);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n7652, CK => CLK, Q => 
                           n6679, QN => n1523);
   OUT1_reg_20_inst : DFF_X1 port map( D => n7651, CK => CLK, Q => n6680, QN =>
                           n1460);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n7650, CK => CLK, Q => 
                           n6681, QN => n1524);
   OUT1_reg_19_inst : DFF_X1 port map( D => n7649, CK => CLK, Q => n6682, QN =>
                           n1461);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n7648, CK => CLK, Q => 
                           n6683, QN => n1525);
   OUT1_reg_18_inst : DFF_X1 port map( D => n7647, CK => CLK, Q => n6684, QN =>
                           n1462);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n7646, CK => CLK, Q => 
                           n6685, QN => n1526);
   OUT1_reg_17_inst : DFF_X1 port map( D => n7645, CK => CLK, Q => n6686, QN =>
                           n1463);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n7644, CK => CLK, Q => 
                           n6687, QN => n1527);
   OUT1_reg_16_inst : DFF_X1 port map( D => n7643, CK => CLK, Q => n6688, QN =>
                           n1464);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n7642, CK => CLK, Q => 
                           n6689, QN => n1528);
   OUT1_reg_15_inst : DFF_X1 port map( D => n7641, CK => CLK, Q => n6690, QN =>
                           n1465);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n7640, CK => CLK, Q => 
                           n6691, QN => n1529);
   OUT1_reg_14_inst : DFF_X1 port map( D => n7639, CK => CLK, Q => n6692, QN =>
                           n1466);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n7638, CK => CLK, Q => 
                           n6693, QN => n1530);
   OUT1_reg_13_inst : DFF_X1 port map( D => n7637, CK => CLK, Q => n6694, QN =>
                           n1467);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n7636, CK => CLK, Q => 
                           n6695, QN => n1531);
   OUT1_reg_12_inst : DFF_X1 port map( D => n7635, CK => CLK, Q => n6696, QN =>
                           n1468);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n7634, CK => CLK, Q => 
                           n6697, QN => n1532);
   OUT1_reg_11_inst : DFF_X1 port map( D => n7633, CK => CLK, Q => n6698, QN =>
                           n1469);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n7632, CK => CLK, Q => 
                           n6699, QN => n1533);
   OUT1_reg_10_inst : DFF_X1 port map( D => n7631, CK => CLK, Q => n6700, QN =>
                           n1470);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n7630, CK => CLK, Q => 
                           n6701, QN => n1534);
   OUT1_reg_9_inst : DFF_X1 port map( D => n7629, CK => CLK, Q => n6702, QN => 
                           n1471);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n7628, CK => CLK, Q => 
                           n6703, QN => n1535);
   OUT1_reg_8_inst : DFF_X1 port map( D => n7627, CK => CLK, Q => n6704, QN => 
                           n1472);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n7626, CK => CLK, Q => 
                           n6705, QN => n1536);
   OUT1_reg_7_inst : DFF_X1 port map( D => n7625, CK => CLK, Q => n6706, QN => 
                           n1473);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n7624, CK => CLK, Q => 
                           n6707, QN => n1537);
   OUT1_reg_6_inst : DFF_X1 port map( D => n7623, CK => CLK, Q => n6708, QN => 
                           n1474);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n7622, CK => CLK, Q => 
                           n6709, QN => n1538);
   OUT1_reg_5_inst : DFF_X1 port map( D => n7621, CK => CLK, Q => n6710, QN => 
                           n1475);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n7620, CK => CLK, Q => 
                           n6711, QN => n1539);
   OUT1_reg_4_inst : DFF_X1 port map( D => n7619, CK => CLK, Q => n6712, QN => 
                           n1476);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n7618, CK => CLK, Q => 
                           n6713, QN => n1540);
   OUT1_reg_3_inst : DFF_X1 port map( D => n7617, CK => CLK, Q => n6714, QN => 
                           n1477);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n7616, CK => CLK, Q => 
                           n6715, QN => n1541);
   OUT1_reg_2_inst : DFF_X1 port map( D => n7615, CK => CLK, Q => n6716, QN => 
                           n1478);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n7614, CK => CLK, Q => 
                           n6717, QN => n1542);
   OUT1_reg_1_inst : DFF_X1 port map( D => n7613, CK => CLK, Q => n6718, QN => 
                           n1479);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n7612, CK => CLK, Q => 
                           n6719, QN => n1543);
   OUT1_reg_0_inst : DFF_X1 port map( D => n7611, CK => CLK, Q => n6720, QN => 
                           n1480);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n7610, CK => CLK, Q => 
                           n6721, QN => n1544);
   OUT2_reg_31_inst : DFF_X1 port map( D => n7609, CK => CLK, Q => n6722, QN =>
                           n1481);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n7608, CK => CLK, Q => 
                           n6723, QN => n1545);
   OUT2_reg_30_inst : DFF_X1 port map( D => n7607, CK => CLK, Q => n6724, QN =>
                           n1482);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n7606, CK => CLK, Q => 
                           n6725, QN => n1546);
   OUT2_reg_29_inst : DFF_X1 port map( D => n7605, CK => CLK, Q => n6726, QN =>
                           n1483);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n7604, CK => CLK, Q => 
                           n6727, QN => n1547);
   OUT2_reg_28_inst : DFF_X1 port map( D => n7603, CK => CLK, Q => n6728, QN =>
                           n1484);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n7602, CK => CLK, Q => 
                           n6729, QN => n1548);
   OUT2_reg_27_inst : DFF_X1 port map( D => n7601, CK => CLK, Q => n6730, QN =>
                           n1485);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n7600, CK => CLK, Q => 
                           n6731, QN => n1549);
   OUT2_reg_26_inst : DFF_X1 port map( D => n7599, CK => CLK, Q => n6732, QN =>
                           n1486);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n7598, CK => CLK, Q => 
                           n6733, QN => n1550);
   OUT2_reg_25_inst : DFF_X1 port map( D => n7597, CK => CLK, Q => n6734, QN =>
                           n1487);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n7596, CK => CLK, Q => 
                           n6735, QN => n1551);
   OUT2_reg_24_inst : DFF_X1 port map( D => n7595, CK => CLK, Q => n6736, QN =>
                           n1488);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n7594, CK => CLK, Q => 
                           n6737, QN => n1552);
   OUT2_reg_23_inst : DFF_X1 port map( D => n7593, CK => CLK, Q => n6738, QN =>
                           n1489);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n7592, CK => CLK, Q => 
                           n6739, QN => n1553);
   OUT2_reg_22_inst : DFF_X1 port map( D => n7591, CK => CLK, Q => n6740, QN =>
                           n1490);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n7590, CK => CLK, Q => 
                           n6741, QN => n1554);
   OUT2_reg_21_inst : DFF_X1 port map( D => n7589, CK => CLK, Q => n6742, QN =>
                           n1491);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n7588, CK => CLK, Q => 
                           n6743, QN => n1555);
   OUT2_reg_20_inst : DFF_X1 port map( D => n7587, CK => CLK, Q => n6744, QN =>
                           n1492);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n7586, CK => CLK, Q => 
                           n6745, QN => n1556);
   OUT2_reg_19_inst : DFF_X1 port map( D => n7585, CK => CLK, Q => n6746, QN =>
                           n1493);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n7584, CK => CLK, Q => 
                           n6747, QN => n1557);
   OUT2_reg_18_inst : DFF_X1 port map( D => n7583, CK => CLK, Q => n6748, QN =>
                           n1494);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n7582, CK => CLK, Q => 
                           n6749, QN => n1558);
   OUT2_reg_17_inst : DFF_X1 port map( D => n7581, CK => CLK, Q => n6750, QN =>
                           n1495);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n7580, CK => CLK, Q => 
                           n6751, QN => n1559);
   OUT2_reg_16_inst : DFF_X1 port map( D => n7579, CK => CLK, Q => n6752, QN =>
                           n1496);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n7578, CK => CLK, Q => 
                           n6753, QN => n1560);
   OUT2_reg_15_inst : DFF_X1 port map( D => n7577, CK => CLK, Q => n6754, QN =>
                           n1497);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n7576, CK => CLK, Q => 
                           n6755, QN => n1561);
   OUT2_reg_14_inst : DFF_X1 port map( D => n7575, CK => CLK, Q => n6756, QN =>
                           n1498);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n7574, CK => CLK, Q => 
                           n6757, QN => n1562);
   OUT2_reg_13_inst : DFF_X1 port map( D => n7573, CK => CLK, Q => n6758, QN =>
                           n1499);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n7572, CK => CLK, Q => 
                           n6759, QN => n1563);
   OUT2_reg_12_inst : DFF_X1 port map( D => n7571, CK => CLK, Q => n6760, QN =>
                           n1500);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n7570, CK => CLK, Q => 
                           n6761, QN => n1564);
   OUT2_reg_11_inst : DFF_X1 port map( D => n7569, CK => CLK, Q => n6762, QN =>
                           n1501);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n7568, CK => CLK, Q => 
                           n6763, QN => n1565);
   OUT2_reg_10_inst : DFF_X1 port map( D => n7567, CK => CLK, Q => n6764, QN =>
                           n1502);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n7566, CK => CLK, Q => 
                           n6765, QN => n1566);
   OUT2_reg_9_inst : DFF_X1 port map( D => n7565, CK => CLK, Q => n6766, QN => 
                           n1503);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n7564, CK => CLK, Q => 
                           n6767, QN => n1567);
   OUT2_reg_8_inst : DFF_X1 port map( D => n7563, CK => CLK, Q => n6768, QN => 
                           n1504);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n7562, CK => CLK, Q => 
                           n6769, QN => n1568);
   OUT2_reg_7_inst : DFF_X1 port map( D => n7561, CK => CLK, Q => n6770, QN => 
                           n1505);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n7560, CK => CLK, Q => 
                           n6771, QN => n1569);
   OUT2_reg_6_inst : DFF_X1 port map( D => n7559, CK => CLK, Q => n6772, QN => 
                           n1506);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n7558, CK => CLK, Q => 
                           n6773, QN => n1570);
   OUT2_reg_5_inst : DFF_X1 port map( D => n7557, CK => CLK, Q => n6774, QN => 
                           n1507);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n7556, CK => CLK, Q => 
                           n6775, QN => n1571);
   OUT2_reg_4_inst : DFF_X1 port map( D => n7555, CK => CLK, Q => n6776, QN => 
                           n1508);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n7554, CK => CLK, Q => 
                           n6777, QN => n1572);
   OUT2_reg_3_inst : DFF_X1 port map( D => n7553, CK => CLK, Q => n6778, QN => 
                           n1509);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n7552, CK => CLK, Q => 
                           n6779, QN => n1573);
   OUT2_reg_2_inst : DFF_X1 port map( D => n7551, CK => CLK, Q => n6780, QN => 
                           n1510);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n7550, CK => CLK, Q => 
                           n6781, QN => n1574);
   OUT2_reg_1_inst : DFF_X1 port map( D => n7549, CK => CLK, Q => n6782, QN => 
                           n1511);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n7548, CK => CLK, Q => 
                           n6783, QN => n1575);
   OUT2_reg_0_inst : DFF_X1 port map( D => n7547, CK => CLK, Q => n6784, QN => 
                           n1512);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n7546, CK => CLK, Q => 
                           n6785, QN => n1576);
   OUT2_tri_0_inst : TBUF_X1 port map( A => n6784, EN => n6785, Z => OUT2(0));
   OUT2_tri_1_inst : TBUF_X1 port map( A => n6782, EN => n6783, Z => OUT2(1));
   OUT2_tri_2_inst : TBUF_X1 port map( A => n6780, EN => n6781, Z => OUT2(2));
   OUT2_tri_3_inst : TBUF_X1 port map( A => n6778, EN => n6779, Z => OUT2(3));
   OUT2_tri_4_inst : TBUF_X1 port map( A => n6776, EN => n6777, Z => OUT2(4));
   OUT2_tri_5_inst : TBUF_X1 port map( A => n6774, EN => n6775, Z => OUT2(5));
   OUT2_tri_6_inst : TBUF_X1 port map( A => n6772, EN => n6773, Z => OUT2(6));
   OUT2_tri_7_inst : TBUF_X1 port map( A => n6770, EN => n6771, Z => OUT2(7));
   OUT2_tri_8_inst : TBUF_X1 port map( A => n6768, EN => n6769, Z => OUT2(8));
   OUT2_tri_9_inst : TBUF_X1 port map( A => n6766, EN => n6767, Z => OUT2(9));
   OUT2_tri_10_inst : TBUF_X1 port map( A => n6764, EN => n6765, Z => OUT2(10))
                           ;
   OUT2_tri_11_inst : TBUF_X1 port map( A => n6762, EN => n6763, Z => OUT2(11))
                           ;
   OUT2_tri_12_inst : TBUF_X1 port map( A => n6760, EN => n6761, Z => OUT2(12))
                           ;
   OUT2_tri_13_inst : TBUF_X1 port map( A => n6758, EN => n6759, Z => OUT2(13))
                           ;
   OUT2_tri_14_inst : TBUF_X1 port map( A => n6756, EN => n6757, Z => OUT2(14))
                           ;
   OUT2_tri_15_inst : TBUF_X1 port map( A => n6754, EN => n6755, Z => OUT2(15))
                           ;
   OUT2_tri_16_inst : TBUF_X1 port map( A => n6752, EN => n6753, Z => OUT2(16))
                           ;
   OUT2_tri_17_inst : TBUF_X1 port map( A => n6750, EN => n6751, Z => OUT2(17))
                           ;
   OUT2_tri_18_inst : TBUF_X1 port map( A => n6748, EN => n6749, Z => OUT2(18))
                           ;
   OUT2_tri_19_inst : TBUF_X1 port map( A => n6746, EN => n6747, Z => OUT2(19))
                           ;
   OUT2_tri_20_inst : TBUF_X1 port map( A => n6744, EN => n6745, Z => OUT2(20))
                           ;
   OUT2_tri_21_inst : TBUF_X1 port map( A => n6742, EN => n6743, Z => OUT2(21))
                           ;
   OUT2_tri_22_inst : TBUF_X1 port map( A => n6740, EN => n6741, Z => OUT2(22))
                           ;
   OUT2_tri_23_inst : TBUF_X1 port map( A => n6738, EN => n6739, Z => OUT2(23))
                           ;
   OUT2_tri_24_inst : TBUF_X1 port map( A => n6736, EN => n6737, Z => OUT2(24))
                           ;
   OUT2_tri_25_inst : TBUF_X1 port map( A => n6734, EN => n6735, Z => OUT2(25))
                           ;
   OUT2_tri_26_inst : TBUF_X1 port map( A => n6732, EN => n6733, Z => OUT2(26))
                           ;
   OUT2_tri_27_inst : TBUF_X1 port map( A => n6730, EN => n6731, Z => OUT2(27))
                           ;
   OUT2_tri_28_inst : TBUF_X1 port map( A => n6728, EN => n6729, Z => OUT2(28))
                           ;
   OUT2_tri_29_inst : TBUF_X1 port map( A => n6726, EN => n6727, Z => OUT2(29))
                           ;
   OUT2_tri_30_inst : TBUF_X1 port map( A => n6724, EN => n6725, Z => OUT2(30))
                           ;
   OUT2_tri_31_inst : TBUF_X1 port map( A => n6722, EN => n6723, Z => OUT2(31))
                           ;
   OUT1_tri_0_inst : TBUF_X1 port map( A => n6720, EN => n6721, Z => OUT1(0));
   OUT1_tri_1_inst : TBUF_X1 port map( A => n6718, EN => n6719, Z => OUT1(1));
   OUT1_tri_2_inst : TBUF_X1 port map( A => n6716, EN => n6717, Z => OUT1(2));
   OUT1_tri_3_inst : TBUF_X1 port map( A => n6714, EN => n6715, Z => OUT1(3));
   OUT1_tri_4_inst : TBUF_X1 port map( A => n6712, EN => n6713, Z => OUT1(4));
   OUT1_tri_5_inst : TBUF_X1 port map( A => n6710, EN => n6711, Z => OUT1(5));
   OUT1_tri_6_inst : TBUF_X1 port map( A => n6708, EN => n6709, Z => OUT1(6));
   OUT1_tri_7_inst : TBUF_X1 port map( A => n6706, EN => n6707, Z => OUT1(7));
   OUT1_tri_8_inst : TBUF_X1 port map( A => n6704, EN => n6705, Z => OUT1(8));
   OUT1_tri_9_inst : TBUF_X1 port map( A => n6702, EN => n6703, Z => OUT1(9));
   OUT1_tri_10_inst : TBUF_X1 port map( A => n6700, EN => n6701, Z => OUT1(10))
                           ;
   OUT1_tri_11_inst : TBUF_X1 port map( A => n6698, EN => n6699, Z => OUT1(11))
                           ;
   OUT1_tri_12_inst : TBUF_X1 port map( A => n6696, EN => n6697, Z => OUT1(12))
                           ;
   OUT1_tri_13_inst : TBUF_X1 port map( A => n6694, EN => n6695, Z => OUT1(13))
                           ;
   OUT1_tri_14_inst : TBUF_X1 port map( A => n6692, EN => n6693, Z => OUT1(14))
                           ;
   OUT1_tri_15_inst : TBUF_X1 port map( A => n6690, EN => n6691, Z => OUT1(15))
                           ;
   OUT1_tri_16_inst : TBUF_X1 port map( A => n6688, EN => n6689, Z => OUT1(16))
                           ;
   OUT1_tri_17_inst : TBUF_X1 port map( A => n6686, EN => n6687, Z => OUT1(17))
                           ;
   OUT1_tri_18_inst : TBUF_X1 port map( A => n6684, EN => n6685, Z => OUT1(18))
                           ;
   OUT1_tri_19_inst : TBUF_X1 port map( A => n6682, EN => n6683, Z => OUT1(19))
                           ;
   OUT1_tri_20_inst : TBUF_X1 port map( A => n6680, EN => n6681, Z => OUT1(20))
                           ;
   OUT1_tri_21_inst : TBUF_X1 port map( A => n6678, EN => n6679, Z => OUT1(21))
                           ;
   OUT1_tri_22_inst : TBUF_X1 port map( A => n6676, EN => n6677, Z => OUT1(22))
                           ;
   OUT1_tri_23_inst : TBUF_X1 port map( A => n6674, EN => n6675, Z => OUT1(23))
                           ;
   OUT1_tri_24_inst : TBUF_X1 port map( A => n6672, EN => n6673, Z => OUT1(24))
                           ;
   OUT1_tri_25_inst : TBUF_X1 port map( A => n6670, EN => n6671, Z => OUT1(25))
                           ;
   OUT1_tri_26_inst : TBUF_X1 port map( A => n6668, EN => n6669, Z => OUT1(26))
                           ;
   OUT1_tri_27_inst : TBUF_X1 port map( A => n6666, EN => n6667, Z => OUT1(27))
                           ;
   OUT1_tri_28_inst : TBUF_X1 port map( A => n6664, EN => n6665, Z => OUT1(28))
                           ;
   OUT1_tri_29_inst : TBUF_X1 port map( A => n6662, EN => n6663, Z => OUT1(29))
                           ;
   OUT1_tri_30_inst : TBUF_X1 port map( A => n6660, EN => n6661, Z => OUT1(30))
                           ;
   OUT1_tri_31_inst : TBUF_X1 port map( A => n6658, EN => n6659, Z => OUT1(31))
                           ;
   U3 : AND2_X1 port map( A1 => DATAIN(23), A2 => n1946, ZN => n385);
   U4 : AND2_X1 port map( A1 => DATAIN(22), A2 => n1946, ZN => n386);
   U5 : AND2_X1 port map( A1 => DATAIN(21), A2 => n1946, ZN => n387);
   U6 : AND2_X1 port map( A1 => DATAIN(20), A2 => n1946, ZN => n388);
   U7 : AND2_X1 port map( A1 => DATAIN(19), A2 => n1946, ZN => n389);
   U8 : AND2_X1 port map( A1 => DATAIN(18), A2 => n1946, ZN => n390);
   U9 : AND2_X1 port map( A1 => DATAIN(17), A2 => n1946, ZN => n391);
   U10 : AND2_X1 port map( A1 => DATAIN(16), A2 => n1946, ZN => n392);
   U11 : AND2_X1 port map( A1 => DATAIN(15), A2 => n1946, ZN => n393);
   U12 : AND2_X1 port map( A1 => DATAIN(14), A2 => n1946, ZN => n394);
   U13 : AND2_X1 port map( A1 => DATAIN(13), A2 => n1946, ZN => n395);
   U14 : AND2_X1 port map( A1 => DATAIN(12), A2 => n1946, ZN => n396);
   U15 : AND2_X1 port map( A1 => DATAIN(11), A2 => n1946, ZN => n397);
   U16 : AND2_X1 port map( A1 => DATAIN(10), A2 => n1946, ZN => n398);
   U17 : AND2_X1 port map( A1 => DATAIN(9), A2 => n1946, ZN => n399);
   U18 : AND2_X1 port map( A1 => DATAIN(8), A2 => n1946, ZN => n400);
   U19 : AND2_X1 port map( A1 => DATAIN(7), A2 => n1946, ZN => n401);
   U20 : AND2_X1 port map( A1 => DATAIN(6), A2 => n1946, ZN => n402);
   U21 : AND2_X1 port map( A1 => DATAIN(5), A2 => n1946, ZN => n403);
   U22 : AND2_X1 port map( A1 => DATAIN(4), A2 => n1946, ZN => n404);
   U23 : AND2_X1 port map( A1 => DATAIN(3), A2 => n1946, ZN => n405);
   U24 : AND2_X1 port map( A1 => DATAIN(2), A2 => n1946, ZN => n406);
   U25 : AND2_X1 port map( A1 => DATAIN(1), A2 => n1946, ZN => n407);
   U26 : AND2_X1 port map( A1 => n1816, A2 => n1772, ZN => n408);
   U27 : AND2_X1 port map( A1 => n3216, A2 => n3207, ZN => n409);
   U28 : AND2_X1 port map( A1 => n4500, A2 => n4491, ZN => n410);
   U29 : NAND2_X2 port map( A1 => n3246, A2 => n3211, ZN => n411);
   U30 : NAND2_X2 port map( A1 => n3203, A2 => n3212, ZN => n412);
   U31 : NAND2_X2 port map( A1 => n4490, A2 => n4495, ZN => n413);
   U32 : NAND2_X2 port map( A1 => n4500, A2 => n4488, ZN => n414);
   U33 : NAND2_X2 port map( A1 => n4487, A2 => n4497, ZN => n415);
   U34 : NAND2_X2 port map( A1 => n3223, A2 => n3212, ZN => n416);
   U35 : NAND2_X2 port map( A1 => n3224, A2 => n1750, ZN => n417);
   U36 : NAND2_X2 port map( A1 => n3234, A2 => n3208, ZN => n418);
   U37 : NAND2_X2 port map( A1 => n3236, A2 => n3211, ZN => n419);
   U38 : AND2_X1 port map( A1 => n3207, A2 => ADD_RD1(6), ZN => n420);
   U39 : NAND2_X2 port map( A1 => n4487, A2 => n4488, ZN => n421);
   U40 : NAND2_X2 port map( A1 => n4508, A2 => n4495, ZN => n422);
   U41 : NAND2_X2 port map( A1 => n4518, A2 => n4492, ZN => n423);
   U42 : NAND2_X2 port map( A1 => n4530, A2 => n4493, ZN => n424);
   U43 : NOR3_X2 port map( A1 => n3248, A2 => ADD_RD1(1), A3 => n3249, ZN => 
                           n3208);
   U44 : NOR3_X2 port map( A1 => n4534, A2 => n4532, A3 => n4533, ZN => n4491);
   U45 : NOR3_X2 port map( A1 => n3250, A2 => n3248, A3 => n3249, ZN => n3207);
   U46 : NOR3_X2 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n3248, ZN 
                           => n3204);
   U47 : NOR3_X2 port map( A1 => n4532, A2 => ADD_RD2(1), A3 => n4533, ZN => 
                           n4492);
   U48 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n4534, ZN 
                           => n4495);
   U49 : NOR3_X2 port map( A1 => n4534, A2 => ADD_RD2(0), A3 => n4533, ZN => 
                           n4493);
   U50 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n4532, ZN 
                           => n4488);
   U51 : AND2_X2 port map( A1 => n3211, A2 => ADD_RD1(6), ZN => n2032);
   U52 : AND2_X2 port map( A1 => n4490, A2 => n4497, ZN => n3280);
   U53 : AND2_X2 port map( A1 => n4507, A2 => n4489, ZN => n3297);
   U54 : INV_X2 port map( A => n420, ZN => n1577);
   U55 : NAND2_X2 port map( A1 => n1951, A2 => n1948, ZN => n1950);
   U56 : INV_X2 port map( A => n409, ZN => n1578);
   U57 : NAND2_X2 port map( A1 => n3266, A2 => n3263, ZN => n3265);
   U58 : INV_X2 port map( A => n410, ZN => n1579);
   U59 : NAND2_X2 port map( A1 => n1819, A2 => n1811, ZN => n1844);
   U60 : NAND2_X2 port map( A1 => n1819, A2 => n1814, ZN => n1846);
   U61 : NAND2_X2 port map( A1 => n1819, A2 => n1816, ZN => n1848);
   U62 : NAND2_X2 port map( A1 => n1853, A2 => n1771, ZN => n1851);
   U63 : NAND2_X2 port map( A1 => n1853, A2 => n1775, ZN => n1854);
   U64 : NAND2_X2 port map( A1 => n1853, A2 => n1778, ZN => n1856);
   U65 : NAND2_X2 port map( A1 => n1853, A2 => n1781, ZN => n1858);
   U66 : NAND2_X2 port map( A1 => n1853, A2 => n1784, ZN => n1860);
   U67 : NAND2_X2 port map( A1 => n1853, A2 => n1787, ZN => n1862);
   U68 : NAND2_X2 port map( A1 => n1853, A2 => n1790, ZN => n1864);
   U69 : NAND2_X2 port map( A1 => n1853, A2 => n1793, ZN => n1866);
   U70 : NAND2_X2 port map( A1 => n1853, A2 => n1796, ZN => n1868);
   U71 : NAND2_X2 port map( A1 => n1853, A2 => n1799, ZN => n1870);
   U72 : NAND2_X2 port map( A1 => n1853, A2 => n1802, ZN => n1872);
   U73 : NAND2_X2 port map( A1 => n1853, A2 => n1805, ZN => n1874);
   U74 : NAND2_X2 port map( A1 => n1853, A2 => n1808, ZN => n1876);
   U75 : NAND2_X2 port map( A1 => n1853, A2 => n1811, ZN => n1878);
   U76 : NAND2_X2 port map( A1 => n1853, A2 => n1814, ZN => n1880);
   U77 : NAND2_X2 port map( A1 => n1853, A2 => n1816, ZN => n1882);
   U78 : NOR3_X4 port map( A1 => ADD_WR(4), A2 => ADD_WR(6), A3 => n1884, ZN =>
                           n1853);
   U79 : NAND2_X2 port map( A1 => n1887, A2 => n1771, ZN => n1885);
   U80 : NAND2_X2 port map( A1 => n1887, A2 => n1775, ZN => n1888);
   U81 : NAND2_X2 port map( A1 => n1887, A2 => n1778, ZN => n1890);
   U82 : NAND2_X2 port map( A1 => n1887, A2 => n1781, ZN => n1892);
   U83 : NAND2_X2 port map( A1 => n1887, A2 => n1784, ZN => n1894);
   U84 : NAND2_X2 port map( A1 => n1887, A2 => n1787, ZN => n1896);
   U85 : NAND2_X2 port map( A1 => n1887, A2 => n1790, ZN => n1898);
   U86 : NAND2_X2 port map( A1 => n1887, A2 => n1793, ZN => n1900);
   U87 : NAND2_X2 port map( A1 => n1887, A2 => n1796, ZN => n1902);
   U88 : NAND2_X2 port map( A1 => n1887, A2 => n1799, ZN => n1906);
   U89 : NAND2_X2 port map( A1 => n1887, A2 => n1802, ZN => n1909);
   U90 : NAND2_X2 port map( A1 => n1887, A2 => n1805, ZN => n1912);
   U91 : NAND2_X2 port map( A1 => n1887, A2 => n1808, ZN => n1916);
   U92 : NAND2_X2 port map( A1 => n1887, A2 => n1811, ZN => n1919);
   U93 : NAND2_X2 port map( A1 => n1887, A2 => n1814, ZN => n1921);
   U94 : NAND2_X2 port map( A1 => n1887, A2 => n1816, ZN => n1923);
   U95 : NOR3_X4 port map( A1 => n1850, A2 => ADD_WR(6), A3 => n1884, ZN => 
                           n1887);
   U96 : NAND2_X2 port map( A1 => n1819, A2 => n1805, ZN => n1840);
   U97 : NAND2_X2 port map( A1 => n1819, A2 => n1808, ZN => n1842);
   U98 : NAND2_X2 port map( A1 => n1819, A2 => n1799, ZN => n1836);
   U99 : NAND2_X2 port map( A1 => n1819, A2 => n1802, ZN => n1838);
   U100 : NAND2_X2 port map( A1 => n1819, A2 => n1793, ZN => n1832);
   U101 : NAND2_X2 port map( A1 => n1819, A2 => n1796, ZN => n1834);
   U102 : NAND2_X2 port map( A1 => n1819, A2 => n1787, ZN => n1828);
   U103 : NAND2_X2 port map( A1 => n1819, A2 => n1790, ZN => n1830);
   U104 : NAND2_X2 port map( A1 => n1819, A2 => n1781, ZN => n1824);
   U105 : NAND2_X2 port map( A1 => n1819, A2 => n1784, ZN => n1826);
   U106 : NAND2_X2 port map( A1 => n1819, A2 => n1775, ZN => n1820);
   U107 : NAND2_X2 port map( A1 => n1819, A2 => n1778, ZN => n1822);
   U108 : INV_X2 port map( A => n408, ZN => n1580);
   U109 : NAND2_X2 port map( A1 => n1819, A2 => n1771, ZN => n1817);
   U110 : NOR3_X4 port map( A1 => ADD_WR(5), A2 => ADD_WR(6), A3 => n1850, ZN 
                           => n1819);
   U111 : NAND2_X2 port map( A1 => n1811, A2 => n1772, ZN => n1809);
   U112 : NAND2_X2 port map( A1 => n1814, A2 => n1772, ZN => n1812);
   U113 : NAND2_X2 port map( A1 => n1805, A2 => n1772, ZN => n1803);
   U114 : NAND2_X2 port map( A1 => n1808, A2 => n1772, ZN => n1806);
   U115 : NAND2_X2 port map( A1 => n1799, A2 => n1772, ZN => n1797);
   U116 : NAND2_X2 port map( A1 => n1802, A2 => n1772, ZN => n1800);
   U117 : NAND2_X2 port map( A1 => n1793, A2 => n1772, ZN => n1791);
   U118 : NAND2_X2 port map( A1 => n1796, A2 => n1772, ZN => n1794);
   U119 : NAND2_X2 port map( A1 => n1787, A2 => n1772, ZN => n1785);
   U120 : NAND2_X2 port map( A1 => n1790, A2 => n1772, ZN => n1788);
   U121 : NAND2_X2 port map( A1 => n1781, A2 => n1772, ZN => n1779);
   U122 : NAND2_X2 port map( A1 => n1784, A2 => n1772, ZN => n1782);
   U123 : NAND2_X2 port map( A1 => n1775, A2 => n1772, ZN => n1773);
   U124 : NAND2_X2 port map( A1 => n1778, A2 => n1772, ZN => n1776);
   U125 : NAND2_X2 port map( A1 => n1771, A2 => n1772, ZN => n1758);
   U126 : NOR3_X4 port map( A1 => ADD_WR(5), A2 => ADD_WR(6), A3 => ADD_WR(4), 
                           ZN => n1772);
   U127 : INV_X1 port map( A => n1942, ZN => n1581);
   U128 : INV_X2 port map( A => n1581, ZN => n1582);
   U129 : INV_X1 port map( A => n1944, ZN => n1583);
   U130 : INV_X2 port map( A => n1583, ZN => n1584);
   U131 : INV_X1 port map( A => n1932, ZN => n1585);
   U132 : INV_X2 port map( A => n1585, ZN => n1586);
   U133 : INV_X1 port map( A => n1939, ZN => n1587);
   U134 : INV_X2 port map( A => n1587, ZN => n1588);
   U135 : INV_X1 port map( A => n1922, ZN => n1589);
   U136 : INV_X2 port map( A => n1589, ZN => n1590);
   U137 : INV_X1 port map( A => n1930, ZN => n1591);
   U138 : INV_X2 port map( A => n1591, ZN => n1592);
   U139 : INV_X1 port map( A => n1917, ZN => n1593);
   U140 : INV_X2 port map( A => n1593, ZN => n1594);
   U141 : INV_X1 port map( A => n1920, ZN => n1595);
   U142 : INV_X2 port map( A => n1595, ZN => n1596);
   U143 : INV_X1 port map( A => n1899, ZN => n1597);
   U144 : INV_X2 port map( A => n1597, ZN => n1598);
   U145 : INV_X1 port map( A => n1901, ZN => n1599);
   U146 : INV_X2 port map( A => n1599, ZN => n1600);
   U147 : INV_X1 port map( A => n1895, ZN => n1601);
   U148 : INV_X2 port map( A => n1601, ZN => n1602);
   U149 : INV_X1 port map( A => n1897, ZN => n1603);
   U150 : INV_X2 port map( A => n1603, ZN => n1604);
   U151 : INV_X1 port map( A => n1886, ZN => n1605);
   U152 : INV_X2 port map( A => n1605, ZN => n1606);
   U153 : INV_X1 port map( A => n1893, ZN => n1607);
   U154 : INV_X2 port map( A => n1607, ZN => n1608);
   U155 : INV_X1 port map( A => n1877, ZN => n1609);
   U156 : INV_X2 port map( A => n1609, ZN => n1610);
   U157 : INV_X1 port map( A => n1883, ZN => n1611);
   U158 : INV_X2 port map( A => n1611, ZN => n1612);
   U159 : INV_X1 port map( A => n1873, ZN => n1613);
   U160 : INV_X2 port map( A => n1613, ZN => n1614);
   U161 : INV_X1 port map( A => n1875, ZN => n1615);
   U162 : INV_X2 port map( A => n1615, ZN => n1616);
   U163 : INV_X1 port map( A => n1865, ZN => n1617);
   U164 : INV_X2 port map( A => n1617, ZN => n1618);
   U165 : INV_X1 port map( A => n1867, ZN => n1619);
   U166 : INV_X2 port map( A => n1619, ZN => n1620);
   U167 : INV_X1 port map( A => n1857, ZN => n1621);
   U168 : INV_X2 port map( A => n1621, ZN => n1622);
   U169 : INV_X1 port map( A => n1859, ZN => n1623);
   U170 : INV_X2 port map( A => n1623, ZN => n1624);
   U171 : INV_X1 port map( A => n1847, ZN => n1625);
   U172 : INV_X2 port map( A => n1625, ZN => n1626);
   U173 : INV_X1 port map( A => n1855, ZN => n1627);
   U174 : INV_X2 port map( A => n1627, ZN => n1628);
   U175 : INV_X1 port map( A => n1839, ZN => n1629);
   U176 : INV_X2 port map( A => n1629, ZN => n1630);
   U177 : INV_X1 port map( A => n1845, ZN => n1631);
   U178 : INV_X2 port map( A => n1631, ZN => n1632);
   U179 : INV_X1 port map( A => n1835, ZN => n1633);
   U180 : INV_X2 port map( A => n1633, ZN => n1634);
   U181 : INV_X1 port map( A => n1837, ZN => n1635);
   U182 : INV_X2 port map( A => n1635, ZN => n1636);
   U183 : INV_X1 port map( A => n1827, ZN => n1637);
   U184 : INV_X2 port map( A => n1637, ZN => n1638);
   U185 : INV_X1 port map( A => n1829, ZN => n1639);
   U186 : INV_X2 port map( A => n1639, ZN => n1640);
   U187 : INV_X1 port map( A => n1818, ZN => n1641);
   U188 : INV_X2 port map( A => n1641, ZN => n1642);
   U189 : INV_X1 port map( A => n1821, ZN => n1643);
   U190 : INV_X2 port map( A => n1643, ZN => n1644);
   U191 : INV_X1 port map( A => n1807, ZN => n1645);
   U192 : INV_X2 port map( A => n1645, ZN => n1646);
   U193 : INV_X1 port map( A => n1815, ZN => n1647);
   U194 : INV_X2 port map( A => n1647, ZN => n1648);
   U195 : INV_X1 port map( A => n1795, ZN => n1649);
   U196 : INV_X2 port map( A => n1649, ZN => n1650);
   U197 : INV_X1 port map( A => n1804, ZN => n1651);
   U198 : INV_X2 port map( A => n1651, ZN => n1652);
   U199 : INV_X1 port map( A => n1789, ZN => n1653);
   U200 : INV_X2 port map( A => n1653, ZN => n1654);
   U201 : INV_X1 port map( A => n1792, ZN => n1655);
   U202 : INV_X2 port map( A => n1655, ZN => n1656);
   U203 : INV_X1 port map( A => n1777, ZN => n1657);
   U204 : INV_X2 port map( A => n1657, ZN => n1658);
   U205 : INV_X1 port map( A => n1780, ZN => n1659);
   U206 : INV_X2 port map( A => n1659, ZN => n1660);
   U207 : INV_X1 port map( A => n1934, ZN => n1661);
   U208 : INV_X2 port map( A => n1661, ZN => n1662);
   U209 : INV_X1 port map( A => n1936, ZN => n1663);
   U210 : INV_X2 port map( A => n1663, ZN => n1664);
   U211 : INV_X1 port map( A => n1924, ZN => n1665);
   U212 : INV_X2 port map( A => n1665, ZN => n1666);
   U213 : INV_X1 port map( A => n1926, ZN => n1667);
   U214 : INV_X2 port map( A => n1667, ZN => n1668);
   U215 : INV_X1 port map( A => n1910, ZN => n1669);
   U216 : INV_X2 port map( A => n1669, ZN => n1670);
   U217 : INV_X1 port map( A => n1913, ZN => n1671);
   U218 : INV_X2 port map( A => n1671, ZN => n1672);
   U219 : INV_X1 port map( A => n1903, ZN => n1673);
   U220 : INV_X2 port map( A => n1673, ZN => n1674);
   U221 : INV_X1 port map( A => n1907, ZN => n1675);
   U222 : INV_X2 port map( A => n1675, ZN => n1676);
   U223 : INV_X1 port map( A => n1889, ZN => n1677);
   U224 : INV_X2 port map( A => n1677, ZN => n1678);
   U225 : INV_X1 port map( A => n1891, ZN => n1679);
   U226 : INV_X2 port map( A => n1679, ZN => n1680);
   U227 : INV_X1 port map( A => n1879, ZN => n1681);
   U228 : INV_X2 port map( A => n1681, ZN => n1682);
   U229 : INV_X1 port map( A => n1881, ZN => n1683);
   U230 : INV_X2 port map( A => n1683, ZN => n1684);
   U231 : INV_X1 port map( A => n1869, ZN => n1685);
   U232 : INV_X2 port map( A => n1685, ZN => n1686);
   U233 : INV_X1 port map( A => n1871, ZN => n1687);
   U234 : INV_X2 port map( A => n1687, ZN => n1688);
   U235 : INV_X1 port map( A => n1861, ZN => n1689);
   U236 : INV_X2 port map( A => n1689, ZN => n1690);
   U237 : INV_X1 port map( A => n1863, ZN => n1691);
   U238 : INV_X2 port map( A => n1691, ZN => n1692);
   U239 : INV_X1 port map( A => n1849, ZN => n1693);
   U240 : INV_X2 port map( A => n1693, ZN => n1694);
   U241 : INV_X1 port map( A => n1852, ZN => n1695);
   U242 : INV_X2 port map( A => n1695, ZN => n1696);
   U243 : INV_X1 port map( A => n1841, ZN => n1697);
   U244 : INV_X2 port map( A => n1697, ZN => n1698);
   U245 : INV_X1 port map( A => n1843, ZN => n1699);
   U246 : INV_X2 port map( A => n1699, ZN => n1700);
   U247 : INV_X1 port map( A => n1831, ZN => n1701);
   U248 : INV_X2 port map( A => n1701, ZN => n1702);
   U249 : INV_X1 port map( A => n1833, ZN => n1703);
   U250 : INV_X2 port map( A => n1703, ZN => n1704);
   U251 : INV_X1 port map( A => n1823, ZN => n1705);
   U252 : INV_X2 port map( A => n1705, ZN => n1706);
   U253 : INV_X1 port map( A => n1825, ZN => n1707);
   U254 : INV_X2 port map( A => n1707, ZN => n1708);
   U255 : INV_X1 port map( A => n1810, ZN => n1709);
   U256 : INV_X2 port map( A => n1709, ZN => n1710);
   U257 : INV_X1 port map( A => n1813, ZN => n1711);
   U258 : INV_X2 port map( A => n1711, ZN => n1712);
   U259 : INV_X1 port map( A => n1798, ZN => n1713);
   U260 : INV_X2 port map( A => n1713, ZN => n1714);
   U261 : INV_X1 port map( A => n1801, ZN => n1715);
   U262 : INV_X2 port map( A => n1715, ZN => n1716);
   U263 : INV_X1 port map( A => n1783, ZN => n1717);
   U264 : INV_X2 port map( A => n1717, ZN => n1718);
   U265 : INV_X1 port map( A => n1786, ZN => n1719);
   U266 : INV_X2 port map( A => n1719, ZN => n1720);
   U267 : INV_X1 port map( A => n1760, ZN => n1721);
   U268 : INV_X2 port map( A => n1721, ZN => n1722);
   U269 : INV_X1 port map( A => n1774, ZN => n1723);
   U270 : INV_X2 port map( A => n1723, ZN => n1724);
   U271 : INV_X4 port map( A => n407, ZN => n1725);
   U272 : INV_X4 port map( A => RESET, ZN => n1770);
   U273 : NAND2_X4 port map( A1 => ENABLE, A2 => n3262, ZN => n1951);
   U274 : NAND2_X4 port map( A1 => ENABLE, A2 => n4545, ZN => n3266);
   U275 : INV_X4 port map( A => n403, ZN => n1726);
   U276 : INV_X4 port map( A => n404, ZN => n1727);
   U277 : INV_X4 port map( A => n405, ZN => n1728);
   U278 : INV_X4 port map( A => n406, ZN => n1729);
   U279 : INV_X4 port map( A => n399, ZN => n1730);
   U280 : INV_X4 port map( A => n400, ZN => n1731);
   U281 : INV_X4 port map( A => n401, ZN => n1732);
   U282 : INV_X4 port map( A => n402, ZN => n1733);
   U283 : INV_X4 port map( A => n395, ZN => n1734);
   U284 : INV_X4 port map( A => n396, ZN => n1735);
   U285 : INV_X4 port map( A => n397, ZN => n1736);
   U286 : INV_X4 port map( A => n398, ZN => n1737);
   U287 : INV_X4 port map( A => n391, ZN => n1738);
   U288 : INV_X4 port map( A => n392, ZN => n1739);
   U289 : INV_X4 port map( A => n393, ZN => n1740);
   U290 : INV_X4 port map( A => n394, ZN => n1741);
   U291 : INV_X4 port map( A => n387, ZN => n1742);
   U292 : INV_X4 port map( A => n388, ZN => n1743);
   U293 : INV_X4 port map( A => n389, ZN => n1744);
   U294 : INV_X4 port map( A => n390, ZN => n1745);
   U295 : INV_X4 port map( A => n385, ZN => n1746);
   U296 : INV_X4 port map( A => n386, ZN => n1747);
   U297 : NAND2_X4 port map( A1 => DATAIN(25), A2 => n1946, ZN => n1766);
   U298 : NAND2_X4 port map( A1 => DATAIN(24), A2 => n1946, ZN => n1767);
   U299 : NAND2_X4 port map( A1 => DATAIN(29), A2 => n1946, ZN => n1762);
   U300 : NAND2_X4 port map( A1 => DATAIN(28), A2 => n1946, ZN => n1763);
   U301 : NAND2_X4 port map( A1 => DATAIN(27), A2 => n1946, ZN => n1764);
   U302 : NAND2_X4 port map( A1 => DATAIN(26), A2 => n1946, ZN => n1765);
   U303 : INV_X2 port map( A => n1769, ZN => n1946);
   U304 : NAND2_X4 port map( A1 => WR, A2 => ENABLE, ZN => n1769);
   U305 : NAND2_X4 port map( A1 => DATAIN(0), A2 => n1946, ZN => n1768);
   U306 : NAND2_X4 port map( A1 => DATAIN(31), A2 => n1946, ZN => n1759);
   U307 : NAND2_X4 port map( A1 => DATAIN(30), A2 => n1946, ZN => n1761);
   U308 : NAND2_X2 port map( A1 => n3216, A2 => n3212, ZN => n1980);
   U309 : NOR3_X2 port map( A1 => n3248, A2 => ADD_RD1(2), A3 => n3250, ZN => 
                           n3212);
   U310 : NOR3_X2 port map( A1 => n4532, A2 => ADD_RD2(2), A3 => n4534, ZN => 
                           n4497);
   U311 : NOR3_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n3249, ZN
                           => n3211);
   U312 : AND2_X2 port map( A1 => n3216, A2 => n3208, ZN => n1971);
   U313 : AND2_X2 port map( A1 => n3234, A2 => n1750, ZN => n2008);
   U314 : CLKBUF_X1 port map( A => n3275, Z => n1748);
   U315 : AND2_X2 port map( A1 => n4518, A2 => n4495, ZN => n3321);
   U316 : CLKBUF_X1 port map( A => n2047, Z => n1749);
   U317 : AND2_X2 port map( A1 => n4487, A2 => n4496, ZN => n3313);
   U318 : AND2_X2 port map( A1 => n4508, A2 => n4492, ZN => n3303);
   U319 : AND2_X2 port map( A1 => n4520, A2 => n4488, ZN => n3331);
   U320 : AND2_X2 port map( A1 => n4530, A2 => n4489, ZN => n3362);
   U321 : CLKBUF_X1 port map( A => n3213, Z => n1750);
   U322 : AND2_X2 port map( A1 => n3206, A2 => n1750, ZN => n1966);
   U323 : AND2_X2 port map( A1 => n4500, A2 => n4495, ZN => n3289);
   U324 : AND2_X2 port map( A1 => n4496, A2 => ADD_RD2(6), ZN => n3346);
   U325 : AND2_X2 port map( A1 => n3203, A2 => n3211, ZN => n2000);
   U326 : CLKBUF_X1 port map( A => n2018, Z => n1751);
   U327 : CLKBUF_X1 port map( A => n2042, Z => n1752);
   U328 : AND2_X2 port map( A1 => n4507, A2 => n4493, ZN => n3337);
   U329 : AND2_X2 port map( A1 => n4520, A2 => n4491, ZN => n3326);
   U330 : CLKBUF_X1 port map( A => n3357, Z => n1753);
   U331 : NAND2_X2 port map( A1 => n3206, A2 => n1755, ZN => n1975);
   U332 : NAND2_X2 port map( A1 => n1927, A2 => n1775, ZN => n1929);
   U333 : NAND2_X2 port map( A1 => n4500, A2 => n4489, ZN => n3292);
   U334 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n4489);
   U335 : AND2_X2 port map( A1 => n3216, A2 => n3204, ZN => n1976);
   U336 : CLKBUF_X1 port map( A => n3284, Z => n1754);
   U337 : AND2_X2 port map( A1 => n3203, A2 => n3207, ZN => n1995);
   U338 : NAND2_X2 port map( A1 => n4507, A2 => n4497, ZN => n3302);
   U339 : NAND2_X2 port map( A1 => n3246, A2 => n1757, ZN => n2046);
   U340 : NAND2_X2 port map( A1 => n4520, A2 => n4496, ZN => n3336);
   U341 : NAND2_X2 port map( A1 => n3206, A2 => n3212, ZN => n1969);
   U342 : NAND2_X2 port map( A1 => n3223, A2 => n3208, ZN => n2026);
   U343 : NAND2_X2 port map( A1 => n4518, A2 => n4491, ZN => n3365);
   U344 : NAND2_X2 port map( A1 => n4488, A2 => ADD_RD2(6), ZN => n3355);
   U345 : AND2_X2 port map( A1 => n3246, A2 => n1755, ZN => n2048);
   U346 : NOR3_X2 port map( A1 => n3227, A2 => n3215, A3 => n3238, ZN => n3246)
                           ;
   U347 : NAND2_X2 port map( A1 => n1927, A2 => n1778, ZN => n1931);
   U348 : CLKBUF_X1 port map( A => n3205, Z => n1755);
   U349 : AND2_X2 port map( A1 => n1755, A2 => ADD_RD1(6), ZN => n2037);
   U350 : AND2_X2 port map( A1 => n3223, A2 => n1755, ZN => n1985);
   U351 : NAND2_X2 port map( A1 => n4530, A2 => n4496, ZN => n3360);
   U352 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n4533, ZN
                           => n4496);
   U353 : AND2_X2 port map( A1 => n4489, A2 => ADD_RD2(6), ZN => n3352);
   U354 : NAND2_X2 port map( A1 => n3204, A2 => ADD_RD1(6), ZN => n2040);
   U355 : NAND2_X2 port map( A1 => n4507, A2 => n4492, ZN => n3340);
   U356 : NAND2_X2 port map( A1 => n4520, A2 => n4493, ZN => n3329);
   U357 : AND2_X2 port map( A1 => n3216, A2 => n3211, ZN => n1972);
   U358 : AND2_X2 port map( A1 => n3206, A2 => n3208, ZN => n1961);
   U359 : AND2_X2 port map( A1 => n3224, A2 => n3207, ZN => n1986);
   U360 : AND2_X2 port map( A1 => n4508, A2 => n4491, ZN => n3298);
   U361 : AND2_X2 port map( A1 => n3246, A2 => n1750, ZN => n2043);
   U362 : NAND2_X2 port map( A1 => n1927, A2 => n1787, ZN => n1938);
   U363 : NAND2_X2 port map( A1 => n4491, A2 => ADD_RD2(6), ZN => n3351);
   U364 : AND2_X1 port map( A1 => n3216, A2 => n1750, ZN => n1979);
   U365 : INV_X2 port map( A => n1979, ZN => n1756);
   U366 : NAND2_X2 port map( A1 => n3236, A2 => n3207, ZN => n2016);
   U367 : NAND2_X2 port map( A1 => n3234, A2 => n1757, ZN => n2050);
   U368 : AND2_X2 port map( A1 => n3216, A2 => n1755, ZN => n1977);
   U369 : NOR4_X2 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(5), A4 => ADD_RD1(6), ZN => n3216);
   U370 : AND2_X2 port map( A1 => n3206, A2 => n3204, ZN => n1967);
   U371 : AND2_X2 port map( A1 => n4500, A2 => n4497, ZN => n3290);
   U372 : AND2_X2 port map( A1 => n4490, A2 => n4496, ZN => n3281);
   U373 : AND2_X2 port map( A1 => n4518, A2 => n4488, ZN => n3322);
   U374 : AND2_X2 port map( A1 => n3224, A2 => n3208, ZN => n1991);
   U375 : AND2_X2 port map( A1 => n4487, A2 => n4492, ZN => n3314);
   U376 : AND2_X2 port map( A1 => n4508, A2 => n4493, ZN => n3304);
   U377 : AND2_X2 port map( A1 => n4520, A2 => n4489, ZN => n3332);
   U378 : AND2_X2 port map( A1 => n4530, A2 => n4495, ZN => n3358);
   U379 : NAND2_X2 port map( A1 => n1927, A2 => n1790, ZN => n1941);
   U380 : CLKBUF_X1 port map( A => n3209, Z => n1757);
   U381 : AND2_X2 port map( A1 => n3224, A2 => n1757, ZN => n1990);
   U382 : AND2_X2 port map( A1 => n3236, A2 => n1757, ZN => n2013);
   U383 : AND2_X2 port map( A1 => n3223, A2 => n1757, ZN => n2023);
   U384 : NAND2_X2 port map( A1 => n3216, A2 => n1757, ZN => n1974);
   U385 : NAND2_X2 port map( A1 => n4508, A2 => n4496, ZN => n3306);
   U386 : AND2_X2 port map( A1 => n3234, A2 => n3204, ZN => n2009);
   U387 : AND2_X2 port map( A1 => n3212, A2 => ADD_RD1(6), ZN => n2033);
   U388 : AND2_X2 port map( A1 => n4490, A2 => n4492, ZN => n3276);
   U389 : AND2_X2 port map( A1 => n4497, A2 => ADD_RD2(6), ZN => n3347);
   U390 : AND2_X2 port map( A1 => n3203, A2 => n3208, ZN => n2001);
   U391 : AND2_X2 port map( A1 => n3223, A2 => n3207, ZN => n2024);
   U392 : AND2_X2 port map( A1 => n4507, A2 => n4491, ZN => n3338);
   U393 : AND2_X2 port map( A1 => n4518, A2 => n4489, ZN => n3327);
   U394 : AND2_X2 port map( A1 => n4530, A2 => n4488, ZN => n3363);
   U395 : NOR3_X2 port map( A1 => n4511, A2 => n4499, A3 => n4522, ZN => n4530)
                           ;
   U396 : NAND2_X2 port map( A1 => n4500, A2 => n4493, ZN => n3287);
   U397 : NAND2_X2 port map( A1 => n3224, A2 => n1755, ZN => n1998);
   U398 : NAND2_X2 port map( A1 => n3236, A2 => n1750, ZN => n2021);
   U399 : NAND2_X2 port map( A1 => n3206, A2 => n3211, ZN => n1970);
   U400 : NAND2_X2 port map( A1 => n4487, A2 => n4495, ZN => n3316);
   U401 : NAND2_X2 port map( A1 => n1927, A2 => n1771, ZN => n1925);
   U402 : AND2_X2 port map( A1 => n3206, A2 => n1757, ZN => n1960);
   U403 : NOR3_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), A3 => n3215, ZN
                           => n3206);
   U404 : AND2_X2 port map( A1 => n4487, A2 => n4491, ZN => n3308);
   U405 : AND2_X2 port map( A1 => n4500, A2 => n4496, ZN => n3285);
   U406 : NOR4_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(5), A4 => ADD_RD2(6), ZN => n4500);
   U407 : AND2_X2 port map( A1 => n3236, A2 => n1755, ZN => n2019);
   U408 : AND2_X2 port map( A1 => n3246, A2 => n3207, ZN => n2038);
   U409 : AND2_X2 port map( A1 => n4487, A2 => n4493, ZN => n3309);
   U410 : NOR3_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(5), A3 => n4511, ZN
                           => n4487);
   U411 : NAND2_X2 port map( A1 => n3223, A2 => n3204, ZN => n1988);
   U412 : NAND2_X2 port map( A1 => n3234, A2 => n3212, ZN => n2011);
   U413 : NAND2_X2 port map( A1 => n3208, A2 => ADD_RD1(6), ZN => n2035);
   U414 : NAND2_X2 port map( A1 => n4507, A2 => n4488, ZN => n3300);
   U415 : NAND2_X2 port map( A1 => n4518, A2 => n4497, ZN => n3324);
   U416 : NAND2_X2 port map( A1 => n4492, A2 => ADD_RD2(6), ZN => n3349);
   U417 : NAND2_X2 port map( A1 => n4508, A2 => n4489, ZN => n3311);
   U418 : NAND2_X2 port map( A1 => n4520, A2 => n4495, ZN => n3334);
   U419 : NAND2_X2 port map( A1 => n3203, A2 => n1750, ZN => n2003);
   U420 : NAND2_X2 port map( A1 => n3224, A2 => n3211, ZN => n1994);
   U421 : NAND2_X2 port map( A1 => n1927, A2 => n1781, ZN => n1933);
   U422 : NAND2_X2 port map( A1 => n3203, A2 => n3204, ZN => n1965);
   U423 : NAND2_X2 port map( A1 => n4490, A2 => n4489, ZN => n3288);
   U424 : NAND2_X2 port map( A1 => n3224, A2 => n3212, ZN => n1993);
   U425 : AND2_X2 port map( A1 => n3203, A2 => n1757, ZN => n1996);
   U426 : NOR3_X2 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(5), A3 => n3227, ZN
                           => n3203);
   U427 : AND2_X2 port map( A1 => n3236, A2 => n3208, ZN => n2014);
   U428 : NOR3_X2 port map( A1 => n3215, A2 => ADD_RD1(4), A3 => n3238, ZN => 
                           n3236);
   U429 : AND2_X2 port map( A1 => n4530, A2 => n4491, ZN => n3353);
   U430 : NAND2_X2 port map( A1 => n3206, A2 => n3207, ZN => n1963);
   U431 : NAND2_X2 port map( A1 => n3223, A2 => n3211, ZN => n2027);
   U432 : NAND2_X2 port map( A1 => n3234, A2 => n1755, ZN => n2017);
   U433 : NAND2_X2 port map( A1 => n1750, A2 => ADD_RD1(6), ZN => n2041);
   U434 : NAND2_X2 port map( A1 => n4508, A2 => n4497, ZN => n3307);
   U435 : NAND2_X2 port map( A1 => n4507, A2 => n4496, ZN => n3341);
   U436 : NAND2_X2 port map( A1 => n4520, A2 => n4492, ZN => n3330);
   U437 : NAND2_X2 port map( A1 => n4518, A2 => n4493, ZN => n3366);
   U438 : NAND2_X2 port map( A1 => n4495, A2 => ADD_RD2(6), ZN => n3356);
   U439 : NAND2_X2 port map( A1 => n4490, A2 => n4488, ZN => n3283);
   U440 : NOR3_X2 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), A3 => n4499, ZN
                           => n4490);
   U441 : NAND2_X2 port map( A1 => n1927, A2 => n1784, ZN => n1935);
   U442 : NAND4_X2 port map( A1 => n3252, A2 => n3253, A3 => n3254, A4 => n3255
                           , ZN => n1948);
   U443 : NAND2_X2 port map( A1 => n4490, A2 => n4491, ZN => n3278);
   U444 : NAND2_X2 port map( A1 => n3234, A2 => n3207, ZN => n2051);
   U445 : NAND2_X2 port map( A1 => n3203, A2 => n1755, ZN => n1964);
   U446 : NAND2_X2 port map( A1 => n3223, A2 => n1750, ZN => n1989);
   U447 : NOR3_X2 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n3238, ZN
                           => n3223);
   U448 : NAND2_X2 port map( A1 => n3234, A2 => n3211, ZN => n2012);
   U449 : NOR3_X2 port map( A1 => n3227, A2 => ADD_RD1(3), A3 => n3238, ZN => 
                           n3234);
   U450 : NAND2_X2 port map( A1 => n1757, A2 => ADD_RD1(6), ZN => n2036);
   U451 : NAND2_X2 port map( A1 => n4487, A2 => n4489, ZN => n3279);
   U452 : NAND2_X2 port map( A1 => n4507, A2 => n4495, ZN => n3301);
   U453 : NOR3_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n4522, ZN
                           => n4507);
   U454 : NAND2_X2 port map( A1 => n4518, A2 => n4496, ZN => n3325);
   U455 : NOR3_X2 port map( A1 => n4511, A2 => ADD_RD2(3), A3 => n4522, ZN => 
                           n4518);
   U456 : NAND2_X2 port map( A1 => n4493, A2 => ADD_RD2(6), ZN => n3350);
   U457 : NAND2_X2 port map( A1 => n3224, A2 => n3204, ZN => n1999);
   U458 : NOR3_X2 port map( A1 => n3215, A2 => ADD_RD1(5), A3 => n3227, ZN => 
                           n3224);
   U459 : NAND2_X2 port map( A1 => n3236, A2 => n3212, ZN => n2022);
   U460 : NAND2_X2 port map( A1 => n3246, A2 => n3208, ZN => n2045);
   U461 : NAND2_X2 port map( A1 => n4508, A2 => n4488, ZN => n3312);
   U462 : NOR3_X2 port map( A1 => n4499, A2 => ADD_RD2(5), A3 => n4511, ZN => 
                           n4508);
   U463 : NAND2_X2 port map( A1 => n4520, A2 => n4497, ZN => n3335);
   U464 : NOR3_X2 port map( A1 => n4499, A2 => ADD_RD2(4), A3 => n4522, ZN => 
                           n4520);
   U465 : NAND2_X2 port map( A1 => n4530, A2 => n4492, ZN => n3361);
   U466 : NAND2_X2 port map( A1 => n1927, A2 => n1793, ZN => n1945);
   U467 : NAND4_X2 port map( A1 => n4536, A2 => n4537, A3 => n4538, A4 => n4539
                           , ZN => n3263);
   U468 : OAI22_X1 port map( A1 => n1758, A2 => n1759, B1 => n1722, B2 => n618,
                           ZN => n9977);
   U469 : OAI22_X1 port map( A1 => n1758, A2 => n1761, B1 => n1722, B2 => n621,
                           ZN => n9976);
   U470 : OAI22_X1 port map( A1 => n1758, A2 => n1762, B1 => n1722, B2 => n624,
                           ZN => n9975);
   U471 : OAI22_X1 port map( A1 => n1758, A2 => n1763, B1 => n1722, B2 => n627,
                           ZN => n9974);
   U472 : OAI22_X1 port map( A1 => n1758, A2 => n1764, B1 => n1722, B2 => n630,
                           ZN => n9973);
   U473 : OAI22_X1 port map( A1 => n1758, A2 => n1765, B1 => n1722, B2 => n633,
                           ZN => n9972);
   U474 : OAI22_X1 port map( A1 => n1758, A2 => n1766, B1 => n1722, B2 => n636,
                           ZN => n9971);
   U475 : OAI22_X1 port map( A1 => n1758, A2 => n1767, B1 => n1722, B2 => n639,
                           ZN => n9970);
   U476 : OAI22_X1 port map( A1 => n1758, A2 => n1746, B1 => n1722, B2 => n642,
                           ZN => n9969);
   U477 : OAI22_X1 port map( A1 => n1758, A2 => n1747, B1 => n1722, B2 => n645,
                           ZN => n9968);
   U478 : OAI22_X1 port map( A1 => n1758, A2 => n1742, B1 => n1722, B2 => n648,
                           ZN => n9967);
   U479 : OAI22_X1 port map( A1 => n1758, A2 => n1743, B1 => n1722, B2 => n651,
                           ZN => n9966);
   U480 : OAI22_X1 port map( A1 => n1758, A2 => n1744, B1 => n1722, B2 => n654,
                           ZN => n9965);
   U481 : OAI22_X1 port map( A1 => n1758, A2 => n1745, B1 => n1722, B2 => n657,
                           ZN => n9964);
   U482 : OAI22_X1 port map( A1 => n1758, A2 => n1738, B1 => n1722, B2 => n660,
                           ZN => n9963);
   U483 : OAI22_X1 port map( A1 => n1758, A2 => n1739, B1 => n1722, B2 => n663,
                           ZN => n9962);
   U484 : OAI22_X1 port map( A1 => n1758, A2 => n1740, B1 => n1722, B2 => n666,
                           ZN => n9961);
   U485 : OAI22_X1 port map( A1 => n1758, A2 => n1741, B1 => n1722, B2 => n669,
                           ZN => n9960);
   U486 : OAI22_X1 port map( A1 => n1758, A2 => n1734, B1 => n1722, B2 => n672,
                           ZN => n9959);
   U487 : OAI22_X1 port map( A1 => n1758, A2 => n1735, B1 => n1722, B2 => n675,
                           ZN => n9958);
   U488 : OAI22_X1 port map( A1 => n1758, A2 => n1736, B1 => n1722, B2 => n678,
                           ZN => n9957);
   U489 : OAI22_X1 port map( A1 => n1758, A2 => n1737, B1 => n1722, B2 => n681,
                           ZN => n9956);
   U490 : OAI22_X1 port map( A1 => n1758, A2 => n1730, B1 => n1722, B2 => n684,
                           ZN => n9955);
   U491 : OAI22_X1 port map( A1 => n1758, A2 => n1731, B1 => n1722, B2 => n687,
                           ZN => n9954);
   U492 : OAI22_X1 port map( A1 => n1758, A2 => n1732, B1 => n1722, B2 => n690,
                           ZN => n9953);
   U493 : OAI22_X1 port map( A1 => n1758, A2 => n1733, B1 => n1722, B2 => n693,
                           ZN => n9952);
   U494 : OAI22_X1 port map( A1 => n1758, A2 => n1726, B1 => n1722, B2 => n696,
                           ZN => n9951);
   U495 : OAI22_X1 port map( A1 => n1758, A2 => n1727, B1 => n1722, B2 => n699,
                           ZN => n9950);
   U496 : OAI22_X1 port map( A1 => n1758, A2 => n1728, B1 => n1722, B2 => n702,
                           ZN => n9949);
   U497 : OAI22_X1 port map( A1 => n1758, A2 => n1729, B1 => n1722, B2 => n705,
                           ZN => n9948);
   U498 : OAI22_X1 port map( A1 => n1758, A2 => n1725, B1 => n1722, B2 => n708,
                           ZN => n9947);
   U499 : OAI22_X1 port map( A1 => n1758, A2 => n1768, B1 => n1722, B2 => n711,
                           ZN => n9946);
   U500 : OAI21_X1 port map( B1 => n1758, B2 => n1769, A => n1770, ZN => n1760)
                           ;
   U501 : OAI22_X1 port map( A1 => n1759, A2 => n1773, B1 => n1724, B2 => n194,
                           ZN => n9945);
   U502 : OAI22_X1 port map( A1 => n1761, A2 => n1773, B1 => n1724, B2 => n197,
                           ZN => n9944);
   U503 : OAI22_X1 port map( A1 => n1762, A2 => n1773, B1 => n1724, B2 => n200,
                           ZN => n9943);
   U504 : OAI22_X1 port map( A1 => n1763, A2 => n1773, B1 => n1724, B2 => n203,
                           ZN => n9942);
   U505 : OAI22_X1 port map( A1 => n1764, A2 => n1773, B1 => n1724, B2 => n206,
                           ZN => n9941);
   U506 : OAI22_X1 port map( A1 => n1765, A2 => n1773, B1 => n1724, B2 => n209,
                           ZN => n9940);
   U507 : OAI22_X1 port map( A1 => n1766, A2 => n1773, B1 => n1724, B2 => n212,
                           ZN => n9939);
   U508 : OAI22_X1 port map( A1 => n1767, A2 => n1773, B1 => n1724, B2 => n215,
                           ZN => n9938);
   U509 : OAI22_X1 port map( A1 => n1746, A2 => n1773, B1 => n1724, B2 => n218,
                           ZN => n9937);
   U510 : OAI22_X1 port map( A1 => n1747, A2 => n1773, B1 => n1724, B2 => n221,
                           ZN => n9936);
   U511 : OAI22_X1 port map( A1 => n1742, A2 => n1773, B1 => n1724, B2 => n224,
                           ZN => n9935);
   U512 : OAI22_X1 port map( A1 => n1743, A2 => n1773, B1 => n1724, B2 => n227,
                           ZN => n9934);
   U513 : OAI22_X1 port map( A1 => n1744, A2 => n1773, B1 => n1724, B2 => n230,
                           ZN => n9933);
   U514 : OAI22_X1 port map( A1 => n1745, A2 => n1773, B1 => n1724, B2 => n233,
                           ZN => n9932);
   U515 : OAI22_X1 port map( A1 => n1738, A2 => n1773, B1 => n1724, B2 => n236,
                           ZN => n9931);
   U516 : OAI22_X1 port map( A1 => n1739, A2 => n1773, B1 => n1724, B2 => n239,
                           ZN => n9930);
   U517 : OAI22_X1 port map( A1 => n1740, A2 => n1773, B1 => n1724, B2 => n242,
                           ZN => n9929);
   U518 : OAI22_X1 port map( A1 => n1741, A2 => n1773, B1 => n1724, B2 => n245,
                           ZN => n9928);
   U519 : OAI22_X1 port map( A1 => n1734, A2 => n1773, B1 => n1724, B2 => n248,
                           ZN => n9927);
   U520 : OAI22_X1 port map( A1 => n1735, A2 => n1773, B1 => n1724, B2 => n251,
                           ZN => n9926);
   U521 : OAI22_X1 port map( A1 => n1736, A2 => n1773, B1 => n1724, B2 => n254,
                           ZN => n9925);
   U522 : OAI22_X1 port map( A1 => n1737, A2 => n1773, B1 => n1724, B2 => n257,
                           ZN => n9924);
   U523 : OAI22_X1 port map( A1 => n1730, A2 => n1773, B1 => n1724, B2 => n260,
                           ZN => n9923);
   U524 : OAI22_X1 port map( A1 => n1731, A2 => n1773, B1 => n1724, B2 => n263,
                           ZN => n9922);
   U525 : OAI22_X1 port map( A1 => n1732, A2 => n1773, B1 => n1724, B2 => n266,
                           ZN => n9921);
   U526 : OAI22_X1 port map( A1 => n1733, A2 => n1773, B1 => n1724, B2 => n269,
                           ZN => n9920);
   U527 : OAI22_X1 port map( A1 => n1726, A2 => n1773, B1 => n1724, B2 => n272,
                           ZN => n9919);
   U528 : OAI22_X1 port map( A1 => n1727, A2 => n1773, B1 => n1724, B2 => n275,
                           ZN => n9918);
   U529 : OAI22_X1 port map( A1 => n1728, A2 => n1773, B1 => n1724, B2 => n278,
                           ZN => n9917);
   U530 : OAI22_X1 port map( A1 => n1729, A2 => n1773, B1 => n1724, B2 => n281,
                           ZN => n9916);
   U531 : OAI22_X1 port map( A1 => n1725, A2 => n1773, B1 => n1724, B2 => n284,
                           ZN => n9915);
   U532 : OAI22_X1 port map( A1 => n1768, A2 => n1773, B1 => n1724, B2 => n287,
                           ZN => n9914);
   U533 : OAI21_X1 port map( B1 => n1769, B2 => n1773, A => n1770, ZN => n1774)
                           ;
   U534 : OAI22_X1 port map( A1 => n1759, A2 => n1776, B1 => n5696, B2 => n1658
                           , ZN => n9913);
   U535 : OAI22_X1 port map( A1 => n1761, A2 => n1776, B1 => n5686, B2 => n1658
                           , ZN => n9912);
   U536 : OAI22_X1 port map( A1 => n1762, A2 => n1776, B1 => n5676, B2 => n1658
                           , ZN => n9911);
   U537 : OAI22_X1 port map( A1 => n1763, A2 => n1776, B1 => n5666, B2 => n1658
                           , ZN => n9910);
   U538 : OAI22_X1 port map( A1 => n1764, A2 => n1776, B1 => n5656, B2 => n1658
                           , ZN => n9909);
   U539 : OAI22_X1 port map( A1 => n1765, A2 => n1776, B1 => n5646, B2 => n1658
                           , ZN => n9908);
   U540 : OAI22_X1 port map( A1 => n1766, A2 => n1776, B1 => n5636, B2 => n1658
                           , ZN => n9907);
   U541 : OAI22_X1 port map( A1 => n1767, A2 => n1776, B1 => n5626, B2 => n1658
                           , ZN => n9906);
   U542 : OAI22_X1 port map( A1 => n1746, A2 => n1776, B1 => n5616, B2 => n1658
                           , ZN => n9905);
   U543 : OAI22_X1 port map( A1 => n1747, A2 => n1776, B1 => n5606, B2 => n1658
                           , ZN => n9904);
   U544 : OAI22_X1 port map( A1 => n1742, A2 => n1776, B1 => n5596, B2 => n1658
                           , ZN => n9903);
   U545 : OAI22_X1 port map( A1 => n1743, A2 => n1776, B1 => n5586, B2 => n1658
                           , ZN => n9902);
   U546 : OAI22_X1 port map( A1 => n1744, A2 => n1776, B1 => n5576, B2 => n1658
                           , ZN => n9901);
   U547 : OAI22_X1 port map( A1 => n1745, A2 => n1776, B1 => n5566, B2 => n1658
                           , ZN => n9900);
   U548 : OAI22_X1 port map( A1 => n1738, A2 => n1776, B1 => n5556, B2 => n1658
                           , ZN => n9899);
   U549 : OAI22_X1 port map( A1 => n1739, A2 => n1776, B1 => n5546, B2 => n1658
                           , ZN => n9898);
   U550 : OAI22_X1 port map( A1 => n1740, A2 => n1776, B1 => n5536, B2 => n1658
                           , ZN => n9897);
   U551 : OAI22_X1 port map( A1 => n1741, A2 => n1776, B1 => n5526, B2 => n1658
                           , ZN => n9896);
   U552 : OAI22_X1 port map( A1 => n1734, A2 => n1776, B1 => n5516, B2 => n1658
                           , ZN => n9895);
   U553 : OAI22_X1 port map( A1 => n1735, A2 => n1776, B1 => n5506, B2 => n1658
                           , ZN => n9894);
   U554 : OAI22_X1 port map( A1 => n1736, A2 => n1776, B1 => n5496, B2 => n1658
                           , ZN => n9893);
   U555 : OAI22_X1 port map( A1 => n1737, A2 => n1776, B1 => n5486, B2 => n1658
                           , ZN => n9892);
   U556 : OAI22_X1 port map( A1 => n1730, A2 => n1776, B1 => n5476, B2 => n1658
                           , ZN => n9891);
   U557 : OAI22_X1 port map( A1 => n1731, A2 => n1776, B1 => n5466, B2 => n1658
                           , ZN => n9890);
   U558 : OAI22_X1 port map( A1 => n1732, A2 => n1776, B1 => n5456, B2 => n1658
                           , ZN => n9889);
   U559 : OAI22_X1 port map( A1 => n1733, A2 => n1776, B1 => n5446, B2 => n1658
                           , ZN => n9888);
   U560 : OAI22_X1 port map( A1 => n1726, A2 => n1776, B1 => n5436, B2 => n1658
                           , ZN => n9887);
   U561 : OAI22_X1 port map( A1 => n1727, A2 => n1776, B1 => n5426, B2 => n1658
                           , ZN => n9886);
   U562 : OAI22_X1 port map( A1 => n1728, A2 => n1776, B1 => n5416, B2 => n1658
                           , ZN => n9885);
   U563 : OAI22_X1 port map( A1 => n1729, A2 => n1776, B1 => n5406, B2 => n1658
                           , ZN => n9884);
   U564 : OAI22_X1 port map( A1 => n1725, A2 => n1776, B1 => n5396, B2 => n1658
                           , ZN => n9883);
   U565 : OAI22_X1 port map( A1 => n1768, A2 => n1776, B1 => n5386, B2 => n1658
                           , ZN => n9882);
   U566 : OAI21_X1 port map( B1 => n1769, B2 => n1776, A => n1770, ZN => n1777)
                           ;
   U567 : OAI22_X1 port map( A1 => n1759, A2 => n1779, B1 => n5697, B2 => n1660
                           , ZN => n9881);
   U568 : OAI22_X1 port map( A1 => n1761, A2 => n1779, B1 => n5687, B2 => n1660
                           , ZN => n9880);
   U569 : OAI22_X1 port map( A1 => n1762, A2 => n1779, B1 => n5677, B2 => n1660
                           , ZN => n9879);
   U570 : OAI22_X1 port map( A1 => n1763, A2 => n1779, B1 => n5667, B2 => n1660
                           , ZN => n9878);
   U571 : OAI22_X1 port map( A1 => n1764, A2 => n1779, B1 => n5657, B2 => n1660
                           , ZN => n9877);
   U572 : OAI22_X1 port map( A1 => n1765, A2 => n1779, B1 => n5647, B2 => n1660
                           , ZN => n9876);
   U573 : OAI22_X1 port map( A1 => n1766, A2 => n1779, B1 => n5637, B2 => n1660
                           , ZN => n9875);
   U574 : OAI22_X1 port map( A1 => n1767, A2 => n1779, B1 => n5627, B2 => n1660
                           , ZN => n9874);
   U575 : OAI22_X1 port map( A1 => n1746, A2 => n1779, B1 => n5617, B2 => n1660
                           , ZN => n9873);
   U576 : OAI22_X1 port map( A1 => n1747, A2 => n1779, B1 => n5607, B2 => n1660
                           , ZN => n9872);
   U577 : OAI22_X1 port map( A1 => n1742, A2 => n1779, B1 => n5597, B2 => n1660
                           , ZN => n9871);
   U578 : OAI22_X1 port map( A1 => n1743, A2 => n1779, B1 => n5587, B2 => n1660
                           , ZN => n9870);
   U579 : OAI22_X1 port map( A1 => n1744, A2 => n1779, B1 => n5577, B2 => n1660
                           , ZN => n9869);
   U580 : OAI22_X1 port map( A1 => n1745, A2 => n1779, B1 => n5567, B2 => n1660
                           , ZN => n9868);
   U581 : OAI22_X1 port map( A1 => n1738, A2 => n1779, B1 => n5557, B2 => n1660
                           , ZN => n9867);
   U582 : OAI22_X1 port map( A1 => n1739, A2 => n1779, B1 => n5547, B2 => n1660
                           , ZN => n9866);
   U583 : OAI22_X1 port map( A1 => n1740, A2 => n1779, B1 => n5537, B2 => n1660
                           , ZN => n9865);
   U584 : OAI22_X1 port map( A1 => n1741, A2 => n1779, B1 => n5527, B2 => n1660
                           , ZN => n9864);
   U585 : OAI22_X1 port map( A1 => n1734, A2 => n1779, B1 => n5517, B2 => n1660
                           , ZN => n9863);
   U586 : OAI22_X1 port map( A1 => n1735, A2 => n1779, B1 => n5507, B2 => n1660
                           , ZN => n9862);
   U587 : OAI22_X1 port map( A1 => n1736, A2 => n1779, B1 => n5497, B2 => n1660
                           , ZN => n9861);
   U588 : OAI22_X1 port map( A1 => n1737, A2 => n1779, B1 => n5487, B2 => n1660
                           , ZN => n9860);
   U589 : OAI22_X1 port map( A1 => n1730, A2 => n1779, B1 => n5477, B2 => n1660
                           , ZN => n9859);
   U590 : OAI22_X1 port map( A1 => n1731, A2 => n1779, B1 => n5467, B2 => n1660
                           , ZN => n9858);
   U591 : OAI22_X1 port map( A1 => n1732, A2 => n1779, B1 => n5457, B2 => n1660
                           , ZN => n9857);
   U592 : OAI22_X1 port map( A1 => n1733, A2 => n1779, B1 => n5447, B2 => n1660
                           , ZN => n9856);
   U593 : OAI22_X1 port map( A1 => n1726, A2 => n1779, B1 => n5437, B2 => n1660
                           , ZN => n9855);
   U594 : OAI22_X1 port map( A1 => n1727, A2 => n1779, B1 => n5427, B2 => n1660
                           , ZN => n9854);
   U595 : OAI22_X1 port map( A1 => n1728, A2 => n1779, B1 => n5417, B2 => n1660
                           , ZN => n9853);
   U596 : OAI22_X1 port map( A1 => n1729, A2 => n1779, B1 => n5407, B2 => n1660
                           , ZN => n9852);
   U597 : OAI22_X1 port map( A1 => n1725, A2 => n1779, B1 => n5397, B2 => n1660
                           , ZN => n9851);
   U598 : OAI22_X1 port map( A1 => n1768, A2 => n1779, B1 => n5387, B2 => n1660
                           , ZN => n9850);
   U599 : OAI21_X1 port map( B1 => n1769, B2 => n1779, A => n1770, ZN => n1780)
                           ;
   U600 : OAI22_X1 port map( A1 => n1759, A2 => n1782, B1 => n1718, B2 => n809,
                           ZN => n9849);
   U601 : OAI22_X1 port map( A1 => n1761, A2 => n1782, B1 => n1718, B2 => n810,
                           ZN => n9848);
   U602 : OAI22_X1 port map( A1 => n1762, A2 => n1782, B1 => n1718, B2 => n811,
                           ZN => n9847);
   U603 : OAI22_X1 port map( A1 => n1763, A2 => n1782, B1 => n1718, B2 => n812,
                           ZN => n9846);
   U604 : OAI22_X1 port map( A1 => n1764, A2 => n1782, B1 => n1718, B2 => n813,
                           ZN => n9845);
   U605 : OAI22_X1 port map( A1 => n1765, A2 => n1782, B1 => n1718, B2 => n814,
                           ZN => n9844);
   U606 : OAI22_X1 port map( A1 => n1766, A2 => n1782, B1 => n1718, B2 => n815,
                           ZN => n9843);
   U607 : OAI22_X1 port map( A1 => n1767, A2 => n1782, B1 => n1718, B2 => n816,
                           ZN => n9842);
   U608 : OAI22_X1 port map( A1 => n1746, A2 => n1782, B1 => n1718, B2 => n817,
                           ZN => n9841);
   U609 : OAI22_X1 port map( A1 => n1747, A2 => n1782, B1 => n1718, B2 => n818,
                           ZN => n9840);
   U610 : OAI22_X1 port map( A1 => n1742, A2 => n1782, B1 => n1718, B2 => n819,
                           ZN => n9839);
   U611 : OAI22_X1 port map( A1 => n1743, A2 => n1782, B1 => n1718, B2 => n820,
                           ZN => n9838);
   U612 : OAI22_X1 port map( A1 => n1744, A2 => n1782, B1 => n1718, B2 => n821,
                           ZN => n9837);
   U613 : OAI22_X1 port map( A1 => n1745, A2 => n1782, B1 => n1718, B2 => n822,
                           ZN => n9836);
   U614 : OAI22_X1 port map( A1 => n1738, A2 => n1782, B1 => n1718, B2 => n823,
                           ZN => n9835);
   U615 : OAI22_X1 port map( A1 => n1739, A2 => n1782, B1 => n1718, B2 => n824,
                           ZN => n9834);
   U616 : OAI22_X1 port map( A1 => n1740, A2 => n1782, B1 => n1718, B2 => n825,
                           ZN => n9833);
   U617 : OAI22_X1 port map( A1 => n1741, A2 => n1782, B1 => n1718, B2 => n826,
                           ZN => n9832);
   U618 : OAI22_X1 port map( A1 => n1734, A2 => n1782, B1 => n1718, B2 => n827,
                           ZN => n9831);
   U619 : OAI22_X1 port map( A1 => n1735, A2 => n1782, B1 => n1718, B2 => n828,
                           ZN => n9830);
   U620 : OAI22_X1 port map( A1 => n1736, A2 => n1782, B1 => n1718, B2 => n829,
                           ZN => n9829);
   U621 : OAI22_X1 port map( A1 => n1737, A2 => n1782, B1 => n1718, B2 => n830,
                           ZN => n9828);
   U622 : OAI22_X1 port map( A1 => n1730, A2 => n1782, B1 => n1718, B2 => n831,
                           ZN => n9827);
   U623 : OAI22_X1 port map( A1 => n1731, A2 => n1782, B1 => n1718, B2 => n832,
                           ZN => n9826);
   U624 : OAI22_X1 port map( A1 => n1732, A2 => n1782, B1 => n1718, B2 => n833,
                           ZN => n9825);
   U625 : OAI22_X1 port map( A1 => n1733, A2 => n1782, B1 => n1718, B2 => n834,
                           ZN => n9824);
   U626 : OAI22_X1 port map( A1 => n1726, A2 => n1782, B1 => n1718, B2 => n835,
                           ZN => n9823);
   U627 : OAI22_X1 port map( A1 => n1727, A2 => n1782, B1 => n1718, B2 => n836,
                           ZN => n9822);
   U628 : OAI22_X1 port map( A1 => n1728, A2 => n1782, B1 => n1718, B2 => n837,
                           ZN => n9821);
   U629 : OAI22_X1 port map( A1 => n1729, A2 => n1782, B1 => n1718, B2 => n838,
                           ZN => n9820);
   U630 : OAI22_X1 port map( A1 => n1725, A2 => n1782, B1 => n1718, B2 => n839,
                           ZN => n9819);
   U631 : OAI22_X1 port map( A1 => n1768, A2 => n1782, B1 => n1718, B2 => n840,
                           ZN => n9818);
   U632 : OAI21_X1 port map( B1 => n1769, B2 => n1782, A => n1770, ZN => n1783)
                           ;
   U633 : OAI22_X1 port map( A1 => n1759, A2 => n1785, B1 => n1720, B2 => n1161
                           , ZN => n9817);
   U634 : OAI22_X1 port map( A1 => n1761, A2 => n1785, B1 => n1720, B2 => n1162
                           , ZN => n9816);
   U635 : OAI22_X1 port map( A1 => n1762, A2 => n1785, B1 => n1720, B2 => n1163
                           , ZN => n9815);
   U636 : OAI22_X1 port map( A1 => n1763, A2 => n1785, B1 => n1720, B2 => n1164
                           , ZN => n9814);
   U637 : OAI22_X1 port map( A1 => n1764, A2 => n1785, B1 => n1720, B2 => n1165
                           , ZN => n9813);
   U638 : OAI22_X1 port map( A1 => n1765, A2 => n1785, B1 => n1720, B2 => n1166
                           , ZN => n9812);
   U639 : OAI22_X1 port map( A1 => n1766, A2 => n1785, B1 => n1720, B2 => n1167
                           , ZN => n9811);
   U640 : OAI22_X1 port map( A1 => n1767, A2 => n1785, B1 => n1720, B2 => n1168
                           , ZN => n9810);
   U641 : OAI22_X1 port map( A1 => n1746, A2 => n1785, B1 => n1720, B2 => n1169
                           , ZN => n9809);
   U642 : OAI22_X1 port map( A1 => n1747, A2 => n1785, B1 => n1720, B2 => n1170
                           , ZN => n9808);
   U643 : OAI22_X1 port map( A1 => n1742, A2 => n1785, B1 => n1720, B2 => n1171
                           , ZN => n9807);
   U644 : OAI22_X1 port map( A1 => n1743, A2 => n1785, B1 => n1720, B2 => n1172
                           , ZN => n9806);
   U645 : OAI22_X1 port map( A1 => n1744, A2 => n1785, B1 => n1720, B2 => n1173
                           , ZN => n9805);
   U646 : OAI22_X1 port map( A1 => n1745, A2 => n1785, B1 => n1720, B2 => n1174
                           , ZN => n9804);
   U647 : OAI22_X1 port map( A1 => n1738, A2 => n1785, B1 => n1720, B2 => n1175
                           , ZN => n9803);
   U648 : OAI22_X1 port map( A1 => n1739, A2 => n1785, B1 => n1720, B2 => n1176
                           , ZN => n9802);
   U649 : OAI22_X1 port map( A1 => n1740, A2 => n1785, B1 => n1720, B2 => n1177
                           , ZN => n9801);
   U650 : OAI22_X1 port map( A1 => n1741, A2 => n1785, B1 => n1720, B2 => n1178
                           , ZN => n9800);
   U651 : OAI22_X1 port map( A1 => n1734, A2 => n1785, B1 => n1720, B2 => n1179
                           , ZN => n9799);
   U652 : OAI22_X1 port map( A1 => n1735, A2 => n1785, B1 => n1720, B2 => n1180
                           , ZN => n9798);
   U653 : OAI22_X1 port map( A1 => n1736, A2 => n1785, B1 => n1720, B2 => n1181
                           , ZN => n9797);
   U654 : OAI22_X1 port map( A1 => n1737, A2 => n1785, B1 => n1720, B2 => n1182
                           , ZN => n9796);
   U655 : OAI22_X1 port map( A1 => n1730, A2 => n1785, B1 => n1720, B2 => n1183
                           , ZN => n9795);
   U656 : OAI22_X1 port map( A1 => n1731, A2 => n1785, B1 => n1720, B2 => n1184
                           , ZN => n9794);
   U657 : OAI22_X1 port map( A1 => n1732, A2 => n1785, B1 => n1720, B2 => n1185
                           , ZN => n9793);
   U658 : OAI22_X1 port map( A1 => n1733, A2 => n1785, B1 => n1720, B2 => n1186
                           , ZN => n9792);
   U659 : OAI22_X1 port map( A1 => n1726, A2 => n1785, B1 => n1720, B2 => n1187
                           , ZN => n9791);
   U660 : OAI22_X1 port map( A1 => n1727, A2 => n1785, B1 => n1720, B2 => n1188
                           , ZN => n9790);
   U661 : OAI22_X1 port map( A1 => n1728, A2 => n1785, B1 => n1720, B2 => n1189
                           , ZN => n9789);
   U662 : OAI22_X1 port map( A1 => n1729, A2 => n1785, B1 => n1720, B2 => n1190
                           , ZN => n9788);
   U663 : OAI22_X1 port map( A1 => n1725, A2 => n1785, B1 => n1720, B2 => n1191
                           , ZN => n9787);
   U664 : OAI22_X1 port map( A1 => n1768, A2 => n1785, B1 => n1720, B2 => n1192
                           , ZN => n9786);
   U665 : OAI21_X1 port map( B1 => n1769, B2 => n1785, A => n1770, ZN => n1786)
                           ;
   U666 : OAI22_X1 port map( A1 => n1759, A2 => n1788, B1 => n5377, B2 => n1654
                           , ZN => n9785);
   U667 : OAI22_X1 port map( A1 => n1761, A2 => n1788, B1 => n5376, B2 => n1654
                           , ZN => n9784);
   U668 : OAI22_X1 port map( A1 => n1762, A2 => n1788, B1 => n5375, B2 => n1654
                           , ZN => n9783);
   U669 : OAI22_X1 port map( A1 => n1763, A2 => n1788, B1 => n5374, B2 => n1654
                           , ZN => n9782);
   U670 : OAI22_X1 port map( A1 => n1764, A2 => n1788, B1 => n5373, B2 => n1654
                           , ZN => n9781);
   U671 : OAI22_X1 port map( A1 => n1765, A2 => n1788, B1 => n5372, B2 => n1654
                           , ZN => n9780);
   U672 : OAI22_X1 port map( A1 => n1766, A2 => n1788, B1 => n5371, B2 => n1654
                           , ZN => n9779);
   U673 : OAI22_X1 port map( A1 => n1767, A2 => n1788, B1 => n5370, B2 => n1654
                           , ZN => n9778);
   U674 : OAI22_X1 port map( A1 => n1746, A2 => n1788, B1 => n5369, B2 => n1654
                           , ZN => n9777);
   U675 : OAI22_X1 port map( A1 => n1747, A2 => n1788, B1 => n5368, B2 => n1654
                           , ZN => n9776);
   U676 : OAI22_X1 port map( A1 => n1742, A2 => n1788, B1 => n5367, B2 => n1654
                           , ZN => n9775);
   U677 : OAI22_X1 port map( A1 => n1743, A2 => n1788, B1 => n5366, B2 => n1654
                           , ZN => n9774);
   U678 : OAI22_X1 port map( A1 => n1744, A2 => n1788, B1 => n5365, B2 => n1654
                           , ZN => n9773);
   U679 : OAI22_X1 port map( A1 => n1745, A2 => n1788, B1 => n5364, B2 => n1654
                           , ZN => n9772);
   U680 : OAI22_X1 port map( A1 => n1738, A2 => n1788, B1 => n5363, B2 => n1654
                           , ZN => n9771);
   U681 : OAI22_X1 port map( A1 => n1739, A2 => n1788, B1 => n5362, B2 => n1654
                           , ZN => n9770);
   U682 : OAI22_X1 port map( A1 => n1740, A2 => n1788, B1 => n5361, B2 => n1654
                           , ZN => n9769);
   U683 : OAI22_X1 port map( A1 => n1741, A2 => n1788, B1 => n5360, B2 => n1654
                           , ZN => n9768);
   U684 : OAI22_X1 port map( A1 => n1734, A2 => n1788, B1 => n5359, B2 => n1654
                           , ZN => n9767);
   U685 : OAI22_X1 port map( A1 => n1735, A2 => n1788, B1 => n5358, B2 => n1654
                           , ZN => n9766);
   U686 : OAI22_X1 port map( A1 => n1736, A2 => n1788, B1 => n5357, B2 => n1654
                           , ZN => n9765);
   U687 : OAI22_X1 port map( A1 => n1737, A2 => n1788, B1 => n5356, B2 => n1654
                           , ZN => n9764);
   U688 : OAI22_X1 port map( A1 => n1730, A2 => n1788, B1 => n5355, B2 => n1654
                           , ZN => n9763);
   U689 : OAI22_X1 port map( A1 => n1731, A2 => n1788, B1 => n5354, B2 => n1654
                           , ZN => n9762);
   U690 : OAI22_X1 port map( A1 => n1732, A2 => n1788, B1 => n5353, B2 => n1654
                           , ZN => n9761);
   U691 : OAI22_X1 port map( A1 => n1733, A2 => n1788, B1 => n5352, B2 => n1654
                           , ZN => n9760);
   U692 : OAI22_X1 port map( A1 => n1726, A2 => n1788, B1 => n5351, B2 => n1654
                           , ZN => n9759);
   U693 : OAI22_X1 port map( A1 => n1727, A2 => n1788, B1 => n5350, B2 => n1654
                           , ZN => n9758);
   U694 : OAI22_X1 port map( A1 => n1728, A2 => n1788, B1 => n5349, B2 => n1654
                           , ZN => n9757);
   U695 : OAI22_X1 port map( A1 => n1729, A2 => n1788, B1 => n5348, B2 => n1654
                           , ZN => n9756);
   U696 : OAI22_X1 port map( A1 => n1725, A2 => n1788, B1 => n5347, B2 => n1654
                           , ZN => n9755);
   U697 : OAI22_X1 port map( A1 => n1768, A2 => n1788, B1 => n5346, B2 => n1654
                           , ZN => n9754);
   U698 : OAI21_X1 port map( B1 => n1769, B2 => n1788, A => n1770, ZN => n1789)
                           ;
   U699 : OAI22_X1 port map( A1 => n1759, A2 => n1791, B1 => n5345, B2 => n1656
                           , ZN => n9753);
   U700 : OAI22_X1 port map( A1 => n1761, A2 => n1791, B1 => n5344, B2 => n1656
                           , ZN => n9752);
   U701 : OAI22_X1 port map( A1 => n1762, A2 => n1791, B1 => n5343, B2 => n1656
                           , ZN => n9751);
   U702 : OAI22_X1 port map( A1 => n1763, A2 => n1791, B1 => n5342, B2 => n1656
                           , ZN => n9750);
   U703 : OAI22_X1 port map( A1 => n1764, A2 => n1791, B1 => n5341, B2 => n1656
                           , ZN => n9749);
   U704 : OAI22_X1 port map( A1 => n1765, A2 => n1791, B1 => n5340, B2 => n1656
                           , ZN => n9748);
   U705 : OAI22_X1 port map( A1 => n1766, A2 => n1791, B1 => n5339, B2 => n1656
                           , ZN => n9747);
   U706 : OAI22_X1 port map( A1 => n1767, A2 => n1791, B1 => n5338, B2 => n1656
                           , ZN => n9746);
   U707 : OAI22_X1 port map( A1 => n1746, A2 => n1791, B1 => n5337, B2 => n1656
                           , ZN => n9745);
   U708 : OAI22_X1 port map( A1 => n1747, A2 => n1791, B1 => n5336, B2 => n1656
                           , ZN => n9744);
   U709 : OAI22_X1 port map( A1 => n1742, A2 => n1791, B1 => n5335, B2 => n1656
                           , ZN => n9743);
   U710 : OAI22_X1 port map( A1 => n1743, A2 => n1791, B1 => n5334, B2 => n1656
                           , ZN => n9742);
   U711 : OAI22_X1 port map( A1 => n1744, A2 => n1791, B1 => n5333, B2 => n1656
                           , ZN => n9741);
   U712 : OAI22_X1 port map( A1 => n1745, A2 => n1791, B1 => n5332, B2 => n1656
                           , ZN => n9740);
   U713 : OAI22_X1 port map( A1 => n1738, A2 => n1791, B1 => n5331, B2 => n1656
                           , ZN => n9739);
   U714 : OAI22_X1 port map( A1 => n1739, A2 => n1791, B1 => n5330, B2 => n1656
                           , ZN => n9738);
   U715 : OAI22_X1 port map( A1 => n1740, A2 => n1791, B1 => n5329, B2 => n1656
                           , ZN => n9737);
   U716 : OAI22_X1 port map( A1 => n1741, A2 => n1791, B1 => n5328, B2 => n1656
                           , ZN => n9736);
   U717 : OAI22_X1 port map( A1 => n1734, A2 => n1791, B1 => n5327, B2 => n1656
                           , ZN => n9735);
   U718 : OAI22_X1 port map( A1 => n1735, A2 => n1791, B1 => n5326, B2 => n1656
                           , ZN => n9734);
   U719 : OAI22_X1 port map( A1 => n1736, A2 => n1791, B1 => n5325, B2 => n1656
                           , ZN => n9733);
   U720 : OAI22_X1 port map( A1 => n1737, A2 => n1791, B1 => n5324, B2 => n1656
                           , ZN => n9732);
   U721 : OAI22_X1 port map( A1 => n1730, A2 => n1791, B1 => n5323, B2 => n1656
                           , ZN => n9731);
   U722 : OAI22_X1 port map( A1 => n1731, A2 => n1791, B1 => n5322, B2 => n1656
                           , ZN => n9730);
   U723 : OAI22_X1 port map( A1 => n1732, A2 => n1791, B1 => n5321, B2 => n1656
                           , ZN => n9729);
   U724 : OAI22_X1 port map( A1 => n1733, A2 => n1791, B1 => n5320, B2 => n1656
                           , ZN => n9728);
   U725 : OAI22_X1 port map( A1 => n1726, A2 => n1791, B1 => n5319, B2 => n1656
                           , ZN => n9727);
   U726 : OAI22_X1 port map( A1 => n1727, A2 => n1791, B1 => n5318, B2 => n1656
                           , ZN => n9726);
   U727 : OAI22_X1 port map( A1 => n1728, A2 => n1791, B1 => n5317, B2 => n1656
                           , ZN => n9725);
   U728 : OAI22_X1 port map( A1 => n1729, A2 => n1791, B1 => n5316, B2 => n1656
                           , ZN => n9724);
   U729 : OAI22_X1 port map( A1 => n1725, A2 => n1791, B1 => n5315, B2 => n1656
                           , ZN => n9723);
   U730 : OAI22_X1 port map( A1 => n1768, A2 => n1791, B1 => n5314, B2 => n1656
                           , ZN => n9722);
   U731 : OAI21_X1 port map( B1 => n1769, B2 => n1791, A => n1770, ZN => n1792)
                           ;
   U732 : OAI22_X1 port map( A1 => n1759, A2 => n1794, B1 => n5313, B2 => n1650
                           , ZN => n9721);
   U733 : OAI22_X1 port map( A1 => n1761, A2 => n1794, B1 => n5312, B2 => n1650
                           , ZN => n9720);
   U734 : OAI22_X1 port map( A1 => n1762, A2 => n1794, B1 => n5311, B2 => n1650
                           , ZN => n9719);
   U735 : OAI22_X1 port map( A1 => n1763, A2 => n1794, B1 => n5310, B2 => n1650
                           , ZN => n9718);
   U736 : OAI22_X1 port map( A1 => n1764, A2 => n1794, B1 => n5309, B2 => n1650
                           , ZN => n9717);
   U737 : OAI22_X1 port map( A1 => n1765, A2 => n1794, B1 => n5308, B2 => n1650
                           , ZN => n9716);
   U738 : OAI22_X1 port map( A1 => n1766, A2 => n1794, B1 => n5307, B2 => n1650
                           , ZN => n9715);
   U739 : OAI22_X1 port map( A1 => n1767, A2 => n1794, B1 => n5306, B2 => n1650
                           , ZN => n9714);
   U740 : OAI22_X1 port map( A1 => n1746, A2 => n1794, B1 => n5305, B2 => n1650
                           , ZN => n9713);
   U741 : OAI22_X1 port map( A1 => n1747, A2 => n1794, B1 => n5304, B2 => n1650
                           , ZN => n9712);
   U742 : OAI22_X1 port map( A1 => n1742, A2 => n1794, B1 => n5303, B2 => n1650
                           , ZN => n9711);
   U743 : OAI22_X1 port map( A1 => n1743, A2 => n1794, B1 => n5302, B2 => n1650
                           , ZN => n9710);
   U744 : OAI22_X1 port map( A1 => n1744, A2 => n1794, B1 => n5301, B2 => n1650
                           , ZN => n9709);
   U745 : OAI22_X1 port map( A1 => n1745, A2 => n1794, B1 => n5300, B2 => n1650
                           , ZN => n9708);
   U746 : OAI22_X1 port map( A1 => n1738, A2 => n1794, B1 => n5299, B2 => n1650
                           , ZN => n9707);
   U747 : OAI22_X1 port map( A1 => n1739, A2 => n1794, B1 => n5298, B2 => n1650
                           , ZN => n9706);
   U748 : OAI22_X1 port map( A1 => n1740, A2 => n1794, B1 => n5297, B2 => n1650
                           , ZN => n9705);
   U749 : OAI22_X1 port map( A1 => n1741, A2 => n1794, B1 => n5296, B2 => n1650
                           , ZN => n9704);
   U750 : OAI22_X1 port map( A1 => n1734, A2 => n1794, B1 => n5295, B2 => n1650
                           , ZN => n9703);
   U751 : OAI22_X1 port map( A1 => n1735, A2 => n1794, B1 => n5294, B2 => n1650
                           , ZN => n9702);
   U752 : OAI22_X1 port map( A1 => n1736, A2 => n1794, B1 => n5293, B2 => n1650
                           , ZN => n9701);
   U753 : OAI22_X1 port map( A1 => n1737, A2 => n1794, B1 => n5292, B2 => n1650
                           , ZN => n9700);
   U754 : OAI22_X1 port map( A1 => n1730, A2 => n1794, B1 => n5291, B2 => n1650
                           , ZN => n9699);
   U755 : OAI22_X1 port map( A1 => n1731, A2 => n1794, B1 => n5290, B2 => n1650
                           , ZN => n9698);
   U756 : OAI22_X1 port map( A1 => n1732, A2 => n1794, B1 => n5289, B2 => n1650
                           , ZN => n9697);
   U757 : OAI22_X1 port map( A1 => n1733, A2 => n1794, B1 => n5288, B2 => n1650
                           , ZN => n9696);
   U758 : OAI22_X1 port map( A1 => n1726, A2 => n1794, B1 => n5287, B2 => n1650
                           , ZN => n9695);
   U759 : OAI22_X1 port map( A1 => n1727, A2 => n1794, B1 => n5286, B2 => n1650
                           , ZN => n9694);
   U760 : OAI22_X1 port map( A1 => n1728, A2 => n1794, B1 => n5285, B2 => n1650
                           , ZN => n9693);
   U761 : OAI22_X1 port map( A1 => n1729, A2 => n1794, B1 => n5284, B2 => n1650
                           , ZN => n9692);
   U762 : OAI22_X1 port map( A1 => n1725, A2 => n1794, B1 => n5283, B2 => n1650
                           , ZN => n9691);
   U763 : OAI22_X1 port map( A1 => n1768, A2 => n1794, B1 => n5282, B2 => n1650
                           , ZN => n9690);
   U764 : OAI21_X1 port map( B1 => n1769, B2 => n1794, A => n1770, ZN => n1795)
                           ;
   U765 : OAI22_X1 port map( A1 => n1759, A2 => n1797, B1 => n1714, B2 => n617,
                           ZN => n9689);
   U766 : OAI22_X1 port map( A1 => n1761, A2 => n1797, B1 => n1714, B2 => n620,
                           ZN => n9688);
   U767 : OAI22_X1 port map( A1 => n1762, A2 => n1797, B1 => n1714, B2 => n623,
                           ZN => n9687);
   U768 : OAI22_X1 port map( A1 => n1763, A2 => n1797, B1 => n1714, B2 => n626,
                           ZN => n9686);
   U769 : OAI22_X1 port map( A1 => n1764, A2 => n1797, B1 => n1714, B2 => n629,
                           ZN => n9685);
   U770 : OAI22_X1 port map( A1 => n1765, A2 => n1797, B1 => n1714, B2 => n632,
                           ZN => n9684);
   U771 : OAI22_X1 port map( A1 => n1766, A2 => n1797, B1 => n1714, B2 => n635,
                           ZN => n9683);
   U772 : OAI22_X1 port map( A1 => n1767, A2 => n1797, B1 => n1714, B2 => n638,
                           ZN => n9682);
   U773 : OAI22_X1 port map( A1 => n1746, A2 => n1797, B1 => n1714, B2 => n641,
                           ZN => n9681);
   U774 : OAI22_X1 port map( A1 => n1747, A2 => n1797, B1 => n1714, B2 => n644,
                           ZN => n9680);
   U775 : OAI22_X1 port map( A1 => n1742, A2 => n1797, B1 => n1714, B2 => n647,
                           ZN => n9679);
   U776 : OAI22_X1 port map( A1 => n1743, A2 => n1797, B1 => n1714, B2 => n650,
                           ZN => n9678);
   U777 : OAI22_X1 port map( A1 => n1744, A2 => n1797, B1 => n1714, B2 => n653,
                           ZN => n9677);
   U778 : OAI22_X1 port map( A1 => n1745, A2 => n1797, B1 => n1714, B2 => n656,
                           ZN => n9676);
   U779 : OAI22_X1 port map( A1 => n1738, A2 => n1797, B1 => n1714, B2 => n659,
                           ZN => n9675);
   U780 : OAI22_X1 port map( A1 => n1739, A2 => n1797, B1 => n1714, B2 => n662,
                           ZN => n9674);
   U781 : OAI22_X1 port map( A1 => n1740, A2 => n1797, B1 => n1714, B2 => n665,
                           ZN => n9673);
   U782 : OAI22_X1 port map( A1 => n1741, A2 => n1797, B1 => n1714, B2 => n668,
                           ZN => n9672);
   U783 : OAI22_X1 port map( A1 => n1734, A2 => n1797, B1 => n1714, B2 => n671,
                           ZN => n9671);
   U784 : OAI22_X1 port map( A1 => n1735, A2 => n1797, B1 => n1714, B2 => n674,
                           ZN => n9670);
   U785 : OAI22_X1 port map( A1 => n1736, A2 => n1797, B1 => n1714, B2 => n677,
                           ZN => n9669);
   U786 : OAI22_X1 port map( A1 => n1737, A2 => n1797, B1 => n1714, B2 => n680,
                           ZN => n9668);
   U787 : OAI22_X1 port map( A1 => n1730, A2 => n1797, B1 => n1714, B2 => n683,
                           ZN => n9667);
   U788 : OAI22_X1 port map( A1 => n1731, A2 => n1797, B1 => n1714, B2 => n686,
                           ZN => n9666);
   U789 : OAI22_X1 port map( A1 => n1732, A2 => n1797, B1 => n1714, B2 => n689,
                           ZN => n9665);
   U790 : OAI22_X1 port map( A1 => n1733, A2 => n1797, B1 => n1714, B2 => n692,
                           ZN => n9664);
   U791 : OAI22_X1 port map( A1 => n1726, A2 => n1797, B1 => n1714, B2 => n695,
                           ZN => n9663);
   U792 : OAI22_X1 port map( A1 => n1727, A2 => n1797, B1 => n1714, B2 => n698,
                           ZN => n9662);
   U793 : OAI22_X1 port map( A1 => n1728, A2 => n1797, B1 => n1714, B2 => n701,
                           ZN => n9661);
   U794 : OAI22_X1 port map( A1 => n1729, A2 => n1797, B1 => n1714, B2 => n704,
                           ZN => n9660);
   U795 : OAI22_X1 port map( A1 => n1725, A2 => n1797, B1 => n1714, B2 => n707,
                           ZN => n9659);
   U796 : OAI22_X1 port map( A1 => n1768, A2 => n1797, B1 => n1714, B2 => n710,
                           ZN => n9658);
   U797 : OAI21_X1 port map( B1 => n1769, B2 => n1797, A => n1770, ZN => n1798)
                           ;
   U798 : OAI22_X1 port map( A1 => n1759, A2 => n1800, B1 => n1716, B2 => n193,
                           ZN => n9657);
   U799 : OAI22_X1 port map( A1 => n1761, A2 => n1800, B1 => n1716, B2 => n196,
                           ZN => n9656);
   U800 : OAI22_X1 port map( A1 => n1762, A2 => n1800, B1 => n1716, B2 => n199,
                           ZN => n9655);
   U801 : OAI22_X1 port map( A1 => n1763, A2 => n1800, B1 => n1716, B2 => n202,
                           ZN => n9654);
   U802 : OAI22_X1 port map( A1 => n1764, A2 => n1800, B1 => n1716, B2 => n205,
                           ZN => n9653);
   U803 : OAI22_X1 port map( A1 => n1765, A2 => n1800, B1 => n1716, B2 => n208,
                           ZN => n9652);
   U804 : OAI22_X1 port map( A1 => n1766, A2 => n1800, B1 => n1716, B2 => n211,
                           ZN => n9651);
   U805 : OAI22_X1 port map( A1 => n1767, A2 => n1800, B1 => n1716, B2 => n214,
                           ZN => n9650);
   U806 : OAI22_X1 port map( A1 => n1746, A2 => n1800, B1 => n1716, B2 => n217,
                           ZN => n9649);
   U807 : OAI22_X1 port map( A1 => n1747, A2 => n1800, B1 => n1716, B2 => n220,
                           ZN => n9648);
   U808 : OAI22_X1 port map( A1 => n1742, A2 => n1800, B1 => n1716, B2 => n223,
                           ZN => n9647);
   U809 : OAI22_X1 port map( A1 => n1743, A2 => n1800, B1 => n1716, B2 => n226,
                           ZN => n9646);
   U810 : OAI22_X1 port map( A1 => n1744, A2 => n1800, B1 => n1716, B2 => n229,
                           ZN => n9645);
   U811 : OAI22_X1 port map( A1 => n1745, A2 => n1800, B1 => n1716, B2 => n232,
                           ZN => n9644);
   U812 : OAI22_X1 port map( A1 => n1738, A2 => n1800, B1 => n1716, B2 => n235,
                           ZN => n9643);
   U813 : OAI22_X1 port map( A1 => n1739, A2 => n1800, B1 => n1716, B2 => n238,
                           ZN => n9642);
   U814 : OAI22_X1 port map( A1 => n1740, A2 => n1800, B1 => n1716, B2 => n241,
                           ZN => n9641);
   U815 : OAI22_X1 port map( A1 => n1741, A2 => n1800, B1 => n1716, B2 => n244,
                           ZN => n9640);
   U816 : OAI22_X1 port map( A1 => n1734, A2 => n1800, B1 => n1716, B2 => n247,
                           ZN => n9639);
   U817 : OAI22_X1 port map( A1 => n1735, A2 => n1800, B1 => n1716, B2 => n250,
                           ZN => n9638);
   U818 : OAI22_X1 port map( A1 => n1736, A2 => n1800, B1 => n1716, B2 => n253,
                           ZN => n9637);
   U819 : OAI22_X1 port map( A1 => n1737, A2 => n1800, B1 => n1716, B2 => n256,
                           ZN => n9636);
   U820 : OAI22_X1 port map( A1 => n1730, A2 => n1800, B1 => n1716, B2 => n259,
                           ZN => n9635);
   U821 : OAI22_X1 port map( A1 => n1731, A2 => n1800, B1 => n1716, B2 => n262,
                           ZN => n9634);
   U822 : OAI22_X1 port map( A1 => n1732, A2 => n1800, B1 => n1716, B2 => n265,
                           ZN => n9633);
   U823 : OAI22_X1 port map( A1 => n1733, A2 => n1800, B1 => n1716, B2 => n268,
                           ZN => n9632);
   U824 : OAI22_X1 port map( A1 => n1726, A2 => n1800, B1 => n1716, B2 => n271,
                           ZN => n9631);
   U825 : OAI22_X1 port map( A1 => n1727, A2 => n1800, B1 => n1716, B2 => n274,
                           ZN => n9630);
   U826 : OAI22_X1 port map( A1 => n1728, A2 => n1800, B1 => n1716, B2 => n277,
                           ZN => n9629);
   U827 : OAI22_X1 port map( A1 => n1729, A2 => n1800, B1 => n1716, B2 => n280,
                           ZN => n9628);
   U828 : OAI22_X1 port map( A1 => n1725, A2 => n1800, B1 => n1716, B2 => n283,
                           ZN => n9627);
   U829 : OAI22_X1 port map( A1 => n1768, A2 => n1800, B1 => n1716, B2 => n286,
                           ZN => n9626);
   U830 : OAI21_X1 port map( B1 => n1769, B2 => n1800, A => n1770, ZN => n1801)
                           ;
   U831 : OAI22_X1 port map( A1 => n1759, A2 => n1803, B1 => n5694, B2 => n1652
                           , ZN => n9625);
   U832 : OAI22_X1 port map( A1 => n1761, A2 => n1803, B1 => n5684, B2 => n1652
                           , ZN => n9624);
   U833 : OAI22_X1 port map( A1 => n1762, A2 => n1803, B1 => n5674, B2 => n1652
                           , ZN => n9623);
   U834 : OAI22_X1 port map( A1 => n1763, A2 => n1803, B1 => n5664, B2 => n1652
                           , ZN => n9622);
   U835 : OAI22_X1 port map( A1 => n1764, A2 => n1803, B1 => n5654, B2 => n1652
                           , ZN => n9621);
   U836 : OAI22_X1 port map( A1 => n1765, A2 => n1803, B1 => n5644, B2 => n1652
                           , ZN => n9620);
   U837 : OAI22_X1 port map( A1 => n1766, A2 => n1803, B1 => n5634, B2 => n1652
                           , ZN => n9619);
   U838 : OAI22_X1 port map( A1 => n1767, A2 => n1803, B1 => n5624, B2 => n1652
                           , ZN => n9618);
   U839 : OAI22_X1 port map( A1 => n1746, A2 => n1803, B1 => n5614, B2 => n1652
                           , ZN => n9617);
   U840 : OAI22_X1 port map( A1 => n1747, A2 => n1803, B1 => n5604, B2 => n1652
                           , ZN => n9616);
   U841 : OAI22_X1 port map( A1 => n1742, A2 => n1803, B1 => n5594, B2 => n1652
                           , ZN => n9615);
   U842 : OAI22_X1 port map( A1 => n1743, A2 => n1803, B1 => n5584, B2 => n1652
                           , ZN => n9614);
   U843 : OAI22_X1 port map( A1 => n1744, A2 => n1803, B1 => n5574, B2 => n1652
                           , ZN => n9613);
   U844 : OAI22_X1 port map( A1 => n1745, A2 => n1803, B1 => n5564, B2 => n1652
                           , ZN => n9612);
   U845 : OAI22_X1 port map( A1 => n1738, A2 => n1803, B1 => n5554, B2 => n1652
                           , ZN => n9611);
   U846 : OAI22_X1 port map( A1 => n1739, A2 => n1803, B1 => n5544, B2 => n1652
                           , ZN => n9610);
   U847 : OAI22_X1 port map( A1 => n1740, A2 => n1803, B1 => n5534, B2 => n1652
                           , ZN => n9609);
   U848 : OAI22_X1 port map( A1 => n1741, A2 => n1803, B1 => n5524, B2 => n1652
                           , ZN => n9608);
   U849 : OAI22_X1 port map( A1 => n1734, A2 => n1803, B1 => n5514, B2 => n1652
                           , ZN => n9607);
   U850 : OAI22_X1 port map( A1 => n1735, A2 => n1803, B1 => n5504, B2 => n1652
                           , ZN => n9606);
   U851 : OAI22_X1 port map( A1 => n1736, A2 => n1803, B1 => n5494, B2 => n1652
                           , ZN => n9605);
   U852 : OAI22_X1 port map( A1 => n1737, A2 => n1803, B1 => n5484, B2 => n1652
                           , ZN => n9604);
   U853 : OAI22_X1 port map( A1 => n1730, A2 => n1803, B1 => n5474, B2 => n1652
                           , ZN => n9603);
   U854 : OAI22_X1 port map( A1 => n1731, A2 => n1803, B1 => n5464, B2 => n1652
                           , ZN => n9602);
   U855 : OAI22_X1 port map( A1 => n1732, A2 => n1803, B1 => n5454, B2 => n1652
                           , ZN => n9601);
   U856 : OAI22_X1 port map( A1 => n1733, A2 => n1803, B1 => n5444, B2 => n1652
                           , ZN => n9600);
   U857 : OAI22_X1 port map( A1 => n1726, A2 => n1803, B1 => n5434, B2 => n1652
                           , ZN => n9599);
   U858 : OAI22_X1 port map( A1 => n1727, A2 => n1803, B1 => n5424, B2 => n1652
                           , ZN => n9598);
   U859 : OAI22_X1 port map( A1 => n1728, A2 => n1803, B1 => n5414, B2 => n1652
                           , ZN => n9597);
   U860 : OAI22_X1 port map( A1 => n1729, A2 => n1803, B1 => n5404, B2 => n1652
                           , ZN => n9596);
   U861 : OAI22_X1 port map( A1 => n1725, A2 => n1803, B1 => n5394, B2 => n1652
                           , ZN => n9595);
   U862 : OAI22_X1 port map( A1 => n1768, A2 => n1803, B1 => n5384, B2 => n1652
                           , ZN => n9594);
   U863 : OAI21_X1 port map( B1 => n1769, B2 => n1803, A => n1770, ZN => n1804)
                           ;
   U864 : OAI22_X1 port map( A1 => n1759, A2 => n1806, B1 => n5695, B2 => n1646
                           , ZN => n9593);
   U865 : OAI22_X1 port map( A1 => n1761, A2 => n1806, B1 => n5685, B2 => n1646
                           , ZN => n9592);
   U866 : OAI22_X1 port map( A1 => n1762, A2 => n1806, B1 => n5675, B2 => n1646
                           , ZN => n9591);
   U867 : OAI22_X1 port map( A1 => n1763, A2 => n1806, B1 => n5665, B2 => n1646
                           , ZN => n9590);
   U868 : OAI22_X1 port map( A1 => n1764, A2 => n1806, B1 => n5655, B2 => n1646
                           , ZN => n9589);
   U869 : OAI22_X1 port map( A1 => n1765, A2 => n1806, B1 => n5645, B2 => n1646
                           , ZN => n9588);
   U870 : OAI22_X1 port map( A1 => n1766, A2 => n1806, B1 => n5635, B2 => n1646
                           , ZN => n9587);
   U871 : OAI22_X1 port map( A1 => n1767, A2 => n1806, B1 => n5625, B2 => n1646
                           , ZN => n9586);
   U872 : OAI22_X1 port map( A1 => n1746, A2 => n1806, B1 => n5615, B2 => n1646
                           , ZN => n9585);
   U873 : OAI22_X1 port map( A1 => n1747, A2 => n1806, B1 => n5605, B2 => n1646
                           , ZN => n9584);
   U874 : OAI22_X1 port map( A1 => n1742, A2 => n1806, B1 => n5595, B2 => n1646
                           , ZN => n9583);
   U875 : OAI22_X1 port map( A1 => n1743, A2 => n1806, B1 => n5585, B2 => n1646
                           , ZN => n9582);
   U876 : OAI22_X1 port map( A1 => n1744, A2 => n1806, B1 => n5575, B2 => n1646
                           , ZN => n9581);
   U877 : OAI22_X1 port map( A1 => n1745, A2 => n1806, B1 => n5565, B2 => n1646
                           , ZN => n9580);
   U878 : OAI22_X1 port map( A1 => n1738, A2 => n1806, B1 => n5555, B2 => n1646
                           , ZN => n9579);
   U879 : OAI22_X1 port map( A1 => n1739, A2 => n1806, B1 => n5545, B2 => n1646
                           , ZN => n9578);
   U880 : OAI22_X1 port map( A1 => n1740, A2 => n1806, B1 => n5535, B2 => n1646
                           , ZN => n9577);
   U881 : OAI22_X1 port map( A1 => n1741, A2 => n1806, B1 => n5525, B2 => n1646
                           , ZN => n9576);
   U882 : OAI22_X1 port map( A1 => n1734, A2 => n1806, B1 => n5515, B2 => n1646
                           , ZN => n9575);
   U883 : OAI22_X1 port map( A1 => n1735, A2 => n1806, B1 => n5505, B2 => n1646
                           , ZN => n9574);
   U884 : OAI22_X1 port map( A1 => n1736, A2 => n1806, B1 => n5495, B2 => n1646
                           , ZN => n9573);
   U885 : OAI22_X1 port map( A1 => n1737, A2 => n1806, B1 => n5485, B2 => n1646
                           , ZN => n9572);
   U886 : OAI22_X1 port map( A1 => n1730, A2 => n1806, B1 => n5475, B2 => n1646
                           , ZN => n9571);
   U887 : OAI22_X1 port map( A1 => n1731, A2 => n1806, B1 => n5465, B2 => n1646
                           , ZN => n9570);
   U888 : OAI22_X1 port map( A1 => n1732, A2 => n1806, B1 => n5455, B2 => n1646
                           , ZN => n9569);
   U889 : OAI22_X1 port map( A1 => n1733, A2 => n1806, B1 => n5445, B2 => n1646
                           , ZN => n9568);
   U890 : OAI22_X1 port map( A1 => n1726, A2 => n1806, B1 => n5435, B2 => n1646
                           , ZN => n9567);
   U891 : OAI22_X1 port map( A1 => n1727, A2 => n1806, B1 => n5425, B2 => n1646
                           , ZN => n9566);
   U892 : OAI22_X1 port map( A1 => n1728, A2 => n1806, B1 => n5415, B2 => n1646
                           , ZN => n9565);
   U893 : OAI22_X1 port map( A1 => n1729, A2 => n1806, B1 => n5405, B2 => n1646
                           , ZN => n9564);
   U894 : OAI22_X1 port map( A1 => n1725, A2 => n1806, B1 => n5395, B2 => n1646
                           , ZN => n9563);
   U895 : OAI22_X1 port map( A1 => n1768, A2 => n1806, B1 => n5385, B2 => n1646
                           , ZN => n9562);
   U896 : OAI21_X1 port map( B1 => n1769, B2 => n1806, A => n1770, ZN => n1807)
                           ;
   U897 : OAI22_X1 port map( A1 => n1759, A2 => n1809, B1 => n1710, B2 => n841,
                           ZN => n9561);
   U898 : OAI22_X1 port map( A1 => n1761, A2 => n1809, B1 => n1710, B2 => n842,
                           ZN => n9560);
   U899 : OAI22_X1 port map( A1 => n1762, A2 => n1809, B1 => n1710, B2 => n843,
                           ZN => n9559);
   U900 : OAI22_X1 port map( A1 => n1763, A2 => n1809, B1 => n1710, B2 => n844,
                           ZN => n9558);
   U901 : OAI22_X1 port map( A1 => n1764, A2 => n1809, B1 => n1710, B2 => n845,
                           ZN => n9557);
   U902 : OAI22_X1 port map( A1 => n1765, A2 => n1809, B1 => n1710, B2 => n846,
                           ZN => n9556);
   U903 : OAI22_X1 port map( A1 => n1766, A2 => n1809, B1 => n1710, B2 => n847,
                           ZN => n9555);
   U904 : OAI22_X1 port map( A1 => n1767, A2 => n1809, B1 => n1710, B2 => n848,
                           ZN => n9554);
   U905 : OAI22_X1 port map( A1 => n1746, A2 => n1809, B1 => n1710, B2 => n849,
                           ZN => n9553);
   U906 : OAI22_X1 port map( A1 => n1747, A2 => n1809, B1 => n1710, B2 => n850,
                           ZN => n9552);
   U907 : OAI22_X1 port map( A1 => n1742, A2 => n1809, B1 => n1710, B2 => n851,
                           ZN => n9551);
   U908 : OAI22_X1 port map( A1 => n1743, A2 => n1809, B1 => n1710, B2 => n852,
                           ZN => n9550);
   U909 : OAI22_X1 port map( A1 => n1744, A2 => n1809, B1 => n1710, B2 => n853,
                           ZN => n9549);
   U910 : OAI22_X1 port map( A1 => n1745, A2 => n1809, B1 => n1710, B2 => n854,
                           ZN => n9548);
   U911 : OAI22_X1 port map( A1 => n1738, A2 => n1809, B1 => n1710, B2 => n855,
                           ZN => n9547);
   U912 : OAI22_X1 port map( A1 => n1739, A2 => n1809, B1 => n1710, B2 => n856,
                           ZN => n9546);
   U913 : OAI22_X1 port map( A1 => n1740, A2 => n1809, B1 => n1710, B2 => n857,
                           ZN => n9545);
   U914 : OAI22_X1 port map( A1 => n1741, A2 => n1809, B1 => n1710, B2 => n858,
                           ZN => n9544);
   U915 : OAI22_X1 port map( A1 => n1734, A2 => n1809, B1 => n1710, B2 => n859,
                           ZN => n9543);
   U916 : OAI22_X1 port map( A1 => n1735, A2 => n1809, B1 => n1710, B2 => n860,
                           ZN => n9542);
   U917 : OAI22_X1 port map( A1 => n1736, A2 => n1809, B1 => n1710, B2 => n861,
                           ZN => n9541);
   U918 : OAI22_X1 port map( A1 => n1737, A2 => n1809, B1 => n1710, B2 => n862,
                           ZN => n9540);
   U919 : OAI22_X1 port map( A1 => n1730, A2 => n1809, B1 => n1710, B2 => n863,
                           ZN => n9539);
   U920 : OAI22_X1 port map( A1 => n1731, A2 => n1809, B1 => n1710, B2 => n864,
                           ZN => n9538);
   U921 : OAI22_X1 port map( A1 => n1732, A2 => n1809, B1 => n1710, B2 => n865,
                           ZN => n9537);
   U922 : OAI22_X1 port map( A1 => n1733, A2 => n1809, B1 => n1710, B2 => n866,
                           ZN => n9536);
   U923 : OAI22_X1 port map( A1 => n1726, A2 => n1809, B1 => n1710, B2 => n867,
                           ZN => n9535);
   U924 : OAI22_X1 port map( A1 => n1727, A2 => n1809, B1 => n1710, B2 => n868,
                           ZN => n9534);
   U925 : OAI22_X1 port map( A1 => n1728, A2 => n1809, B1 => n1710, B2 => n869,
                           ZN => n9533);
   U926 : OAI22_X1 port map( A1 => n1729, A2 => n1809, B1 => n1710, B2 => n870,
                           ZN => n9532);
   U927 : OAI22_X1 port map( A1 => n1725, A2 => n1809, B1 => n1710, B2 => n871,
                           ZN => n9531);
   U928 : OAI22_X1 port map( A1 => n1768, A2 => n1809, B1 => n1710, B2 => n872,
                           ZN => n9530);
   U929 : OAI21_X1 port map( B1 => n1769, B2 => n1809, A => n1770, ZN => n1810)
                           ;
   U930 : OAI22_X1 port map( A1 => n1759, A2 => n1812, B1 => n1712, B2 => n1193
                           , ZN => n9529);
   U931 : OAI22_X1 port map( A1 => n1761, A2 => n1812, B1 => n1712, B2 => n1194
                           , ZN => n9528);
   U932 : OAI22_X1 port map( A1 => n1762, A2 => n1812, B1 => n1712, B2 => n1195
                           , ZN => n9527);
   U933 : OAI22_X1 port map( A1 => n1763, A2 => n1812, B1 => n1712, B2 => n1196
                           , ZN => n9526);
   U934 : OAI22_X1 port map( A1 => n1764, A2 => n1812, B1 => n1712, B2 => n1197
                           , ZN => n9525);
   U935 : OAI22_X1 port map( A1 => n1765, A2 => n1812, B1 => n1712, B2 => n1198
                           , ZN => n9524);
   U936 : OAI22_X1 port map( A1 => n1766, A2 => n1812, B1 => n1712, B2 => n1199
                           , ZN => n9523);
   U937 : OAI22_X1 port map( A1 => n1767, A2 => n1812, B1 => n1712, B2 => n1200
                           , ZN => n9522);
   U938 : OAI22_X1 port map( A1 => n1746, A2 => n1812, B1 => n1712, B2 => n1201
                           , ZN => n9521);
   U939 : OAI22_X1 port map( A1 => n1747, A2 => n1812, B1 => n1712, B2 => n1202
                           , ZN => n9520);
   U940 : OAI22_X1 port map( A1 => n1742, A2 => n1812, B1 => n1712, B2 => n1203
                           , ZN => n9519);
   U941 : OAI22_X1 port map( A1 => n1743, A2 => n1812, B1 => n1712, B2 => n1204
                           , ZN => n9518);
   U942 : OAI22_X1 port map( A1 => n1744, A2 => n1812, B1 => n1712, B2 => n1205
                           , ZN => n9517);
   U943 : OAI22_X1 port map( A1 => n1745, A2 => n1812, B1 => n1712, B2 => n1206
                           , ZN => n9516);
   U944 : OAI22_X1 port map( A1 => n1738, A2 => n1812, B1 => n1712, B2 => n1207
                           , ZN => n9515);
   U945 : OAI22_X1 port map( A1 => n1739, A2 => n1812, B1 => n1712, B2 => n1208
                           , ZN => n9514);
   U946 : OAI22_X1 port map( A1 => n1740, A2 => n1812, B1 => n1712, B2 => n1209
                           , ZN => n9513);
   U947 : OAI22_X1 port map( A1 => n1741, A2 => n1812, B1 => n1712, B2 => n1210
                           , ZN => n9512);
   U948 : OAI22_X1 port map( A1 => n1734, A2 => n1812, B1 => n1712, B2 => n1211
                           , ZN => n9511);
   U949 : OAI22_X1 port map( A1 => n1735, A2 => n1812, B1 => n1712, B2 => n1212
                           , ZN => n9510);
   U950 : OAI22_X1 port map( A1 => n1736, A2 => n1812, B1 => n1712, B2 => n1213
                           , ZN => n9509);
   U951 : OAI22_X1 port map( A1 => n1737, A2 => n1812, B1 => n1712, B2 => n1214
                           , ZN => n9508);
   U952 : OAI22_X1 port map( A1 => n1730, A2 => n1812, B1 => n1712, B2 => n1215
                           , ZN => n9507);
   U953 : OAI22_X1 port map( A1 => n1731, A2 => n1812, B1 => n1712, B2 => n1216
                           , ZN => n9506);
   U954 : OAI22_X1 port map( A1 => n1732, A2 => n1812, B1 => n1712, B2 => n1217
                           , ZN => n9505);
   U955 : OAI22_X1 port map( A1 => n1733, A2 => n1812, B1 => n1712, B2 => n1218
                           , ZN => n9504);
   U956 : OAI22_X1 port map( A1 => n1726, A2 => n1812, B1 => n1712, B2 => n1219
                           , ZN => n9503);
   U957 : OAI22_X1 port map( A1 => n1727, A2 => n1812, B1 => n1712, B2 => n1220
                           , ZN => n9502);
   U958 : OAI22_X1 port map( A1 => n1728, A2 => n1812, B1 => n1712, B2 => n1221
                           , ZN => n9501);
   U959 : OAI22_X1 port map( A1 => n1729, A2 => n1812, B1 => n1712, B2 => n1222
                           , ZN => n9500);
   U960 : OAI22_X1 port map( A1 => n1725, A2 => n1812, B1 => n1712, B2 => n1223
                           , ZN => n9499);
   U961 : OAI22_X1 port map( A1 => n1768, A2 => n1812, B1 => n1712, B2 => n1224
                           , ZN => n9498);
   U962 : OAI21_X1 port map( B1 => n1769, B2 => n1812, A => n1770, ZN => n1813)
                           ;
   U963 : OAI22_X1 port map( A1 => n1759, A2 => n1580, B1 => n5281, B2 => n1648
                           , ZN => n9497);
   U964 : OAI22_X1 port map( A1 => n1761, A2 => n1580, B1 => n5280, B2 => n1648
                           , ZN => n9496);
   U965 : OAI22_X1 port map( A1 => n1762, A2 => n1580, B1 => n5279, B2 => n1648
                           , ZN => n9495);
   U966 : OAI22_X1 port map( A1 => n1763, A2 => n1580, B1 => n5278, B2 => n1648
                           , ZN => n9494);
   U967 : OAI22_X1 port map( A1 => n1764, A2 => n1580, B1 => n5277, B2 => n1648
                           , ZN => n9493);
   U968 : OAI22_X1 port map( A1 => n1765, A2 => n1580, B1 => n5276, B2 => n1648
                           , ZN => n9492);
   U969 : OAI22_X1 port map( A1 => n1766, A2 => n1580, B1 => n5275, B2 => n1648
                           , ZN => n9491);
   U970 : OAI22_X1 port map( A1 => n1767, A2 => n1580, B1 => n5274, B2 => n1648
                           , ZN => n9490);
   U971 : OAI22_X1 port map( A1 => n1746, A2 => n1580, B1 => n5273, B2 => n1648
                           , ZN => n9489);
   U972 : OAI22_X1 port map( A1 => n1747, A2 => n1580, B1 => n5272, B2 => n1648
                           , ZN => n9488);
   U973 : OAI22_X1 port map( A1 => n1742, A2 => n1580, B1 => n5271, B2 => n1648
                           , ZN => n9487);
   U974 : OAI22_X1 port map( A1 => n1743, A2 => n1580, B1 => n5270, B2 => n1648
                           , ZN => n9486);
   U975 : OAI22_X1 port map( A1 => n1744, A2 => n1580, B1 => n5269, B2 => n1648
                           , ZN => n9485);
   U976 : OAI22_X1 port map( A1 => n1745, A2 => n1580, B1 => n5268, B2 => n1648
                           , ZN => n9484);
   U977 : OAI22_X1 port map( A1 => n1738, A2 => n1580, B1 => n5267, B2 => n1648
                           , ZN => n9483);
   U978 : OAI22_X1 port map( A1 => n1739, A2 => n1580, B1 => n5266, B2 => n1648
                           , ZN => n9482);
   U979 : OAI22_X1 port map( A1 => n1740, A2 => n1580, B1 => n5265, B2 => n1648
                           , ZN => n9481);
   U980 : OAI22_X1 port map( A1 => n1741, A2 => n1580, B1 => n5264, B2 => n1648
                           , ZN => n9480);
   U981 : OAI22_X1 port map( A1 => n1734, A2 => n1580, B1 => n5263, B2 => n1648
                           , ZN => n9479);
   U982 : OAI22_X1 port map( A1 => n1735, A2 => n1580, B1 => n5262, B2 => n1648
                           , ZN => n9478);
   U983 : OAI22_X1 port map( A1 => n1736, A2 => n1580, B1 => n5261, B2 => n1648
                           , ZN => n9477);
   U984 : OAI22_X1 port map( A1 => n1737, A2 => n1580, B1 => n5260, B2 => n1648
                           , ZN => n9476);
   U985 : OAI22_X1 port map( A1 => n1730, A2 => n1580, B1 => n5259, B2 => n1648
                           , ZN => n9475);
   U986 : OAI22_X1 port map( A1 => n1731, A2 => n1580, B1 => n5258, B2 => n1648
                           , ZN => n9474);
   U987 : OAI22_X1 port map( A1 => n1732, A2 => n1580, B1 => n5257, B2 => n1648
                           , ZN => n9473);
   U988 : OAI22_X1 port map( A1 => n1733, A2 => n1580, B1 => n5256, B2 => n1648
                           , ZN => n9472);
   U989 : OAI22_X1 port map( A1 => n1726, A2 => n1580, B1 => n5255, B2 => n1648
                           , ZN => n9471);
   U990 : OAI22_X1 port map( A1 => n1727, A2 => n1580, B1 => n5254, B2 => n1648
                           , ZN => n9470);
   U991 : OAI22_X1 port map( A1 => n1728, A2 => n1580, B1 => n5253, B2 => n1648
                           , ZN => n9469);
   U992 : OAI22_X1 port map( A1 => n1729, A2 => n1580, B1 => n5252, B2 => n1648
                           , ZN => n9468);
   U993 : OAI22_X1 port map( A1 => n1725, A2 => n1580, B1 => n5251, B2 => n1648
                           , ZN => n9467);
   U994 : OAI22_X1 port map( A1 => n1768, A2 => n1580, B1 => n5250, B2 => n1648
                           , ZN => n9466);
   U995 : OAI21_X1 port map( B1 => n1769, B2 => n1580, A => n1770, ZN => n1815)
                           ;
   U996 : OAI22_X1 port map( A1 => n1759, A2 => n1817, B1 => n5249, B2 => n1642
                           , ZN => n9465);
   U997 : OAI22_X1 port map( A1 => n1761, A2 => n1817, B1 => n5248, B2 => n1642
                           , ZN => n9464);
   U998 : OAI22_X1 port map( A1 => n1762, A2 => n1817, B1 => n5247, B2 => n1642
                           , ZN => n9463);
   U999 : OAI22_X1 port map( A1 => n1763, A2 => n1817, B1 => n5246, B2 => n1642
                           , ZN => n9462);
   U1000 : OAI22_X1 port map( A1 => n1764, A2 => n1817, B1 => n5245, B2 => 
                           n1642, ZN => n9461);
   U1001 : OAI22_X1 port map( A1 => n1765, A2 => n1817, B1 => n5244, B2 => 
                           n1642, ZN => n9460);
   U1002 : OAI22_X1 port map( A1 => n1766, A2 => n1817, B1 => n5243, B2 => 
                           n1642, ZN => n9459);
   U1003 : OAI22_X1 port map( A1 => n1767, A2 => n1817, B1 => n5242, B2 => 
                           n1642, ZN => n9458);
   U1004 : OAI22_X1 port map( A1 => n1746, A2 => n1817, B1 => n5241, B2 => 
                           n1642, ZN => n9457);
   U1005 : OAI22_X1 port map( A1 => n1747, A2 => n1817, B1 => n5240, B2 => 
                           n1642, ZN => n9456);
   U1006 : OAI22_X1 port map( A1 => n1742, A2 => n1817, B1 => n5239, B2 => 
                           n1642, ZN => n9455);
   U1007 : OAI22_X1 port map( A1 => n1743, A2 => n1817, B1 => n5238, B2 => 
                           n1642, ZN => n9454);
   U1008 : OAI22_X1 port map( A1 => n1744, A2 => n1817, B1 => n5237, B2 => 
                           n1642, ZN => n9453);
   U1009 : OAI22_X1 port map( A1 => n1745, A2 => n1817, B1 => n5236, B2 => 
                           n1642, ZN => n9452);
   U1010 : OAI22_X1 port map( A1 => n1738, A2 => n1817, B1 => n5235, B2 => 
                           n1642, ZN => n9451);
   U1011 : OAI22_X1 port map( A1 => n1739, A2 => n1817, B1 => n5234, B2 => 
                           n1642, ZN => n9450);
   U1012 : OAI22_X1 port map( A1 => n1740, A2 => n1817, B1 => n5233, B2 => 
                           n1642, ZN => n9449);
   U1013 : OAI22_X1 port map( A1 => n1741, A2 => n1817, B1 => n5232, B2 => 
                           n1642, ZN => n9448);
   U1014 : OAI22_X1 port map( A1 => n1734, A2 => n1817, B1 => n5231, B2 => 
                           n1642, ZN => n9447);
   U1015 : OAI22_X1 port map( A1 => n1735, A2 => n1817, B1 => n5230, B2 => 
                           n1642, ZN => n9446);
   U1016 : OAI22_X1 port map( A1 => n1736, A2 => n1817, B1 => n5229, B2 => 
                           n1642, ZN => n9445);
   U1017 : OAI22_X1 port map( A1 => n1737, A2 => n1817, B1 => n5228, B2 => 
                           n1642, ZN => n9444);
   U1018 : OAI22_X1 port map( A1 => n1730, A2 => n1817, B1 => n5227, B2 => 
                           n1642, ZN => n9443);
   U1019 : OAI22_X1 port map( A1 => n1731, A2 => n1817, B1 => n5226, B2 => 
                           n1642, ZN => n9442);
   U1020 : OAI22_X1 port map( A1 => n1732, A2 => n1817, B1 => n5225, B2 => 
                           n1642, ZN => n9441);
   U1021 : OAI22_X1 port map( A1 => n1733, A2 => n1817, B1 => n5224, B2 => 
                           n1642, ZN => n9440);
   U1022 : OAI22_X1 port map( A1 => n1726, A2 => n1817, B1 => n5223, B2 => 
                           n1642, ZN => n9439);
   U1023 : OAI22_X1 port map( A1 => n1727, A2 => n1817, B1 => n5222, B2 => 
                           n1642, ZN => n9438);
   U1024 : OAI22_X1 port map( A1 => n1728, A2 => n1817, B1 => n5221, B2 => 
                           n1642, ZN => n9437);
   U1025 : OAI22_X1 port map( A1 => n1729, A2 => n1817, B1 => n5220, B2 => 
                           n1642, ZN => n9436);
   U1026 : OAI22_X1 port map( A1 => n1725, A2 => n1817, B1 => n5219, B2 => 
                           n1642, ZN => n9435);
   U1027 : OAI22_X1 port map( A1 => n1768, A2 => n1817, B1 => n5218, B2 => 
                           n1642, ZN => n9434);
   U1028 : OAI21_X1 port map( B1 => n1769, B2 => n1817, A => n1770, ZN => n1818
                           );
   U1029 : OAI22_X1 port map( A1 => n1759, A2 => n1820, B1 => n5217, B2 => 
                           n1644, ZN => n9433);
   U1030 : OAI22_X1 port map( A1 => n1761, A2 => n1820, B1 => n5216, B2 => 
                           n1644, ZN => n9432);
   U1031 : OAI22_X1 port map( A1 => n1762, A2 => n1820, B1 => n5215, B2 => 
                           n1644, ZN => n9431);
   U1032 : OAI22_X1 port map( A1 => n1763, A2 => n1820, B1 => n5214, B2 => 
                           n1644, ZN => n9430);
   U1033 : OAI22_X1 port map( A1 => n1764, A2 => n1820, B1 => n5213, B2 => 
                           n1644, ZN => n9429);
   U1034 : OAI22_X1 port map( A1 => n1765, A2 => n1820, B1 => n5212, B2 => 
                           n1644, ZN => n9428);
   U1035 : OAI22_X1 port map( A1 => n1766, A2 => n1820, B1 => n5211, B2 => 
                           n1644, ZN => n9427);
   U1036 : OAI22_X1 port map( A1 => n1767, A2 => n1820, B1 => n5210, B2 => 
                           n1644, ZN => n9426);
   U1037 : OAI22_X1 port map( A1 => n1746, A2 => n1820, B1 => n5209, B2 => 
                           n1644, ZN => n9425);
   U1038 : OAI22_X1 port map( A1 => n1747, A2 => n1820, B1 => n5208, B2 => 
                           n1644, ZN => n9424);
   U1039 : OAI22_X1 port map( A1 => n1742, A2 => n1820, B1 => n5207, B2 => 
                           n1644, ZN => n9423);
   U1040 : OAI22_X1 port map( A1 => n1743, A2 => n1820, B1 => n5206, B2 => 
                           n1644, ZN => n9422);
   U1041 : OAI22_X1 port map( A1 => n1744, A2 => n1820, B1 => n5205, B2 => 
                           n1644, ZN => n9421);
   U1042 : OAI22_X1 port map( A1 => n1745, A2 => n1820, B1 => n5204, B2 => 
                           n1644, ZN => n9420);
   U1043 : OAI22_X1 port map( A1 => n1738, A2 => n1820, B1 => n5203, B2 => 
                           n1644, ZN => n9419);
   U1044 : OAI22_X1 port map( A1 => n1739, A2 => n1820, B1 => n5202, B2 => 
                           n1644, ZN => n9418);
   U1045 : OAI22_X1 port map( A1 => n1740, A2 => n1820, B1 => n5201, B2 => 
                           n1644, ZN => n9417);
   U1046 : OAI22_X1 port map( A1 => n1741, A2 => n1820, B1 => n5200, B2 => 
                           n1644, ZN => n9416);
   U1047 : OAI22_X1 port map( A1 => n1734, A2 => n1820, B1 => n5199, B2 => 
                           n1644, ZN => n9415);
   U1048 : OAI22_X1 port map( A1 => n1735, A2 => n1820, B1 => n5198, B2 => 
                           n1644, ZN => n9414);
   U1049 : OAI22_X1 port map( A1 => n1736, A2 => n1820, B1 => n5197, B2 => 
                           n1644, ZN => n9413);
   U1050 : OAI22_X1 port map( A1 => n1737, A2 => n1820, B1 => n5196, B2 => 
                           n1644, ZN => n9412);
   U1051 : OAI22_X1 port map( A1 => n1730, A2 => n1820, B1 => n5195, B2 => 
                           n1644, ZN => n9411);
   U1052 : OAI22_X1 port map( A1 => n1731, A2 => n1820, B1 => n5194, B2 => 
                           n1644, ZN => n9410);
   U1053 : OAI22_X1 port map( A1 => n1732, A2 => n1820, B1 => n5193, B2 => 
                           n1644, ZN => n9409);
   U1054 : OAI22_X1 port map( A1 => n1733, A2 => n1820, B1 => n5192, B2 => 
                           n1644, ZN => n9408);
   U1055 : OAI22_X1 port map( A1 => n1726, A2 => n1820, B1 => n5191, B2 => 
                           n1644, ZN => n9407);
   U1056 : OAI22_X1 port map( A1 => n1727, A2 => n1820, B1 => n5190, B2 => 
                           n1644, ZN => n9406);
   U1057 : OAI22_X1 port map( A1 => n1728, A2 => n1820, B1 => n5189, B2 => 
                           n1644, ZN => n9405);
   U1058 : OAI22_X1 port map( A1 => n1729, A2 => n1820, B1 => n5188, B2 => 
                           n1644, ZN => n9404);
   U1059 : OAI22_X1 port map( A1 => n1725, A2 => n1820, B1 => n5187, B2 => 
                           n1644, ZN => n9403);
   U1060 : OAI22_X1 port map( A1 => n1768, A2 => n1820, B1 => n5186, B2 => 
                           n1644, ZN => n9402);
   U1061 : OAI21_X1 port map( B1 => n1769, B2 => n1820, A => n1770, ZN => n1821
                           );
   U1062 : OAI22_X1 port map( A1 => n1759, A2 => n1822, B1 => n1706, B2 => n457
                           , ZN => n9401);
   U1063 : OAI22_X1 port map( A1 => n1761, A2 => n1822, B1 => n1706, B2 => n459
                           , ZN => n9400);
   U1064 : OAI22_X1 port map( A1 => n1762, A2 => n1822, B1 => n1706, B2 => n461
                           , ZN => n9399);
   U1065 : OAI22_X1 port map( A1 => n1763, A2 => n1822, B1 => n1706, B2 => n463
                           , ZN => n9398);
   U1066 : OAI22_X1 port map( A1 => n1764, A2 => n1822, B1 => n1706, B2 => n465
                           , ZN => n9397);
   U1067 : OAI22_X1 port map( A1 => n1765, A2 => n1822, B1 => n1706, B2 => n467
                           , ZN => n9396);
   U1068 : OAI22_X1 port map( A1 => n1766, A2 => n1822, B1 => n1706, B2 => n469
                           , ZN => n9395);
   U1069 : OAI22_X1 port map( A1 => n1767, A2 => n1822, B1 => n1706, B2 => n471
                           , ZN => n9394);
   U1070 : OAI22_X1 port map( A1 => n1746, A2 => n1822, B1 => n1706, B2 => n473
                           , ZN => n9393);
   U1071 : OAI22_X1 port map( A1 => n1747, A2 => n1822, B1 => n1706, B2 => n475
                           , ZN => n9392);
   U1072 : OAI22_X1 port map( A1 => n1742, A2 => n1822, B1 => n1706, B2 => n477
                           , ZN => n9391);
   U1073 : OAI22_X1 port map( A1 => n1743, A2 => n1822, B1 => n1706, B2 => n479
                           , ZN => n9390);
   U1074 : OAI22_X1 port map( A1 => n1744, A2 => n1822, B1 => n1706, B2 => n481
                           , ZN => n9389);
   U1075 : OAI22_X1 port map( A1 => n1745, A2 => n1822, B1 => n1706, B2 => n483
                           , ZN => n9388);
   U1076 : OAI22_X1 port map( A1 => n1738, A2 => n1822, B1 => n1706, B2 => n485
                           , ZN => n9387);
   U1077 : OAI22_X1 port map( A1 => n1739, A2 => n1822, B1 => n1706, B2 => n487
                           , ZN => n9386);
   U1078 : OAI22_X1 port map( A1 => n1740, A2 => n1822, B1 => n1706, B2 => n489
                           , ZN => n9385);
   U1079 : OAI22_X1 port map( A1 => n1741, A2 => n1822, B1 => n1706, B2 => n491
                           , ZN => n9384);
   U1080 : OAI22_X1 port map( A1 => n1734, A2 => n1822, B1 => n1706, B2 => n493
                           , ZN => n9383);
   U1081 : OAI22_X1 port map( A1 => n1735, A2 => n1822, B1 => n1706, B2 => n495
                           , ZN => n9382);
   U1082 : OAI22_X1 port map( A1 => n1736, A2 => n1822, B1 => n1706, B2 => n497
                           , ZN => n9381);
   U1083 : OAI22_X1 port map( A1 => n1737, A2 => n1822, B1 => n1706, B2 => n499
                           , ZN => n9380);
   U1084 : OAI22_X1 port map( A1 => n1730, A2 => n1822, B1 => n1706, B2 => n501
                           , ZN => n9379);
   U1085 : OAI22_X1 port map( A1 => n1731, A2 => n1822, B1 => n1706, B2 => n503
                           , ZN => n9378);
   U1086 : OAI22_X1 port map( A1 => n1732, A2 => n1822, B1 => n1706, B2 => n505
                           , ZN => n9377);
   U1087 : OAI22_X1 port map( A1 => n1733, A2 => n1822, B1 => n1706, B2 => n507
                           , ZN => n9376);
   U1088 : OAI22_X1 port map( A1 => n1726, A2 => n1822, B1 => n1706, B2 => n509
                           , ZN => n9375);
   U1089 : OAI22_X1 port map( A1 => n1727, A2 => n1822, B1 => n1706, B2 => n511
                           , ZN => n9374);
   U1090 : OAI22_X1 port map( A1 => n1728, A2 => n1822, B1 => n1706, B2 => n513
                           , ZN => n9373);
   U1091 : OAI22_X1 port map( A1 => n1729, A2 => n1822, B1 => n1706, B2 => n515
                           , ZN => n9372);
   U1092 : OAI22_X1 port map( A1 => n1725, A2 => n1822, B1 => n1706, B2 => n517
                           , ZN => n9371);
   U1093 : OAI22_X1 port map( A1 => n1768, A2 => n1822, B1 => n1706, B2 => n519
                           , ZN => n9370);
   U1094 : OAI21_X1 port map( B1 => n1769, B2 => n1822, A => n1770, ZN => n1823
                           );
   U1095 : OAI22_X1 port map( A1 => n1759, A2 => n1824, B1 => n1708, B2 => n1, 
                           ZN => n9369);
   U1096 : OAI22_X1 port map( A1 => n1761, A2 => n1824, B1 => n1708, B2 => n3, 
                           ZN => n9368);
   U1097 : OAI22_X1 port map( A1 => n1762, A2 => n1824, B1 => n1708, B2 => n5, 
                           ZN => n9367);
   U1098 : OAI22_X1 port map( A1 => n1763, A2 => n1824, B1 => n1708, B2 => n7, 
                           ZN => n9366);
   U1099 : OAI22_X1 port map( A1 => n1764, A2 => n1824, B1 => n1708, B2 => n9, 
                           ZN => n9365);
   U1100 : OAI22_X1 port map( A1 => n1765, A2 => n1824, B1 => n1708, B2 => n11,
                           ZN => n9364);
   U1101 : OAI22_X1 port map( A1 => n1766, A2 => n1824, B1 => n1708, B2 => n13,
                           ZN => n9363);
   U1102 : OAI22_X1 port map( A1 => n1767, A2 => n1824, B1 => n1708, B2 => n15,
                           ZN => n9362);
   U1103 : OAI22_X1 port map( A1 => n1746, A2 => n1824, B1 => n1708, B2 => n17,
                           ZN => n9361);
   U1104 : OAI22_X1 port map( A1 => n1747, A2 => n1824, B1 => n1708, B2 => n19,
                           ZN => n9360);
   U1105 : OAI22_X1 port map( A1 => n1742, A2 => n1824, B1 => n1708, B2 => n21,
                           ZN => n9359);
   U1106 : OAI22_X1 port map( A1 => n1743, A2 => n1824, B1 => n1708, B2 => n23,
                           ZN => n9358);
   U1107 : OAI22_X1 port map( A1 => n1744, A2 => n1824, B1 => n1708, B2 => n25,
                           ZN => n9357);
   U1108 : OAI22_X1 port map( A1 => n1745, A2 => n1824, B1 => n1708, B2 => n27,
                           ZN => n9356);
   U1109 : OAI22_X1 port map( A1 => n1738, A2 => n1824, B1 => n1708, B2 => n29,
                           ZN => n9355);
   U1110 : OAI22_X1 port map( A1 => n1739, A2 => n1824, B1 => n1708, B2 => n31,
                           ZN => n9354);
   U1111 : OAI22_X1 port map( A1 => n1740, A2 => n1824, B1 => n1708, B2 => n33,
                           ZN => n9353);
   U1112 : OAI22_X1 port map( A1 => n1741, A2 => n1824, B1 => n1708, B2 => n35,
                           ZN => n9352);
   U1113 : OAI22_X1 port map( A1 => n1734, A2 => n1824, B1 => n1708, B2 => n37,
                           ZN => n9351);
   U1114 : OAI22_X1 port map( A1 => n1735, A2 => n1824, B1 => n1708, B2 => n39,
                           ZN => n9350);
   U1115 : OAI22_X1 port map( A1 => n1736, A2 => n1824, B1 => n1708, B2 => n41,
                           ZN => n9349);
   U1116 : OAI22_X1 port map( A1 => n1737, A2 => n1824, B1 => n1708, B2 => n43,
                           ZN => n9348);
   U1117 : OAI22_X1 port map( A1 => n1730, A2 => n1824, B1 => n1708, B2 => n45,
                           ZN => n9347);
   U1118 : OAI22_X1 port map( A1 => n1731, A2 => n1824, B1 => n1708, B2 => n47,
                           ZN => n9346);
   U1119 : OAI22_X1 port map( A1 => n1732, A2 => n1824, B1 => n1708, B2 => n49,
                           ZN => n9345);
   U1120 : OAI22_X1 port map( A1 => n1733, A2 => n1824, B1 => n1708, B2 => n51,
                           ZN => n9344);
   U1121 : OAI22_X1 port map( A1 => n1726, A2 => n1824, B1 => n1708, B2 => n53,
                           ZN => n9343);
   U1122 : OAI22_X1 port map( A1 => n1727, A2 => n1824, B1 => n1708, B2 => n55,
                           ZN => n9342);
   U1123 : OAI22_X1 port map( A1 => n1728, A2 => n1824, B1 => n1708, B2 => n57,
                           ZN => n9341);
   U1124 : OAI22_X1 port map( A1 => n1729, A2 => n1824, B1 => n1708, B2 => n59,
                           ZN => n9340);
   U1125 : OAI22_X1 port map( A1 => n1725, A2 => n1824, B1 => n1708, B2 => n61,
                           ZN => n9339);
   U1126 : OAI22_X1 port map( A1 => n1768, A2 => n1824, B1 => n1708, B2 => n63,
                           ZN => n9338);
   U1127 : OAI21_X1 port map( B1 => n1769, B2 => n1824, A => n1770, ZN => n1825
                           );
   U1128 : OAI22_X1 port map( A1 => n1759, A2 => n1826, B1 => n5824, B2 => 
                           n1638, ZN => n9337);
   U1129 : OAI22_X1 port map( A1 => n1761, A2 => n1826, B1 => n5820, B2 => 
                           n1638, ZN => n9336);
   U1130 : OAI22_X1 port map( A1 => n1762, A2 => n1826, B1 => n5816, B2 => 
                           n1638, ZN => n9335);
   U1131 : OAI22_X1 port map( A1 => n1763, A2 => n1826, B1 => n5812, B2 => 
                           n1638, ZN => n9334);
   U1132 : OAI22_X1 port map( A1 => n1764, A2 => n1826, B1 => n5808, B2 => 
                           n1638, ZN => n9333);
   U1133 : OAI22_X1 port map( A1 => n1765, A2 => n1826, B1 => n5804, B2 => 
                           n1638, ZN => n9332);
   U1134 : OAI22_X1 port map( A1 => n1766, A2 => n1826, B1 => n5800, B2 => 
                           n1638, ZN => n9331);
   U1135 : OAI22_X1 port map( A1 => n1767, A2 => n1826, B1 => n5796, B2 => 
                           n1638, ZN => n9330);
   U1136 : OAI22_X1 port map( A1 => n1746, A2 => n1826, B1 => n5792, B2 => 
                           n1638, ZN => n9329);
   U1137 : OAI22_X1 port map( A1 => n1747, A2 => n1826, B1 => n5788, B2 => 
                           n1638, ZN => n9328);
   U1138 : OAI22_X1 port map( A1 => n1742, A2 => n1826, B1 => n5784, B2 => 
                           n1638, ZN => n9327);
   U1139 : OAI22_X1 port map( A1 => n1743, A2 => n1826, B1 => n5780, B2 => 
                           n1638, ZN => n9326);
   U1140 : OAI22_X1 port map( A1 => n1744, A2 => n1826, B1 => n5776, B2 => 
                           n1638, ZN => n9325);
   U1141 : OAI22_X1 port map( A1 => n1745, A2 => n1826, B1 => n5772, B2 => 
                           n1638, ZN => n9324);
   U1142 : OAI22_X1 port map( A1 => n1738, A2 => n1826, B1 => n5768, B2 => 
                           n1638, ZN => n9323);
   U1143 : OAI22_X1 port map( A1 => n1739, A2 => n1826, B1 => n5764, B2 => 
                           n1638, ZN => n9322);
   U1144 : OAI22_X1 port map( A1 => n1740, A2 => n1826, B1 => n5760, B2 => 
                           n1638, ZN => n9321);
   U1145 : OAI22_X1 port map( A1 => n1741, A2 => n1826, B1 => n5756, B2 => 
                           n1638, ZN => n9320);
   U1146 : OAI22_X1 port map( A1 => n1734, A2 => n1826, B1 => n5752, B2 => 
                           n1638, ZN => n9319);
   U1147 : OAI22_X1 port map( A1 => n1735, A2 => n1826, B1 => n5748, B2 => 
                           n1638, ZN => n9318);
   U1148 : OAI22_X1 port map( A1 => n1736, A2 => n1826, B1 => n5744, B2 => 
                           n1638, ZN => n9317);
   U1149 : OAI22_X1 port map( A1 => n1737, A2 => n1826, B1 => n5740, B2 => 
                           n1638, ZN => n9316);
   U1150 : OAI22_X1 port map( A1 => n1730, A2 => n1826, B1 => n5736, B2 => 
                           n1638, ZN => n9315);
   U1151 : OAI22_X1 port map( A1 => n1731, A2 => n1826, B1 => n5732, B2 => 
                           n1638, ZN => n9314);
   U1152 : OAI22_X1 port map( A1 => n1732, A2 => n1826, B1 => n5728, B2 => 
                           n1638, ZN => n9313);
   U1153 : OAI22_X1 port map( A1 => n1733, A2 => n1826, B1 => n5724, B2 => 
                           n1638, ZN => n9312);
   U1154 : OAI22_X1 port map( A1 => n1726, A2 => n1826, B1 => n5720, B2 => 
                           n1638, ZN => n9311);
   U1155 : OAI22_X1 port map( A1 => n1727, A2 => n1826, B1 => n5716, B2 => 
                           n1638, ZN => n9310);
   U1156 : OAI22_X1 port map( A1 => n1728, A2 => n1826, B1 => n5712, B2 => 
                           n1638, ZN => n9309);
   U1157 : OAI22_X1 port map( A1 => n1729, A2 => n1826, B1 => n5708, B2 => 
                           n1638, ZN => n9308);
   U1158 : OAI22_X1 port map( A1 => n1725, A2 => n1826, B1 => n5704, B2 => 
                           n1638, ZN => n9307);
   U1159 : OAI22_X1 port map( A1 => n1768, A2 => n1826, B1 => n5700, B2 => 
                           n1638, ZN => n9306);
   U1160 : OAI21_X1 port map( B1 => n1769, B2 => n1826, A => n1770, ZN => n1827
                           );
   U1161 : OAI22_X1 port map( A1 => n1759, A2 => n1828, B1 => n5825, B2 => 
                           n1640, ZN => n9305);
   U1162 : OAI22_X1 port map( A1 => n1761, A2 => n1828, B1 => n5821, B2 => 
                           n1640, ZN => n9304);
   U1163 : OAI22_X1 port map( A1 => n1762, A2 => n1828, B1 => n5817, B2 => 
                           n1640, ZN => n9303);
   U1164 : OAI22_X1 port map( A1 => n1763, A2 => n1828, B1 => n5813, B2 => 
                           n1640, ZN => n9302);
   U1165 : OAI22_X1 port map( A1 => n1764, A2 => n1828, B1 => n5809, B2 => 
                           n1640, ZN => n9301);
   U1166 : OAI22_X1 port map( A1 => n1765, A2 => n1828, B1 => n5805, B2 => 
                           n1640, ZN => n9300);
   U1167 : OAI22_X1 port map( A1 => n1766, A2 => n1828, B1 => n5801, B2 => 
                           n1640, ZN => n9299);
   U1168 : OAI22_X1 port map( A1 => n1767, A2 => n1828, B1 => n5797, B2 => 
                           n1640, ZN => n9298);
   U1169 : OAI22_X1 port map( A1 => n1746, A2 => n1828, B1 => n5793, B2 => 
                           n1640, ZN => n9297);
   U1170 : OAI22_X1 port map( A1 => n1747, A2 => n1828, B1 => n5789, B2 => 
                           n1640, ZN => n9296);
   U1171 : OAI22_X1 port map( A1 => n1742, A2 => n1828, B1 => n5785, B2 => 
                           n1640, ZN => n9295);
   U1172 : OAI22_X1 port map( A1 => n1743, A2 => n1828, B1 => n5781, B2 => 
                           n1640, ZN => n9294);
   U1173 : OAI22_X1 port map( A1 => n1744, A2 => n1828, B1 => n5777, B2 => 
                           n1640, ZN => n9293);
   U1174 : OAI22_X1 port map( A1 => n1745, A2 => n1828, B1 => n5773, B2 => 
                           n1640, ZN => n9292);
   U1175 : OAI22_X1 port map( A1 => n1738, A2 => n1828, B1 => n5769, B2 => 
                           n1640, ZN => n9291);
   U1176 : OAI22_X1 port map( A1 => n1739, A2 => n1828, B1 => n5765, B2 => 
                           n1640, ZN => n9290);
   U1177 : OAI22_X1 port map( A1 => n1740, A2 => n1828, B1 => n5761, B2 => 
                           n1640, ZN => n9289);
   U1178 : OAI22_X1 port map( A1 => n1741, A2 => n1828, B1 => n5757, B2 => 
                           n1640, ZN => n9288);
   U1179 : OAI22_X1 port map( A1 => n1734, A2 => n1828, B1 => n5753, B2 => 
                           n1640, ZN => n9287);
   U1180 : OAI22_X1 port map( A1 => n1735, A2 => n1828, B1 => n5749, B2 => 
                           n1640, ZN => n9286);
   U1181 : OAI22_X1 port map( A1 => n1736, A2 => n1828, B1 => n5745, B2 => 
                           n1640, ZN => n9285);
   U1182 : OAI22_X1 port map( A1 => n1737, A2 => n1828, B1 => n5741, B2 => 
                           n1640, ZN => n9284);
   U1183 : OAI22_X1 port map( A1 => n1730, A2 => n1828, B1 => n5737, B2 => 
                           n1640, ZN => n9283);
   U1184 : OAI22_X1 port map( A1 => n1731, A2 => n1828, B1 => n5733, B2 => 
                           n1640, ZN => n9282);
   U1185 : OAI22_X1 port map( A1 => n1732, A2 => n1828, B1 => n5729, B2 => 
                           n1640, ZN => n9281);
   U1186 : OAI22_X1 port map( A1 => n1733, A2 => n1828, B1 => n5725, B2 => 
                           n1640, ZN => n9280);
   U1187 : OAI22_X1 port map( A1 => n1726, A2 => n1828, B1 => n5721, B2 => 
                           n1640, ZN => n9279);
   U1188 : OAI22_X1 port map( A1 => n1727, A2 => n1828, B1 => n5717, B2 => 
                           n1640, ZN => n9278);
   U1189 : OAI22_X1 port map( A1 => n1728, A2 => n1828, B1 => n5713, B2 => 
                           n1640, ZN => n9277);
   U1190 : OAI22_X1 port map( A1 => n1729, A2 => n1828, B1 => n5709, B2 => 
                           n1640, ZN => n9276);
   U1191 : OAI22_X1 port map( A1 => n1725, A2 => n1828, B1 => n5705, B2 => 
                           n1640, ZN => n9275);
   U1192 : OAI22_X1 port map( A1 => n1768, A2 => n1828, B1 => n5701, B2 => 
                           n1640, ZN => n9274);
   U1193 : OAI21_X1 port map( B1 => n1769, B2 => n1828, A => n1770, ZN => n1829
                           );
   U1194 : OAI22_X1 port map( A1 => n1759, A2 => n1830, B1 => n1702, B2 => n873
                           , ZN => n9273);
   U1195 : OAI22_X1 port map( A1 => n1761, A2 => n1830, B1 => n1702, B2 => n874
                           , ZN => n9272);
   U1196 : OAI22_X1 port map( A1 => n1762, A2 => n1830, B1 => n1702, B2 => n875
                           , ZN => n9271);
   U1197 : OAI22_X1 port map( A1 => n1763, A2 => n1830, B1 => n1702, B2 => n876
                           , ZN => n9270);
   U1198 : OAI22_X1 port map( A1 => n1764, A2 => n1830, B1 => n1702, B2 => n877
                           , ZN => n9269);
   U1199 : OAI22_X1 port map( A1 => n1765, A2 => n1830, B1 => n1702, B2 => n878
                           , ZN => n9268);
   U1200 : OAI22_X1 port map( A1 => n1766, A2 => n1830, B1 => n1702, B2 => n879
                           , ZN => n9267);
   U1201 : OAI22_X1 port map( A1 => n1767, A2 => n1830, B1 => n1702, B2 => n880
                           , ZN => n9266);
   U1202 : OAI22_X1 port map( A1 => n1746, A2 => n1830, B1 => n1702, B2 => n881
                           , ZN => n9265);
   U1203 : OAI22_X1 port map( A1 => n1747, A2 => n1830, B1 => n1702, B2 => n882
                           , ZN => n9264);
   U1204 : OAI22_X1 port map( A1 => n1742, A2 => n1830, B1 => n1702, B2 => n883
                           , ZN => n9263);
   U1205 : OAI22_X1 port map( A1 => n1743, A2 => n1830, B1 => n1702, B2 => n884
                           , ZN => n9262);
   U1206 : OAI22_X1 port map( A1 => n1744, A2 => n1830, B1 => n1702, B2 => n885
                           , ZN => n9261);
   U1207 : OAI22_X1 port map( A1 => n1745, A2 => n1830, B1 => n1702, B2 => n886
                           , ZN => n9260);
   U1208 : OAI22_X1 port map( A1 => n1738, A2 => n1830, B1 => n1702, B2 => n887
                           , ZN => n9259);
   U1209 : OAI22_X1 port map( A1 => n1739, A2 => n1830, B1 => n1702, B2 => n888
                           , ZN => n9258);
   U1210 : OAI22_X1 port map( A1 => n1740, A2 => n1830, B1 => n1702, B2 => n889
                           , ZN => n9257);
   U1211 : OAI22_X1 port map( A1 => n1741, A2 => n1830, B1 => n1702, B2 => n890
                           , ZN => n9256);
   U1212 : OAI22_X1 port map( A1 => n1734, A2 => n1830, B1 => n1702, B2 => n891
                           , ZN => n9255);
   U1213 : OAI22_X1 port map( A1 => n1735, A2 => n1830, B1 => n1702, B2 => n892
                           , ZN => n9254);
   U1214 : OAI22_X1 port map( A1 => n1736, A2 => n1830, B1 => n1702, B2 => n893
                           , ZN => n9253);
   U1215 : OAI22_X1 port map( A1 => n1737, A2 => n1830, B1 => n1702, B2 => n894
                           , ZN => n9252);
   U1216 : OAI22_X1 port map( A1 => n1730, A2 => n1830, B1 => n1702, B2 => n895
                           , ZN => n9251);
   U1217 : OAI22_X1 port map( A1 => n1731, A2 => n1830, B1 => n1702, B2 => n896
                           , ZN => n9250);
   U1218 : OAI22_X1 port map( A1 => n1732, A2 => n1830, B1 => n1702, B2 => n897
                           , ZN => n9249);
   U1219 : OAI22_X1 port map( A1 => n1733, A2 => n1830, B1 => n1702, B2 => n898
                           , ZN => n9248);
   U1220 : OAI22_X1 port map( A1 => n1726, A2 => n1830, B1 => n1702, B2 => n899
                           , ZN => n9247);
   U1221 : OAI22_X1 port map( A1 => n1727, A2 => n1830, B1 => n1702, B2 => n900
                           , ZN => n9246);
   U1222 : OAI22_X1 port map( A1 => n1728, A2 => n1830, B1 => n1702, B2 => n901
                           , ZN => n9245);
   U1223 : OAI22_X1 port map( A1 => n1729, A2 => n1830, B1 => n1702, B2 => n902
                           , ZN => n9244);
   U1224 : OAI22_X1 port map( A1 => n1725, A2 => n1830, B1 => n1702, B2 => n903
                           , ZN => n9243);
   U1225 : OAI22_X1 port map( A1 => n1768, A2 => n1830, B1 => n1702, B2 => n904
                           , ZN => n9242);
   U1226 : OAI21_X1 port map( B1 => n1769, B2 => n1830, A => n1770, ZN => n1831
                           );
   U1227 : OAI22_X1 port map( A1 => n1759, A2 => n1832, B1 => n1704, B2 => 
                           n1225, ZN => n9241);
   U1228 : OAI22_X1 port map( A1 => n1761, A2 => n1832, B1 => n1704, B2 => 
                           n1226, ZN => n9240);
   U1229 : OAI22_X1 port map( A1 => n1762, A2 => n1832, B1 => n1704, B2 => 
                           n1227, ZN => n9239);
   U1230 : OAI22_X1 port map( A1 => n1763, A2 => n1832, B1 => n1704, B2 => 
                           n1228, ZN => n9238);
   U1231 : OAI22_X1 port map( A1 => n1764, A2 => n1832, B1 => n1704, B2 => 
                           n1229, ZN => n9237);
   U1232 : OAI22_X1 port map( A1 => n1765, A2 => n1832, B1 => n1704, B2 => 
                           n1230, ZN => n9236);
   U1233 : OAI22_X1 port map( A1 => n1766, A2 => n1832, B1 => n1704, B2 => 
                           n1231, ZN => n9235);
   U1234 : OAI22_X1 port map( A1 => n1767, A2 => n1832, B1 => n1704, B2 => 
                           n1232, ZN => n9234);
   U1235 : OAI22_X1 port map( A1 => n1746, A2 => n1832, B1 => n1704, B2 => 
                           n1233, ZN => n9233);
   U1236 : OAI22_X1 port map( A1 => n1747, A2 => n1832, B1 => n1704, B2 => 
                           n1234, ZN => n9232);
   U1237 : OAI22_X1 port map( A1 => n1742, A2 => n1832, B1 => n1704, B2 => 
                           n1235, ZN => n9231);
   U1238 : OAI22_X1 port map( A1 => n1743, A2 => n1832, B1 => n1704, B2 => 
                           n1236, ZN => n9230);
   U1239 : OAI22_X1 port map( A1 => n1744, A2 => n1832, B1 => n1704, B2 => 
                           n1237, ZN => n9229);
   U1240 : OAI22_X1 port map( A1 => n1745, A2 => n1832, B1 => n1704, B2 => 
                           n1238, ZN => n9228);
   U1241 : OAI22_X1 port map( A1 => n1738, A2 => n1832, B1 => n1704, B2 => 
                           n1239, ZN => n9227);
   U1242 : OAI22_X1 port map( A1 => n1739, A2 => n1832, B1 => n1704, B2 => 
                           n1240, ZN => n9226);
   U1243 : OAI22_X1 port map( A1 => n1740, A2 => n1832, B1 => n1704, B2 => 
                           n1241, ZN => n9225);
   U1244 : OAI22_X1 port map( A1 => n1741, A2 => n1832, B1 => n1704, B2 => 
                           n1242, ZN => n9224);
   U1245 : OAI22_X1 port map( A1 => n1734, A2 => n1832, B1 => n1704, B2 => 
                           n1243, ZN => n9223);
   U1246 : OAI22_X1 port map( A1 => n1735, A2 => n1832, B1 => n1704, B2 => 
                           n1244, ZN => n9222);
   U1247 : OAI22_X1 port map( A1 => n1736, A2 => n1832, B1 => n1704, B2 => 
                           n1245, ZN => n9221);
   U1248 : OAI22_X1 port map( A1 => n1737, A2 => n1832, B1 => n1704, B2 => 
                           n1246, ZN => n9220);
   U1249 : OAI22_X1 port map( A1 => n1730, A2 => n1832, B1 => n1704, B2 => 
                           n1247, ZN => n9219);
   U1250 : OAI22_X1 port map( A1 => n1731, A2 => n1832, B1 => n1704, B2 => 
                           n1248, ZN => n9218);
   U1251 : OAI22_X1 port map( A1 => n1732, A2 => n1832, B1 => n1704, B2 => 
                           n1249, ZN => n9217);
   U1252 : OAI22_X1 port map( A1 => n1733, A2 => n1832, B1 => n1704, B2 => 
                           n1250, ZN => n9216);
   U1253 : OAI22_X1 port map( A1 => n1726, A2 => n1832, B1 => n1704, B2 => 
                           n1251, ZN => n9215);
   U1254 : OAI22_X1 port map( A1 => n1727, A2 => n1832, B1 => n1704, B2 => 
                           n1252, ZN => n9214);
   U1255 : OAI22_X1 port map( A1 => n1728, A2 => n1832, B1 => n1704, B2 => 
                           n1253, ZN => n9213);
   U1256 : OAI22_X1 port map( A1 => n1729, A2 => n1832, B1 => n1704, B2 => 
                           n1254, ZN => n9212);
   U1257 : OAI22_X1 port map( A1 => n1725, A2 => n1832, B1 => n1704, B2 => 
                           n1255, ZN => n9211);
   U1258 : OAI22_X1 port map( A1 => n1768, A2 => n1832, B1 => n1704, B2 => 
                           n1256, ZN => n9210);
   U1259 : OAI21_X1 port map( B1 => n1769, B2 => n1832, A => n1770, ZN => n1833
                           );
   U1260 : OAI22_X1 port map( A1 => n1759, A2 => n1834, B1 => n5185, B2 => 
                           n1634, ZN => n9209);
   U1261 : OAI22_X1 port map( A1 => n1761, A2 => n1834, B1 => n5184, B2 => 
                           n1634, ZN => n9208);
   U1262 : OAI22_X1 port map( A1 => n1762, A2 => n1834, B1 => n5183, B2 => 
                           n1634, ZN => n9207);
   U1263 : OAI22_X1 port map( A1 => n1763, A2 => n1834, B1 => n5182, B2 => 
                           n1634, ZN => n9206);
   U1264 : OAI22_X1 port map( A1 => n1764, A2 => n1834, B1 => n5181, B2 => 
                           n1634, ZN => n9205);
   U1265 : OAI22_X1 port map( A1 => n1765, A2 => n1834, B1 => n5180, B2 => 
                           n1634, ZN => n9204);
   U1266 : OAI22_X1 port map( A1 => n1766, A2 => n1834, B1 => n5179, B2 => 
                           n1634, ZN => n9203);
   U1267 : OAI22_X1 port map( A1 => n1767, A2 => n1834, B1 => n5178, B2 => 
                           n1634, ZN => n9202);
   U1268 : OAI22_X1 port map( A1 => n1746, A2 => n1834, B1 => n5177, B2 => 
                           n1634, ZN => n9201);
   U1269 : OAI22_X1 port map( A1 => n1747, A2 => n1834, B1 => n5176, B2 => 
                           n1634, ZN => n9200);
   U1270 : OAI22_X1 port map( A1 => n1742, A2 => n1834, B1 => n5175, B2 => 
                           n1634, ZN => n9199);
   U1271 : OAI22_X1 port map( A1 => n1743, A2 => n1834, B1 => n5174, B2 => 
                           n1634, ZN => n9198);
   U1272 : OAI22_X1 port map( A1 => n1744, A2 => n1834, B1 => n5173, B2 => 
                           n1634, ZN => n9197);
   U1273 : OAI22_X1 port map( A1 => n1745, A2 => n1834, B1 => n5172, B2 => 
                           n1634, ZN => n9196);
   U1274 : OAI22_X1 port map( A1 => n1738, A2 => n1834, B1 => n5171, B2 => 
                           n1634, ZN => n9195);
   U1275 : OAI22_X1 port map( A1 => n1739, A2 => n1834, B1 => n5170, B2 => 
                           n1634, ZN => n9194);
   U1276 : OAI22_X1 port map( A1 => n1740, A2 => n1834, B1 => n5169, B2 => 
                           n1634, ZN => n9193);
   U1277 : OAI22_X1 port map( A1 => n1741, A2 => n1834, B1 => n5168, B2 => 
                           n1634, ZN => n9192);
   U1278 : OAI22_X1 port map( A1 => n1734, A2 => n1834, B1 => n5167, B2 => 
                           n1634, ZN => n9191);
   U1279 : OAI22_X1 port map( A1 => n1735, A2 => n1834, B1 => n5166, B2 => 
                           n1634, ZN => n9190);
   U1280 : OAI22_X1 port map( A1 => n1736, A2 => n1834, B1 => n5165, B2 => 
                           n1634, ZN => n9189);
   U1281 : OAI22_X1 port map( A1 => n1737, A2 => n1834, B1 => n5164, B2 => 
                           n1634, ZN => n9188);
   U1282 : OAI22_X1 port map( A1 => n1730, A2 => n1834, B1 => n5163, B2 => 
                           n1634, ZN => n9187);
   U1283 : OAI22_X1 port map( A1 => n1731, A2 => n1834, B1 => n5162, B2 => 
                           n1634, ZN => n9186);
   U1284 : OAI22_X1 port map( A1 => n1732, A2 => n1834, B1 => n5161, B2 => 
                           n1634, ZN => n9185);
   U1285 : OAI22_X1 port map( A1 => n1733, A2 => n1834, B1 => n5160, B2 => 
                           n1634, ZN => n9184);
   U1286 : OAI22_X1 port map( A1 => n1726, A2 => n1834, B1 => n5159, B2 => 
                           n1634, ZN => n9183);
   U1287 : OAI22_X1 port map( A1 => n1727, A2 => n1834, B1 => n5158, B2 => 
                           n1634, ZN => n9182);
   U1288 : OAI22_X1 port map( A1 => n1728, A2 => n1834, B1 => n5157, B2 => 
                           n1634, ZN => n9181);
   U1289 : OAI22_X1 port map( A1 => n1729, A2 => n1834, B1 => n5156, B2 => 
                           n1634, ZN => n9180);
   U1290 : OAI22_X1 port map( A1 => n1725, A2 => n1834, B1 => n5155, B2 => 
                           n1634, ZN => n9179);
   U1291 : OAI22_X1 port map( A1 => n1768, A2 => n1834, B1 => n5154, B2 => 
                           n1634, ZN => n9178);
   U1292 : OAI21_X1 port map( B1 => n1769, B2 => n1834, A => n1770, ZN => n1835
                           );
   U1293 : OAI22_X1 port map( A1 => n1759, A2 => n1836, B1 => n5153, B2 => 
                           n1636, ZN => n9177);
   U1294 : OAI22_X1 port map( A1 => n1761, A2 => n1836, B1 => n5152, B2 => 
                           n1636, ZN => n9176);
   U1295 : OAI22_X1 port map( A1 => n1762, A2 => n1836, B1 => n5151, B2 => 
                           n1636, ZN => n9175);
   U1296 : OAI22_X1 port map( A1 => n1763, A2 => n1836, B1 => n5150, B2 => 
                           n1636, ZN => n9174);
   U1297 : OAI22_X1 port map( A1 => n1764, A2 => n1836, B1 => n5149, B2 => 
                           n1636, ZN => n9173);
   U1298 : OAI22_X1 port map( A1 => n1765, A2 => n1836, B1 => n5148, B2 => 
                           n1636, ZN => n9172);
   U1299 : OAI22_X1 port map( A1 => n1766, A2 => n1836, B1 => n5147, B2 => 
                           n1636, ZN => n9171);
   U1300 : OAI22_X1 port map( A1 => n1767, A2 => n1836, B1 => n5146, B2 => 
                           n1636, ZN => n9170);
   U1301 : OAI22_X1 port map( A1 => n1746, A2 => n1836, B1 => n5145, B2 => 
                           n1636, ZN => n9169);
   U1302 : OAI22_X1 port map( A1 => n1747, A2 => n1836, B1 => n5144, B2 => 
                           n1636, ZN => n9168);
   U1303 : OAI22_X1 port map( A1 => n1742, A2 => n1836, B1 => n5143, B2 => 
                           n1636, ZN => n9167);
   U1304 : OAI22_X1 port map( A1 => n1743, A2 => n1836, B1 => n5142, B2 => 
                           n1636, ZN => n9166);
   U1305 : OAI22_X1 port map( A1 => n1744, A2 => n1836, B1 => n5141, B2 => 
                           n1636, ZN => n9165);
   U1306 : OAI22_X1 port map( A1 => n1745, A2 => n1836, B1 => n5140, B2 => 
                           n1636, ZN => n9164);
   U1307 : OAI22_X1 port map( A1 => n1738, A2 => n1836, B1 => n5139, B2 => 
                           n1636, ZN => n9163);
   U1308 : OAI22_X1 port map( A1 => n1739, A2 => n1836, B1 => n5138, B2 => 
                           n1636, ZN => n9162);
   U1309 : OAI22_X1 port map( A1 => n1740, A2 => n1836, B1 => n5137, B2 => 
                           n1636, ZN => n9161);
   U1310 : OAI22_X1 port map( A1 => n1741, A2 => n1836, B1 => n5136, B2 => 
                           n1636, ZN => n9160);
   U1311 : OAI22_X1 port map( A1 => n1734, A2 => n1836, B1 => n5135, B2 => 
                           n1636, ZN => n9159);
   U1312 : OAI22_X1 port map( A1 => n1735, A2 => n1836, B1 => n5134, B2 => 
                           n1636, ZN => n9158);
   U1313 : OAI22_X1 port map( A1 => n1736, A2 => n1836, B1 => n5133, B2 => 
                           n1636, ZN => n9157);
   U1314 : OAI22_X1 port map( A1 => n1737, A2 => n1836, B1 => n5132, B2 => 
                           n1636, ZN => n9156);
   U1315 : OAI22_X1 port map( A1 => n1730, A2 => n1836, B1 => n5131, B2 => 
                           n1636, ZN => n9155);
   U1316 : OAI22_X1 port map( A1 => n1731, A2 => n1836, B1 => n5130, B2 => 
                           n1636, ZN => n9154);
   U1317 : OAI22_X1 port map( A1 => n1732, A2 => n1836, B1 => n5129, B2 => 
                           n1636, ZN => n9153);
   U1318 : OAI22_X1 port map( A1 => n1733, A2 => n1836, B1 => n5128, B2 => 
                           n1636, ZN => n9152);
   U1319 : OAI22_X1 port map( A1 => n1726, A2 => n1836, B1 => n5127, B2 => 
                           n1636, ZN => n9151);
   U1320 : OAI22_X1 port map( A1 => n1727, A2 => n1836, B1 => n5126, B2 => 
                           n1636, ZN => n9150);
   U1321 : OAI22_X1 port map( A1 => n1728, A2 => n1836, B1 => n5125, B2 => 
                           n1636, ZN => n9149);
   U1322 : OAI22_X1 port map( A1 => n1729, A2 => n1836, B1 => n5124, B2 => 
                           n1636, ZN => n9148);
   U1323 : OAI22_X1 port map( A1 => n1725, A2 => n1836, B1 => n5123, B2 => 
                           n1636, ZN => n9147);
   U1324 : OAI22_X1 port map( A1 => n1768, A2 => n1836, B1 => n5122, B2 => 
                           n1636, ZN => n9146);
   U1325 : OAI21_X1 port map( B1 => n1769, B2 => n1836, A => n1770, ZN => n1837
                           );
   U1326 : OAI22_X1 port map( A1 => n1759, A2 => n1838, B1 => n5121, B2 => 
                           n1630, ZN => n9145);
   U1327 : OAI22_X1 port map( A1 => n1761, A2 => n1838, B1 => n5120, B2 => 
                           n1630, ZN => n9144);
   U1328 : OAI22_X1 port map( A1 => n1762, A2 => n1838, B1 => n5119, B2 => 
                           n1630, ZN => n9143);
   U1329 : OAI22_X1 port map( A1 => n1763, A2 => n1838, B1 => n5118, B2 => 
                           n1630, ZN => n9142);
   U1330 : OAI22_X1 port map( A1 => n1764, A2 => n1838, B1 => n5117, B2 => 
                           n1630, ZN => n9141);
   U1331 : OAI22_X1 port map( A1 => n1765, A2 => n1838, B1 => n5116, B2 => 
                           n1630, ZN => n9140);
   U1332 : OAI22_X1 port map( A1 => n1766, A2 => n1838, B1 => n5115, B2 => 
                           n1630, ZN => n9139);
   U1333 : OAI22_X1 port map( A1 => n1767, A2 => n1838, B1 => n5114, B2 => 
                           n1630, ZN => n9138);
   U1334 : OAI22_X1 port map( A1 => n1746, A2 => n1838, B1 => n5113, B2 => 
                           n1630, ZN => n9137);
   U1335 : OAI22_X1 port map( A1 => n1747, A2 => n1838, B1 => n5112, B2 => 
                           n1630, ZN => n9136);
   U1336 : OAI22_X1 port map( A1 => n1742, A2 => n1838, B1 => n5111, B2 => 
                           n1630, ZN => n9135);
   U1337 : OAI22_X1 port map( A1 => n1743, A2 => n1838, B1 => n5110, B2 => 
                           n1630, ZN => n9134);
   U1338 : OAI22_X1 port map( A1 => n1744, A2 => n1838, B1 => n5109, B2 => 
                           n1630, ZN => n9133);
   U1339 : OAI22_X1 port map( A1 => n1745, A2 => n1838, B1 => n5108, B2 => 
                           n1630, ZN => n9132);
   U1340 : OAI22_X1 port map( A1 => n1738, A2 => n1838, B1 => n5107, B2 => 
                           n1630, ZN => n9131);
   U1341 : OAI22_X1 port map( A1 => n1739, A2 => n1838, B1 => n5106, B2 => 
                           n1630, ZN => n9130);
   U1342 : OAI22_X1 port map( A1 => n1740, A2 => n1838, B1 => n5105, B2 => 
                           n1630, ZN => n9129);
   U1343 : OAI22_X1 port map( A1 => n1741, A2 => n1838, B1 => n5104, B2 => 
                           n1630, ZN => n9128);
   U1344 : OAI22_X1 port map( A1 => n1734, A2 => n1838, B1 => n5103, B2 => 
                           n1630, ZN => n9127);
   U1345 : OAI22_X1 port map( A1 => n1735, A2 => n1838, B1 => n5102, B2 => 
                           n1630, ZN => n9126);
   U1346 : OAI22_X1 port map( A1 => n1736, A2 => n1838, B1 => n5101, B2 => 
                           n1630, ZN => n9125);
   U1347 : OAI22_X1 port map( A1 => n1737, A2 => n1838, B1 => n5100, B2 => 
                           n1630, ZN => n9124);
   U1348 : OAI22_X1 port map( A1 => n1730, A2 => n1838, B1 => n5099, B2 => 
                           n1630, ZN => n9123);
   U1349 : OAI22_X1 port map( A1 => n1731, A2 => n1838, B1 => n5098, B2 => 
                           n1630, ZN => n9122);
   U1350 : OAI22_X1 port map( A1 => n1732, A2 => n1838, B1 => n5097, B2 => 
                           n1630, ZN => n9121);
   U1351 : OAI22_X1 port map( A1 => n1733, A2 => n1838, B1 => n5096, B2 => 
                           n1630, ZN => n9120);
   U1352 : OAI22_X1 port map( A1 => n1726, A2 => n1838, B1 => n5095, B2 => 
                           n1630, ZN => n9119);
   U1353 : OAI22_X1 port map( A1 => n1727, A2 => n1838, B1 => n5094, B2 => 
                           n1630, ZN => n9118);
   U1354 : OAI22_X1 port map( A1 => n1728, A2 => n1838, B1 => n5093, B2 => 
                           n1630, ZN => n9117);
   U1355 : OAI22_X1 port map( A1 => n1729, A2 => n1838, B1 => n5092, B2 => 
                           n1630, ZN => n9116);
   U1356 : OAI22_X1 port map( A1 => n1725, A2 => n1838, B1 => n5091, B2 => 
                           n1630, ZN => n9115);
   U1357 : OAI22_X1 port map( A1 => n1768, A2 => n1838, B1 => n5090, B2 => 
                           n1630, ZN => n9114);
   U1358 : OAI21_X1 port map( B1 => n1769, B2 => n1838, A => n1770, ZN => n1839
                           );
   U1359 : OAI22_X1 port map( A1 => n1759, A2 => n1840, B1 => n1698, B2 => n65,
                           ZN => n9113);
   U1360 : OAI22_X1 port map( A1 => n1761, A2 => n1840, B1 => n1698, B2 => n66,
                           ZN => n9112);
   U1361 : OAI22_X1 port map( A1 => n1762, A2 => n1840, B1 => n1698, B2 => n67,
                           ZN => n9111);
   U1362 : OAI22_X1 port map( A1 => n1763, A2 => n1840, B1 => n1698, B2 => n68,
                           ZN => n9110);
   U1363 : OAI22_X1 port map( A1 => n1764, A2 => n1840, B1 => n1698, B2 => n69,
                           ZN => n9109);
   U1364 : OAI22_X1 port map( A1 => n1765, A2 => n1840, B1 => n1698, B2 => n70,
                           ZN => n9108);
   U1365 : OAI22_X1 port map( A1 => n1766, A2 => n1840, B1 => n1698, B2 => n71,
                           ZN => n9107);
   U1366 : OAI22_X1 port map( A1 => n1767, A2 => n1840, B1 => n1698, B2 => n72,
                           ZN => n9106);
   U1367 : OAI22_X1 port map( A1 => n1746, A2 => n1840, B1 => n1698, B2 => n73,
                           ZN => n9105);
   U1368 : OAI22_X1 port map( A1 => n1747, A2 => n1840, B1 => n1698, B2 => n74,
                           ZN => n9104);
   U1369 : OAI22_X1 port map( A1 => n1742, A2 => n1840, B1 => n1698, B2 => n75,
                           ZN => n9103);
   U1370 : OAI22_X1 port map( A1 => n1743, A2 => n1840, B1 => n1698, B2 => n76,
                           ZN => n9102);
   U1371 : OAI22_X1 port map( A1 => n1744, A2 => n1840, B1 => n1698, B2 => n77,
                           ZN => n9101);
   U1372 : OAI22_X1 port map( A1 => n1745, A2 => n1840, B1 => n1698, B2 => n78,
                           ZN => n9100);
   U1373 : OAI22_X1 port map( A1 => n1738, A2 => n1840, B1 => n1698, B2 => n79,
                           ZN => n9099);
   U1374 : OAI22_X1 port map( A1 => n1739, A2 => n1840, B1 => n1698, B2 => n80,
                           ZN => n9098);
   U1375 : OAI22_X1 port map( A1 => n1740, A2 => n1840, B1 => n1698, B2 => n81,
                           ZN => n9097);
   U1376 : OAI22_X1 port map( A1 => n1741, A2 => n1840, B1 => n1698, B2 => n82,
                           ZN => n9096);
   U1377 : OAI22_X1 port map( A1 => n1734, A2 => n1840, B1 => n1698, B2 => n83,
                           ZN => n9095);
   U1378 : OAI22_X1 port map( A1 => n1735, A2 => n1840, B1 => n1698, B2 => n84,
                           ZN => n9094);
   U1379 : OAI22_X1 port map( A1 => n1736, A2 => n1840, B1 => n1698, B2 => n85,
                           ZN => n9093);
   U1380 : OAI22_X1 port map( A1 => n1737, A2 => n1840, B1 => n1698, B2 => n86,
                           ZN => n9092);
   U1381 : OAI22_X1 port map( A1 => n1730, A2 => n1840, B1 => n1698, B2 => n87,
                           ZN => n9091);
   U1382 : OAI22_X1 port map( A1 => n1731, A2 => n1840, B1 => n1698, B2 => n88,
                           ZN => n9090);
   U1383 : OAI22_X1 port map( A1 => n1732, A2 => n1840, B1 => n1698, B2 => n89,
                           ZN => n9089);
   U1384 : OAI22_X1 port map( A1 => n1733, A2 => n1840, B1 => n1698, B2 => n90,
                           ZN => n9088);
   U1385 : OAI22_X1 port map( A1 => n1726, A2 => n1840, B1 => n1698, B2 => n91,
                           ZN => n9087);
   U1386 : OAI22_X1 port map( A1 => n1727, A2 => n1840, B1 => n1698, B2 => n92,
                           ZN => n9086);
   U1387 : OAI22_X1 port map( A1 => n1728, A2 => n1840, B1 => n1698, B2 => n93,
                           ZN => n9085);
   U1388 : OAI22_X1 port map( A1 => n1729, A2 => n1840, B1 => n1698, B2 => n94,
                           ZN => n9084);
   U1389 : OAI22_X1 port map( A1 => n1725, A2 => n1840, B1 => n1698, B2 => n95,
                           ZN => n9083);
   U1390 : OAI22_X1 port map( A1 => n1768, A2 => n1840, B1 => n1698, B2 => n96,
                           ZN => n9082);
   U1391 : OAI21_X1 port map( B1 => n1769, B2 => n1840, A => n1770, ZN => n1841
                           );
   U1392 : OAI22_X1 port map( A1 => n1759, A2 => n1842, B1 => n1700, B2 => n425
                           , ZN => n9081);
   U1393 : OAI22_X1 port map( A1 => n1761, A2 => n1842, B1 => n1700, B2 => n426
                           , ZN => n9080);
   U1394 : OAI22_X1 port map( A1 => n1762, A2 => n1842, B1 => n1700, B2 => n427
                           , ZN => n9079);
   U1395 : OAI22_X1 port map( A1 => n1763, A2 => n1842, B1 => n1700, B2 => n428
                           , ZN => n9078);
   U1396 : OAI22_X1 port map( A1 => n1764, A2 => n1842, B1 => n1700, B2 => n429
                           , ZN => n9077);
   U1397 : OAI22_X1 port map( A1 => n1765, A2 => n1842, B1 => n1700, B2 => n430
                           , ZN => n9076);
   U1398 : OAI22_X1 port map( A1 => n1766, A2 => n1842, B1 => n1700, B2 => n431
                           , ZN => n9075);
   U1399 : OAI22_X1 port map( A1 => n1767, A2 => n1842, B1 => n1700, B2 => n432
                           , ZN => n9074);
   U1400 : OAI22_X1 port map( A1 => n1746, A2 => n1842, B1 => n1700, B2 => n433
                           , ZN => n9073);
   U1401 : OAI22_X1 port map( A1 => n1747, A2 => n1842, B1 => n1700, B2 => n434
                           , ZN => n9072);
   U1402 : OAI22_X1 port map( A1 => n1742, A2 => n1842, B1 => n1700, B2 => n435
                           , ZN => n9071);
   U1403 : OAI22_X1 port map( A1 => n1743, A2 => n1842, B1 => n1700, B2 => n436
                           , ZN => n9070);
   U1404 : OAI22_X1 port map( A1 => n1744, A2 => n1842, B1 => n1700, B2 => n437
                           , ZN => n9069);
   U1405 : OAI22_X1 port map( A1 => n1745, A2 => n1842, B1 => n1700, B2 => n438
                           , ZN => n9068);
   U1406 : OAI22_X1 port map( A1 => n1738, A2 => n1842, B1 => n1700, B2 => n439
                           , ZN => n9067);
   U1407 : OAI22_X1 port map( A1 => n1739, A2 => n1842, B1 => n1700, B2 => n440
                           , ZN => n9066);
   U1408 : OAI22_X1 port map( A1 => n1740, A2 => n1842, B1 => n1700, B2 => n441
                           , ZN => n9065);
   U1409 : OAI22_X1 port map( A1 => n1741, A2 => n1842, B1 => n1700, B2 => n442
                           , ZN => n9064);
   U1410 : OAI22_X1 port map( A1 => n1734, A2 => n1842, B1 => n1700, B2 => n443
                           , ZN => n9063);
   U1411 : OAI22_X1 port map( A1 => n1735, A2 => n1842, B1 => n1700, B2 => n444
                           , ZN => n9062);
   U1412 : OAI22_X1 port map( A1 => n1736, A2 => n1842, B1 => n1700, B2 => n445
                           , ZN => n9061);
   U1413 : OAI22_X1 port map( A1 => n1737, A2 => n1842, B1 => n1700, B2 => n446
                           , ZN => n9060);
   U1414 : OAI22_X1 port map( A1 => n1730, A2 => n1842, B1 => n1700, B2 => n447
                           , ZN => n9059);
   U1415 : OAI22_X1 port map( A1 => n1731, A2 => n1842, B1 => n1700, B2 => n448
                           , ZN => n9058);
   U1416 : OAI22_X1 port map( A1 => n1732, A2 => n1842, B1 => n1700, B2 => n449
                           , ZN => n9057);
   U1417 : OAI22_X1 port map( A1 => n1733, A2 => n1842, B1 => n1700, B2 => n450
                           , ZN => n9056);
   U1418 : OAI22_X1 port map( A1 => n1726, A2 => n1842, B1 => n1700, B2 => n451
                           , ZN => n9055);
   U1419 : OAI22_X1 port map( A1 => n1727, A2 => n1842, B1 => n1700, B2 => n452
                           , ZN => n9054);
   U1420 : OAI22_X1 port map( A1 => n1728, A2 => n1842, B1 => n1700, B2 => n453
                           , ZN => n9053);
   U1421 : OAI22_X1 port map( A1 => n1729, A2 => n1842, B1 => n1700, B2 => n454
                           , ZN => n9052);
   U1422 : OAI22_X1 port map( A1 => n1725, A2 => n1842, B1 => n1700, B2 => n455
                           , ZN => n9051);
   U1423 : OAI22_X1 port map( A1 => n1768, A2 => n1842, B1 => n1700, B2 => n456
                           , ZN => n9050);
   U1424 : OAI21_X1 port map( B1 => n1769, B2 => n1842, A => n1770, ZN => n1843
                           );
   U1425 : OAI22_X1 port map( A1 => n1759, A2 => n1844, B1 => n5692, B2 => 
                           n1632, ZN => n9049);
   U1426 : OAI22_X1 port map( A1 => n1761, A2 => n1844, B1 => n5682, B2 => 
                           n1632, ZN => n9048);
   U1427 : OAI22_X1 port map( A1 => n1762, A2 => n1844, B1 => n5672, B2 => 
                           n1632, ZN => n9047);
   U1428 : OAI22_X1 port map( A1 => n1763, A2 => n1844, B1 => n5662, B2 => 
                           n1632, ZN => n9046);
   U1429 : OAI22_X1 port map( A1 => n1764, A2 => n1844, B1 => n5652, B2 => 
                           n1632, ZN => n9045);
   U1430 : OAI22_X1 port map( A1 => n1765, A2 => n1844, B1 => n5642, B2 => 
                           n1632, ZN => n9044);
   U1431 : OAI22_X1 port map( A1 => n1766, A2 => n1844, B1 => n5632, B2 => 
                           n1632, ZN => n9043);
   U1432 : OAI22_X1 port map( A1 => n1767, A2 => n1844, B1 => n5622, B2 => 
                           n1632, ZN => n9042);
   U1433 : OAI22_X1 port map( A1 => n1746, A2 => n1844, B1 => n5612, B2 => 
                           n1632, ZN => n9041);
   U1434 : OAI22_X1 port map( A1 => n1747, A2 => n1844, B1 => n5602, B2 => 
                           n1632, ZN => n9040);
   U1435 : OAI22_X1 port map( A1 => n1742, A2 => n1844, B1 => n5592, B2 => 
                           n1632, ZN => n9039);
   U1436 : OAI22_X1 port map( A1 => n1743, A2 => n1844, B1 => n5582, B2 => 
                           n1632, ZN => n9038);
   U1437 : OAI22_X1 port map( A1 => n1744, A2 => n1844, B1 => n5572, B2 => 
                           n1632, ZN => n9037);
   U1438 : OAI22_X1 port map( A1 => n1745, A2 => n1844, B1 => n5562, B2 => 
                           n1632, ZN => n9036);
   U1439 : OAI22_X1 port map( A1 => n1738, A2 => n1844, B1 => n5552, B2 => 
                           n1632, ZN => n9035);
   U1440 : OAI22_X1 port map( A1 => n1739, A2 => n1844, B1 => n5542, B2 => 
                           n1632, ZN => n9034);
   U1441 : OAI22_X1 port map( A1 => n1740, A2 => n1844, B1 => n5532, B2 => 
                           n1632, ZN => n9033);
   U1442 : OAI22_X1 port map( A1 => n1741, A2 => n1844, B1 => n5522, B2 => 
                           n1632, ZN => n9032);
   U1443 : OAI22_X1 port map( A1 => n1734, A2 => n1844, B1 => n5512, B2 => 
                           n1632, ZN => n9031);
   U1444 : OAI22_X1 port map( A1 => n1735, A2 => n1844, B1 => n5502, B2 => 
                           n1632, ZN => n9030);
   U1445 : OAI22_X1 port map( A1 => n1736, A2 => n1844, B1 => n5492, B2 => 
                           n1632, ZN => n9029);
   U1446 : OAI22_X1 port map( A1 => n1737, A2 => n1844, B1 => n5482, B2 => 
                           n1632, ZN => n9028);
   U1447 : OAI22_X1 port map( A1 => n1730, A2 => n1844, B1 => n5472, B2 => 
                           n1632, ZN => n9027);
   U1448 : OAI22_X1 port map( A1 => n1731, A2 => n1844, B1 => n5462, B2 => 
                           n1632, ZN => n9026);
   U1449 : OAI22_X1 port map( A1 => n1732, A2 => n1844, B1 => n5452, B2 => 
                           n1632, ZN => n9025);
   U1450 : OAI22_X1 port map( A1 => n1733, A2 => n1844, B1 => n5442, B2 => 
                           n1632, ZN => n9024);
   U1451 : OAI22_X1 port map( A1 => n1726, A2 => n1844, B1 => n5432, B2 => 
                           n1632, ZN => n9023);
   U1452 : OAI22_X1 port map( A1 => n1727, A2 => n1844, B1 => n5422, B2 => 
                           n1632, ZN => n9022);
   U1453 : OAI22_X1 port map( A1 => n1728, A2 => n1844, B1 => n5412, B2 => 
                           n1632, ZN => n9021);
   U1454 : OAI22_X1 port map( A1 => n1729, A2 => n1844, B1 => n5402, B2 => 
                           n1632, ZN => n9020);
   U1455 : OAI22_X1 port map( A1 => n1725, A2 => n1844, B1 => n5392, B2 => 
                           n1632, ZN => n9019);
   U1456 : OAI22_X1 port map( A1 => n1768, A2 => n1844, B1 => n5382, B2 => 
                           n1632, ZN => n9018);
   U1457 : OAI21_X1 port map( B1 => n1769, B2 => n1844, A => n1770, ZN => n1845
                           );
   U1458 : OAI22_X1 port map( A1 => n1759, A2 => n1846, B1 => n5693, B2 => 
                           n1626, ZN => n9017);
   U1459 : OAI22_X1 port map( A1 => n1761, A2 => n1846, B1 => n5683, B2 => 
                           n1626, ZN => n9016);
   U1460 : OAI22_X1 port map( A1 => n1762, A2 => n1846, B1 => n5673, B2 => 
                           n1626, ZN => n9015);
   U1461 : OAI22_X1 port map( A1 => n1763, A2 => n1846, B1 => n5663, B2 => 
                           n1626, ZN => n9014);
   U1462 : OAI22_X1 port map( A1 => n1764, A2 => n1846, B1 => n5653, B2 => 
                           n1626, ZN => n9013);
   U1463 : OAI22_X1 port map( A1 => n1765, A2 => n1846, B1 => n5643, B2 => 
                           n1626, ZN => n9012);
   U1464 : OAI22_X1 port map( A1 => n1766, A2 => n1846, B1 => n5633, B2 => 
                           n1626, ZN => n9011);
   U1465 : OAI22_X1 port map( A1 => n1767, A2 => n1846, B1 => n5623, B2 => 
                           n1626, ZN => n9010);
   U1466 : OAI22_X1 port map( A1 => n1746, A2 => n1846, B1 => n5613, B2 => 
                           n1626, ZN => n9009);
   U1467 : OAI22_X1 port map( A1 => n1747, A2 => n1846, B1 => n5603, B2 => 
                           n1626, ZN => n9008);
   U1468 : OAI22_X1 port map( A1 => n1742, A2 => n1846, B1 => n5593, B2 => 
                           n1626, ZN => n9007);
   U1469 : OAI22_X1 port map( A1 => n1743, A2 => n1846, B1 => n5583, B2 => 
                           n1626, ZN => n9006);
   U1470 : OAI22_X1 port map( A1 => n1744, A2 => n1846, B1 => n5573, B2 => 
                           n1626, ZN => n9005);
   U1471 : OAI22_X1 port map( A1 => n1745, A2 => n1846, B1 => n5563, B2 => 
                           n1626, ZN => n9004);
   U1472 : OAI22_X1 port map( A1 => n1738, A2 => n1846, B1 => n5553, B2 => 
                           n1626, ZN => n9003);
   U1473 : OAI22_X1 port map( A1 => n1739, A2 => n1846, B1 => n5543, B2 => 
                           n1626, ZN => n9002);
   U1474 : OAI22_X1 port map( A1 => n1740, A2 => n1846, B1 => n5533, B2 => 
                           n1626, ZN => n9001);
   U1475 : OAI22_X1 port map( A1 => n1741, A2 => n1846, B1 => n5523, B2 => 
                           n1626, ZN => n9000);
   U1476 : OAI22_X1 port map( A1 => n1734, A2 => n1846, B1 => n5513, B2 => 
                           n1626, ZN => n8999);
   U1477 : OAI22_X1 port map( A1 => n1735, A2 => n1846, B1 => n5503, B2 => 
                           n1626, ZN => n8998);
   U1478 : OAI22_X1 port map( A1 => n1736, A2 => n1846, B1 => n5493, B2 => 
                           n1626, ZN => n8997);
   U1479 : OAI22_X1 port map( A1 => n1737, A2 => n1846, B1 => n5483, B2 => 
                           n1626, ZN => n8996);
   U1480 : OAI22_X1 port map( A1 => n1730, A2 => n1846, B1 => n5473, B2 => 
                           n1626, ZN => n8995);
   U1481 : OAI22_X1 port map( A1 => n1731, A2 => n1846, B1 => n5463, B2 => 
                           n1626, ZN => n8994);
   U1482 : OAI22_X1 port map( A1 => n1732, A2 => n1846, B1 => n5453, B2 => 
                           n1626, ZN => n8993);
   U1483 : OAI22_X1 port map( A1 => n1733, A2 => n1846, B1 => n5443, B2 => 
                           n1626, ZN => n8992);
   U1484 : OAI22_X1 port map( A1 => n1726, A2 => n1846, B1 => n5433, B2 => 
                           n1626, ZN => n8991);
   U1485 : OAI22_X1 port map( A1 => n1727, A2 => n1846, B1 => n5423, B2 => 
                           n1626, ZN => n8990);
   U1486 : OAI22_X1 port map( A1 => n1728, A2 => n1846, B1 => n5413, B2 => 
                           n1626, ZN => n8989);
   U1487 : OAI22_X1 port map( A1 => n1729, A2 => n1846, B1 => n5403, B2 => 
                           n1626, ZN => n8988);
   U1488 : OAI22_X1 port map( A1 => n1725, A2 => n1846, B1 => n5393, B2 => 
                           n1626, ZN => n8987);
   U1489 : OAI22_X1 port map( A1 => n1768, A2 => n1846, B1 => n5383, B2 => 
                           n1626, ZN => n8986);
   U1490 : OAI21_X1 port map( B1 => n1769, B2 => n1846, A => n1770, ZN => n1847
                           );
   U1491 : OAI22_X1 port map( A1 => n1759, A2 => n1848, B1 => n1694, B2 => n905
                           , ZN => n8985);
   U1492 : OAI22_X1 port map( A1 => n1761, A2 => n1848, B1 => n1694, B2 => n906
                           , ZN => n8984);
   U1493 : OAI22_X1 port map( A1 => n1762, A2 => n1848, B1 => n1694, B2 => n907
                           , ZN => n8983);
   U1494 : OAI22_X1 port map( A1 => n1763, A2 => n1848, B1 => n1694, B2 => n908
                           , ZN => n8982);
   U1495 : OAI22_X1 port map( A1 => n1764, A2 => n1848, B1 => n1694, B2 => n909
                           , ZN => n8981);
   U1496 : OAI22_X1 port map( A1 => n1765, A2 => n1848, B1 => n1694, B2 => n910
                           , ZN => n8980);
   U1497 : OAI22_X1 port map( A1 => n1766, A2 => n1848, B1 => n1694, B2 => n911
                           , ZN => n8979);
   U1498 : OAI22_X1 port map( A1 => n1767, A2 => n1848, B1 => n1694, B2 => n912
                           , ZN => n8978);
   U1499 : OAI22_X1 port map( A1 => n1746, A2 => n1848, B1 => n1694, B2 => n913
                           , ZN => n8977);
   U1500 : OAI22_X1 port map( A1 => n1747, A2 => n1848, B1 => n1694, B2 => n914
                           , ZN => n8976);
   U1501 : OAI22_X1 port map( A1 => n1742, A2 => n1848, B1 => n1694, B2 => n915
                           , ZN => n8975);
   U1502 : OAI22_X1 port map( A1 => n1743, A2 => n1848, B1 => n1694, B2 => n916
                           , ZN => n8974);
   U1503 : OAI22_X1 port map( A1 => n1744, A2 => n1848, B1 => n1694, B2 => n917
                           , ZN => n8973);
   U1504 : OAI22_X1 port map( A1 => n1745, A2 => n1848, B1 => n1694, B2 => n918
                           , ZN => n8972);
   U1505 : OAI22_X1 port map( A1 => n1738, A2 => n1848, B1 => n1694, B2 => n919
                           , ZN => n8971);
   U1506 : OAI22_X1 port map( A1 => n1739, A2 => n1848, B1 => n1694, B2 => n920
                           , ZN => n8970);
   U1507 : OAI22_X1 port map( A1 => n1740, A2 => n1848, B1 => n1694, B2 => n921
                           , ZN => n8969);
   U1508 : OAI22_X1 port map( A1 => n1741, A2 => n1848, B1 => n1694, B2 => n922
                           , ZN => n8968);
   U1509 : OAI22_X1 port map( A1 => n1734, A2 => n1848, B1 => n1694, B2 => n923
                           , ZN => n8967);
   U1510 : OAI22_X1 port map( A1 => n1735, A2 => n1848, B1 => n1694, B2 => n924
                           , ZN => n8966);
   U1511 : OAI22_X1 port map( A1 => n1736, A2 => n1848, B1 => n1694, B2 => n925
                           , ZN => n8965);
   U1512 : OAI22_X1 port map( A1 => n1737, A2 => n1848, B1 => n1694, B2 => n926
                           , ZN => n8964);
   U1513 : OAI22_X1 port map( A1 => n1730, A2 => n1848, B1 => n1694, B2 => n927
                           , ZN => n8963);
   U1514 : OAI22_X1 port map( A1 => n1731, A2 => n1848, B1 => n1694, B2 => n928
                           , ZN => n8962);
   U1515 : OAI22_X1 port map( A1 => n1732, A2 => n1848, B1 => n1694, B2 => n929
                           , ZN => n8961);
   U1516 : OAI22_X1 port map( A1 => n1733, A2 => n1848, B1 => n1694, B2 => n930
                           , ZN => n8960);
   U1517 : OAI22_X1 port map( A1 => n1726, A2 => n1848, B1 => n1694, B2 => n931
                           , ZN => n8959);
   U1518 : OAI22_X1 port map( A1 => n1727, A2 => n1848, B1 => n1694, B2 => n932
                           , ZN => n8958);
   U1519 : OAI22_X1 port map( A1 => n1728, A2 => n1848, B1 => n1694, B2 => n933
                           , ZN => n8957);
   U1520 : OAI22_X1 port map( A1 => n1729, A2 => n1848, B1 => n1694, B2 => n934
                           , ZN => n8956);
   U1521 : OAI22_X1 port map( A1 => n1725, A2 => n1848, B1 => n1694, B2 => n935
                           , ZN => n8955);
   U1522 : OAI22_X1 port map( A1 => n1768, A2 => n1848, B1 => n1694, B2 => n936
                           , ZN => n8954);
   U1523 : OAI21_X1 port map( B1 => n1769, B2 => n1848, A => n1770, ZN => n1849
                           );
   U1524 : OAI22_X1 port map( A1 => n1759, A2 => n1851, B1 => n1696, B2 => 
                           n1257, ZN => n8953);
   U1525 : OAI22_X1 port map( A1 => n1761, A2 => n1851, B1 => n1696, B2 => 
                           n1258, ZN => n8952);
   U1526 : OAI22_X1 port map( A1 => n1762, A2 => n1851, B1 => n1696, B2 => 
                           n1259, ZN => n8951);
   U1527 : OAI22_X1 port map( A1 => n1763, A2 => n1851, B1 => n1696, B2 => 
                           n1260, ZN => n8950);
   U1528 : OAI22_X1 port map( A1 => n1764, A2 => n1851, B1 => n1696, B2 => 
                           n1261, ZN => n8949);
   U1529 : OAI22_X1 port map( A1 => n1765, A2 => n1851, B1 => n1696, B2 => 
                           n1262, ZN => n8948);
   U1530 : OAI22_X1 port map( A1 => n1766, A2 => n1851, B1 => n1696, B2 => 
                           n1263, ZN => n8947);
   U1531 : OAI22_X1 port map( A1 => n1767, A2 => n1851, B1 => n1696, B2 => 
                           n1264, ZN => n8946);
   U1532 : OAI22_X1 port map( A1 => n1746, A2 => n1851, B1 => n1696, B2 => 
                           n1265, ZN => n8945);
   U1533 : OAI22_X1 port map( A1 => n1747, A2 => n1851, B1 => n1696, B2 => 
                           n1266, ZN => n8944);
   U1534 : OAI22_X1 port map( A1 => n1742, A2 => n1851, B1 => n1696, B2 => 
                           n1267, ZN => n8943);
   U1535 : OAI22_X1 port map( A1 => n1743, A2 => n1851, B1 => n1696, B2 => 
                           n1268, ZN => n8942);
   U1536 : OAI22_X1 port map( A1 => n1744, A2 => n1851, B1 => n1696, B2 => 
                           n1269, ZN => n8941);
   U1537 : OAI22_X1 port map( A1 => n1745, A2 => n1851, B1 => n1696, B2 => 
                           n1270, ZN => n8940);
   U1538 : OAI22_X1 port map( A1 => n1738, A2 => n1851, B1 => n1696, B2 => 
                           n1271, ZN => n8939);
   U1539 : OAI22_X1 port map( A1 => n1739, A2 => n1851, B1 => n1696, B2 => 
                           n1272, ZN => n8938);
   U1540 : OAI22_X1 port map( A1 => n1740, A2 => n1851, B1 => n1696, B2 => 
                           n1273, ZN => n8937);
   U1541 : OAI22_X1 port map( A1 => n1741, A2 => n1851, B1 => n1696, B2 => 
                           n1274, ZN => n8936);
   U1542 : OAI22_X1 port map( A1 => n1734, A2 => n1851, B1 => n1696, B2 => 
                           n1275, ZN => n8935);
   U1543 : OAI22_X1 port map( A1 => n1735, A2 => n1851, B1 => n1696, B2 => 
                           n1276, ZN => n8934);
   U1544 : OAI22_X1 port map( A1 => n1736, A2 => n1851, B1 => n1696, B2 => 
                           n1277, ZN => n8933);
   U1545 : OAI22_X1 port map( A1 => n1737, A2 => n1851, B1 => n1696, B2 => 
                           n1278, ZN => n8932);
   U1546 : OAI22_X1 port map( A1 => n1730, A2 => n1851, B1 => n1696, B2 => 
                           n1279, ZN => n8931);
   U1547 : OAI22_X1 port map( A1 => n1731, A2 => n1851, B1 => n1696, B2 => 
                           n1280, ZN => n8930);
   U1548 : OAI22_X1 port map( A1 => n1732, A2 => n1851, B1 => n1696, B2 => 
                           n1281, ZN => n8929);
   U1549 : OAI22_X1 port map( A1 => n1733, A2 => n1851, B1 => n1696, B2 => 
                           n1282, ZN => n8928);
   U1550 : OAI22_X1 port map( A1 => n1726, A2 => n1851, B1 => n1696, B2 => 
                           n1283, ZN => n8927);
   U1551 : OAI22_X1 port map( A1 => n1727, A2 => n1851, B1 => n1696, B2 => 
                           n1284, ZN => n8926);
   U1552 : OAI22_X1 port map( A1 => n1728, A2 => n1851, B1 => n1696, B2 => 
                           n1285, ZN => n8925);
   U1553 : OAI22_X1 port map( A1 => n1729, A2 => n1851, B1 => n1696, B2 => 
                           n1286, ZN => n8924);
   U1554 : OAI22_X1 port map( A1 => n1725, A2 => n1851, B1 => n1696, B2 => 
                           n1287, ZN => n8923);
   U1555 : OAI22_X1 port map( A1 => n1768, A2 => n1851, B1 => n1696, B2 => 
                           n1288, ZN => n8922);
   U1556 : OAI21_X1 port map( B1 => n1769, B2 => n1851, A => n1770, ZN => n1852
                           );
   U1557 : OAI22_X1 port map( A1 => n1759, A2 => n1854, B1 => n5089, B2 => 
                           n1628, ZN => n8921);
   U1558 : OAI22_X1 port map( A1 => n1761, A2 => n1854, B1 => n5088, B2 => 
                           n1628, ZN => n8920);
   U1559 : OAI22_X1 port map( A1 => n1762, A2 => n1854, B1 => n5087, B2 => 
                           n1628, ZN => n8919);
   U1560 : OAI22_X1 port map( A1 => n1763, A2 => n1854, B1 => n5086, B2 => 
                           n1628, ZN => n8918);
   U1561 : OAI22_X1 port map( A1 => n1764, A2 => n1854, B1 => n5085, B2 => 
                           n1628, ZN => n8917);
   U1562 : OAI22_X1 port map( A1 => n1765, A2 => n1854, B1 => n5084, B2 => 
                           n1628, ZN => n8916);
   U1563 : OAI22_X1 port map( A1 => n1766, A2 => n1854, B1 => n5083, B2 => 
                           n1628, ZN => n8915);
   U1564 : OAI22_X1 port map( A1 => n1767, A2 => n1854, B1 => n5082, B2 => 
                           n1628, ZN => n8914);
   U1565 : OAI22_X1 port map( A1 => n1746, A2 => n1854, B1 => n5081, B2 => 
                           n1628, ZN => n8913);
   U1566 : OAI22_X1 port map( A1 => n1747, A2 => n1854, B1 => n5080, B2 => 
                           n1628, ZN => n8912);
   U1567 : OAI22_X1 port map( A1 => n1742, A2 => n1854, B1 => n5079, B2 => 
                           n1628, ZN => n8911);
   U1568 : OAI22_X1 port map( A1 => n1743, A2 => n1854, B1 => n5078, B2 => 
                           n1628, ZN => n8910);
   U1569 : OAI22_X1 port map( A1 => n1744, A2 => n1854, B1 => n5077, B2 => 
                           n1628, ZN => n8909);
   U1570 : OAI22_X1 port map( A1 => n1745, A2 => n1854, B1 => n5076, B2 => 
                           n1628, ZN => n8908);
   U1571 : OAI22_X1 port map( A1 => n1738, A2 => n1854, B1 => n5075, B2 => 
                           n1628, ZN => n8907);
   U1572 : OAI22_X1 port map( A1 => n1739, A2 => n1854, B1 => n5074, B2 => 
                           n1628, ZN => n8906);
   U1573 : OAI22_X1 port map( A1 => n1740, A2 => n1854, B1 => n5073, B2 => 
                           n1628, ZN => n8905);
   U1574 : OAI22_X1 port map( A1 => n1741, A2 => n1854, B1 => n5072, B2 => 
                           n1628, ZN => n8904);
   U1575 : OAI22_X1 port map( A1 => n1734, A2 => n1854, B1 => n5071, B2 => 
                           n1628, ZN => n8903);
   U1576 : OAI22_X1 port map( A1 => n1735, A2 => n1854, B1 => n5070, B2 => 
                           n1628, ZN => n8902);
   U1577 : OAI22_X1 port map( A1 => n1736, A2 => n1854, B1 => n5069, B2 => 
                           n1628, ZN => n8901);
   U1578 : OAI22_X1 port map( A1 => n1737, A2 => n1854, B1 => n5068, B2 => 
                           n1628, ZN => n8900);
   U1579 : OAI22_X1 port map( A1 => n1730, A2 => n1854, B1 => n5067, B2 => 
                           n1628, ZN => n8899);
   U1580 : OAI22_X1 port map( A1 => n1731, A2 => n1854, B1 => n5066, B2 => 
                           n1628, ZN => n8898);
   U1581 : OAI22_X1 port map( A1 => n1732, A2 => n1854, B1 => n5065, B2 => 
                           n1628, ZN => n8897);
   U1582 : OAI22_X1 port map( A1 => n1733, A2 => n1854, B1 => n5064, B2 => 
                           n1628, ZN => n8896);
   U1583 : OAI22_X1 port map( A1 => n1726, A2 => n1854, B1 => n5063, B2 => 
                           n1628, ZN => n8895);
   U1584 : OAI22_X1 port map( A1 => n1727, A2 => n1854, B1 => n5062, B2 => 
                           n1628, ZN => n8894);
   U1585 : OAI22_X1 port map( A1 => n1728, A2 => n1854, B1 => n5061, B2 => 
                           n1628, ZN => n8893);
   U1586 : OAI22_X1 port map( A1 => n1729, A2 => n1854, B1 => n5060, B2 => 
                           n1628, ZN => n8892);
   U1587 : OAI22_X1 port map( A1 => n1725, A2 => n1854, B1 => n5059, B2 => 
                           n1628, ZN => n8891);
   U1588 : OAI22_X1 port map( A1 => n1768, A2 => n1854, B1 => n5058, B2 => 
                           n1628, ZN => n8890);
   U1589 : OAI21_X1 port map( B1 => n1769, B2 => n1854, A => n1770, ZN => n1855
                           );
   U1590 : OAI22_X1 port map( A1 => n1759, A2 => n1856, B1 => n5057, B2 => 
                           n1622, ZN => n8889);
   U1591 : OAI22_X1 port map( A1 => n1761, A2 => n1856, B1 => n5056, B2 => 
                           n1622, ZN => n8888);
   U1592 : OAI22_X1 port map( A1 => n1762, A2 => n1856, B1 => n5055, B2 => 
                           n1622, ZN => n8887);
   U1593 : OAI22_X1 port map( A1 => n1763, A2 => n1856, B1 => n5054, B2 => 
                           n1622, ZN => n8886);
   U1594 : OAI22_X1 port map( A1 => n1764, A2 => n1856, B1 => n5053, B2 => 
                           n1622, ZN => n8885);
   U1595 : OAI22_X1 port map( A1 => n1765, A2 => n1856, B1 => n5052, B2 => 
                           n1622, ZN => n8884);
   U1596 : OAI22_X1 port map( A1 => n1766, A2 => n1856, B1 => n5051, B2 => 
                           n1622, ZN => n8883);
   U1597 : OAI22_X1 port map( A1 => n1767, A2 => n1856, B1 => n5050, B2 => 
                           n1622, ZN => n8882);
   U1598 : OAI22_X1 port map( A1 => n1746, A2 => n1856, B1 => n5049, B2 => 
                           n1622, ZN => n8881);
   U1599 : OAI22_X1 port map( A1 => n1747, A2 => n1856, B1 => n5048, B2 => 
                           n1622, ZN => n8880);
   U1600 : OAI22_X1 port map( A1 => n1742, A2 => n1856, B1 => n5047, B2 => 
                           n1622, ZN => n8879);
   U1601 : OAI22_X1 port map( A1 => n1743, A2 => n1856, B1 => n5046, B2 => 
                           n1622, ZN => n8878);
   U1602 : OAI22_X1 port map( A1 => n1744, A2 => n1856, B1 => n5045, B2 => 
                           n1622, ZN => n8877);
   U1603 : OAI22_X1 port map( A1 => n1745, A2 => n1856, B1 => n5044, B2 => 
                           n1622, ZN => n8876);
   U1604 : OAI22_X1 port map( A1 => n1738, A2 => n1856, B1 => n5043, B2 => 
                           n1622, ZN => n8875);
   U1605 : OAI22_X1 port map( A1 => n1739, A2 => n1856, B1 => n5042, B2 => 
                           n1622, ZN => n8874);
   U1606 : OAI22_X1 port map( A1 => n1740, A2 => n1856, B1 => n5041, B2 => 
                           n1622, ZN => n8873);
   U1607 : OAI22_X1 port map( A1 => n1741, A2 => n1856, B1 => n5040, B2 => 
                           n1622, ZN => n8872);
   U1608 : OAI22_X1 port map( A1 => n1734, A2 => n1856, B1 => n5039, B2 => 
                           n1622, ZN => n8871);
   U1609 : OAI22_X1 port map( A1 => n1735, A2 => n1856, B1 => n5038, B2 => 
                           n1622, ZN => n8870);
   U1610 : OAI22_X1 port map( A1 => n1736, A2 => n1856, B1 => n5037, B2 => 
                           n1622, ZN => n8869);
   U1611 : OAI22_X1 port map( A1 => n1737, A2 => n1856, B1 => n5036, B2 => 
                           n1622, ZN => n8868);
   U1612 : OAI22_X1 port map( A1 => n1730, A2 => n1856, B1 => n5035, B2 => 
                           n1622, ZN => n8867);
   U1613 : OAI22_X1 port map( A1 => n1731, A2 => n1856, B1 => n5034, B2 => 
                           n1622, ZN => n8866);
   U1614 : OAI22_X1 port map( A1 => n1732, A2 => n1856, B1 => n5033, B2 => 
                           n1622, ZN => n8865);
   U1615 : OAI22_X1 port map( A1 => n1733, A2 => n1856, B1 => n5032, B2 => 
                           n1622, ZN => n8864);
   U1616 : OAI22_X1 port map( A1 => n1726, A2 => n1856, B1 => n5031, B2 => 
                           n1622, ZN => n8863);
   U1617 : OAI22_X1 port map( A1 => n1727, A2 => n1856, B1 => n5030, B2 => 
                           n1622, ZN => n8862);
   U1618 : OAI22_X1 port map( A1 => n1728, A2 => n1856, B1 => n5029, B2 => 
                           n1622, ZN => n8861);
   U1619 : OAI22_X1 port map( A1 => n1729, A2 => n1856, B1 => n5028, B2 => 
                           n1622, ZN => n8860);
   U1620 : OAI22_X1 port map( A1 => n1725, A2 => n1856, B1 => n5027, B2 => 
                           n1622, ZN => n8859);
   U1621 : OAI22_X1 port map( A1 => n1768, A2 => n1856, B1 => n5026, B2 => 
                           n1622, ZN => n8858);
   U1622 : OAI21_X1 port map( B1 => n1769, B2 => n1856, A => n1770, ZN => n1857
                           );
   U1623 : OAI22_X1 port map( A1 => n1759, A2 => n1858, B1 => n5025, B2 => 
                           n1624, ZN => n8857);
   U1624 : OAI22_X1 port map( A1 => n1761, A2 => n1858, B1 => n5024, B2 => 
                           n1624, ZN => n8856);
   U1625 : OAI22_X1 port map( A1 => n1762, A2 => n1858, B1 => n5023, B2 => 
                           n1624, ZN => n8855);
   U1626 : OAI22_X1 port map( A1 => n1763, A2 => n1858, B1 => n5022, B2 => 
                           n1624, ZN => n8854);
   U1627 : OAI22_X1 port map( A1 => n1764, A2 => n1858, B1 => n5021, B2 => 
                           n1624, ZN => n8853);
   U1628 : OAI22_X1 port map( A1 => n1765, A2 => n1858, B1 => n5020, B2 => 
                           n1624, ZN => n8852);
   U1629 : OAI22_X1 port map( A1 => n1766, A2 => n1858, B1 => n5019, B2 => 
                           n1624, ZN => n8851);
   U1630 : OAI22_X1 port map( A1 => n1767, A2 => n1858, B1 => n5018, B2 => 
                           n1624, ZN => n8850);
   U1631 : OAI22_X1 port map( A1 => n1746, A2 => n1858, B1 => n5017, B2 => 
                           n1624, ZN => n8849);
   U1632 : OAI22_X1 port map( A1 => n1747, A2 => n1858, B1 => n5016, B2 => 
                           n1624, ZN => n8848);
   U1633 : OAI22_X1 port map( A1 => n1742, A2 => n1858, B1 => n5015, B2 => 
                           n1624, ZN => n8847);
   U1634 : OAI22_X1 port map( A1 => n1743, A2 => n1858, B1 => n5014, B2 => 
                           n1624, ZN => n8846);
   U1635 : OAI22_X1 port map( A1 => n1744, A2 => n1858, B1 => n5013, B2 => 
                           n1624, ZN => n8845);
   U1636 : OAI22_X1 port map( A1 => n1745, A2 => n1858, B1 => n5012, B2 => 
                           n1624, ZN => n8844);
   U1637 : OAI22_X1 port map( A1 => n1738, A2 => n1858, B1 => n5011, B2 => 
                           n1624, ZN => n8843);
   U1638 : OAI22_X1 port map( A1 => n1739, A2 => n1858, B1 => n5010, B2 => 
                           n1624, ZN => n8842);
   U1639 : OAI22_X1 port map( A1 => n1740, A2 => n1858, B1 => n5009, B2 => 
                           n1624, ZN => n8841);
   U1640 : OAI22_X1 port map( A1 => n1741, A2 => n1858, B1 => n5008, B2 => 
                           n1624, ZN => n8840);
   U1641 : OAI22_X1 port map( A1 => n1734, A2 => n1858, B1 => n5007, B2 => 
                           n1624, ZN => n8839);
   U1642 : OAI22_X1 port map( A1 => n1735, A2 => n1858, B1 => n5006, B2 => 
                           n1624, ZN => n8838);
   U1643 : OAI22_X1 port map( A1 => n1736, A2 => n1858, B1 => n5005, B2 => 
                           n1624, ZN => n8837);
   U1644 : OAI22_X1 port map( A1 => n1737, A2 => n1858, B1 => n5004, B2 => 
                           n1624, ZN => n8836);
   U1645 : OAI22_X1 port map( A1 => n1730, A2 => n1858, B1 => n5003, B2 => 
                           n1624, ZN => n8835);
   U1646 : OAI22_X1 port map( A1 => n1731, A2 => n1858, B1 => n5002, B2 => 
                           n1624, ZN => n8834);
   U1647 : OAI22_X1 port map( A1 => n1732, A2 => n1858, B1 => n5001, B2 => 
                           n1624, ZN => n8833);
   U1648 : OAI22_X1 port map( A1 => n1733, A2 => n1858, B1 => n5000, B2 => 
                           n1624, ZN => n8832);
   U1649 : OAI22_X1 port map( A1 => n1726, A2 => n1858, B1 => n4999, B2 => 
                           n1624, ZN => n8831);
   U1650 : OAI22_X1 port map( A1 => n1727, A2 => n1858, B1 => n4998, B2 => 
                           n1624, ZN => n8830);
   U1651 : OAI22_X1 port map( A1 => n1728, A2 => n1858, B1 => n4997, B2 => 
                           n1624, ZN => n8829);
   U1652 : OAI22_X1 port map( A1 => n1729, A2 => n1858, B1 => n4996, B2 => 
                           n1624, ZN => n8828);
   U1653 : OAI22_X1 port map( A1 => n1725, A2 => n1858, B1 => n4995, B2 => 
                           n1624, ZN => n8827);
   U1654 : OAI22_X1 port map( A1 => n1768, A2 => n1858, B1 => n4994, B2 => 
                           n1624, ZN => n8826);
   U1655 : OAI21_X1 port map( B1 => n1769, B2 => n1858, A => n1770, ZN => n1859
                           );
   U1656 : OAI22_X1 port map( A1 => n1759, A2 => n1860, B1 => n1690, B2 => n458
                           , ZN => n8825);
   U1657 : OAI22_X1 port map( A1 => n1761, A2 => n1860, B1 => n1690, B2 => n460
                           , ZN => n8824);
   U1658 : OAI22_X1 port map( A1 => n1762, A2 => n1860, B1 => n1690, B2 => n462
                           , ZN => n8823);
   U1659 : OAI22_X1 port map( A1 => n1763, A2 => n1860, B1 => n1690, B2 => n464
                           , ZN => n8822);
   U1660 : OAI22_X1 port map( A1 => n1764, A2 => n1860, B1 => n1690, B2 => n466
                           , ZN => n8821);
   U1661 : OAI22_X1 port map( A1 => n1765, A2 => n1860, B1 => n1690, B2 => n468
                           , ZN => n8820);
   U1662 : OAI22_X1 port map( A1 => n1766, A2 => n1860, B1 => n1690, B2 => n470
                           , ZN => n8819);
   U1663 : OAI22_X1 port map( A1 => n1767, A2 => n1860, B1 => n1690, B2 => n472
                           , ZN => n8818);
   U1664 : OAI22_X1 port map( A1 => n1746, A2 => n1860, B1 => n1690, B2 => n474
                           , ZN => n8817);
   U1665 : OAI22_X1 port map( A1 => n1747, A2 => n1860, B1 => n1690, B2 => n476
                           , ZN => n8816);
   U1666 : OAI22_X1 port map( A1 => n1742, A2 => n1860, B1 => n1690, B2 => n478
                           , ZN => n8815);
   U1667 : OAI22_X1 port map( A1 => n1743, A2 => n1860, B1 => n1690, B2 => n480
                           , ZN => n8814);
   U1668 : OAI22_X1 port map( A1 => n1744, A2 => n1860, B1 => n1690, B2 => n482
                           , ZN => n8813);
   U1669 : OAI22_X1 port map( A1 => n1745, A2 => n1860, B1 => n1690, B2 => n484
                           , ZN => n8812);
   U1670 : OAI22_X1 port map( A1 => n1738, A2 => n1860, B1 => n1690, B2 => n486
                           , ZN => n8811);
   U1671 : OAI22_X1 port map( A1 => n1739, A2 => n1860, B1 => n1690, B2 => n488
                           , ZN => n8810);
   U1672 : OAI22_X1 port map( A1 => n1740, A2 => n1860, B1 => n1690, B2 => n490
                           , ZN => n8809);
   U1673 : OAI22_X1 port map( A1 => n1741, A2 => n1860, B1 => n1690, B2 => n492
                           , ZN => n8808);
   U1674 : OAI22_X1 port map( A1 => n1734, A2 => n1860, B1 => n1690, B2 => n494
                           , ZN => n8807);
   U1675 : OAI22_X1 port map( A1 => n1735, A2 => n1860, B1 => n1690, B2 => n496
                           , ZN => n8806);
   U1676 : OAI22_X1 port map( A1 => n1736, A2 => n1860, B1 => n1690, B2 => n498
                           , ZN => n8805);
   U1677 : OAI22_X1 port map( A1 => n1737, A2 => n1860, B1 => n1690, B2 => n500
                           , ZN => n8804);
   U1678 : OAI22_X1 port map( A1 => n1730, A2 => n1860, B1 => n1690, B2 => n502
                           , ZN => n8803);
   U1679 : OAI22_X1 port map( A1 => n1731, A2 => n1860, B1 => n1690, B2 => n504
                           , ZN => n8802);
   U1680 : OAI22_X1 port map( A1 => n1732, A2 => n1860, B1 => n1690, B2 => n506
                           , ZN => n8801);
   U1681 : OAI22_X1 port map( A1 => n1733, A2 => n1860, B1 => n1690, B2 => n508
                           , ZN => n8800);
   U1682 : OAI22_X1 port map( A1 => n1726, A2 => n1860, B1 => n1690, B2 => n510
                           , ZN => n8799);
   U1683 : OAI22_X1 port map( A1 => n1727, A2 => n1860, B1 => n1690, B2 => n512
                           , ZN => n8798);
   U1684 : OAI22_X1 port map( A1 => n1728, A2 => n1860, B1 => n1690, B2 => n514
                           , ZN => n8797);
   U1685 : OAI22_X1 port map( A1 => n1729, A2 => n1860, B1 => n1690, B2 => n516
                           , ZN => n8796);
   U1686 : OAI22_X1 port map( A1 => n1725, A2 => n1860, B1 => n1690, B2 => n518
                           , ZN => n8795);
   U1687 : OAI22_X1 port map( A1 => n1768, A2 => n1860, B1 => n1690, B2 => n520
                           , ZN => n8794);
   U1688 : OAI21_X1 port map( B1 => n1769, B2 => n1860, A => n1770, ZN => n1861
                           );
   U1689 : OAI22_X1 port map( A1 => n1759, A2 => n1862, B1 => n1692, B2 => n2, 
                           ZN => n8793);
   U1690 : OAI22_X1 port map( A1 => n1761, A2 => n1862, B1 => n1692, B2 => n4, 
                           ZN => n8792);
   U1691 : OAI22_X1 port map( A1 => n1762, A2 => n1862, B1 => n1692, B2 => n6, 
                           ZN => n8791);
   U1692 : OAI22_X1 port map( A1 => n1763, A2 => n1862, B1 => n1692, B2 => n8, 
                           ZN => n8790);
   U1693 : OAI22_X1 port map( A1 => n1764, A2 => n1862, B1 => n1692, B2 => n10,
                           ZN => n8789);
   U1694 : OAI22_X1 port map( A1 => n1765, A2 => n1862, B1 => n1692, B2 => n12,
                           ZN => n8788);
   U1695 : OAI22_X1 port map( A1 => n1766, A2 => n1862, B1 => n1692, B2 => n14,
                           ZN => n8787);
   U1696 : OAI22_X1 port map( A1 => n1767, A2 => n1862, B1 => n1692, B2 => n16,
                           ZN => n8786);
   U1697 : OAI22_X1 port map( A1 => n1746, A2 => n1862, B1 => n1692, B2 => n18,
                           ZN => n8785);
   U1698 : OAI22_X1 port map( A1 => n1747, A2 => n1862, B1 => n1692, B2 => n20,
                           ZN => n8784);
   U1699 : OAI22_X1 port map( A1 => n1742, A2 => n1862, B1 => n1692, B2 => n22,
                           ZN => n8783);
   U1700 : OAI22_X1 port map( A1 => n1743, A2 => n1862, B1 => n1692, B2 => n24,
                           ZN => n8782);
   U1701 : OAI22_X1 port map( A1 => n1744, A2 => n1862, B1 => n1692, B2 => n26,
                           ZN => n8781);
   U1702 : OAI22_X1 port map( A1 => n1745, A2 => n1862, B1 => n1692, B2 => n28,
                           ZN => n8780);
   U1703 : OAI22_X1 port map( A1 => n1738, A2 => n1862, B1 => n1692, B2 => n30,
                           ZN => n8779);
   U1704 : OAI22_X1 port map( A1 => n1739, A2 => n1862, B1 => n1692, B2 => n32,
                           ZN => n8778);
   U1705 : OAI22_X1 port map( A1 => n1740, A2 => n1862, B1 => n1692, B2 => n34,
                           ZN => n8777);
   U1706 : OAI22_X1 port map( A1 => n1741, A2 => n1862, B1 => n1692, B2 => n36,
                           ZN => n8776);
   U1707 : OAI22_X1 port map( A1 => n1734, A2 => n1862, B1 => n1692, B2 => n38,
                           ZN => n8775);
   U1708 : OAI22_X1 port map( A1 => n1735, A2 => n1862, B1 => n1692, B2 => n40,
                           ZN => n8774);
   U1709 : OAI22_X1 port map( A1 => n1736, A2 => n1862, B1 => n1692, B2 => n42,
                           ZN => n8773);
   U1710 : OAI22_X1 port map( A1 => n1737, A2 => n1862, B1 => n1692, B2 => n44,
                           ZN => n8772);
   U1711 : OAI22_X1 port map( A1 => n1730, A2 => n1862, B1 => n1692, B2 => n46,
                           ZN => n8771);
   U1712 : OAI22_X1 port map( A1 => n1731, A2 => n1862, B1 => n1692, B2 => n48,
                           ZN => n8770);
   U1713 : OAI22_X1 port map( A1 => n1732, A2 => n1862, B1 => n1692, B2 => n50,
                           ZN => n8769);
   U1714 : OAI22_X1 port map( A1 => n1733, A2 => n1862, B1 => n1692, B2 => n52,
                           ZN => n8768);
   U1715 : OAI22_X1 port map( A1 => n1726, A2 => n1862, B1 => n1692, B2 => n54,
                           ZN => n8767);
   U1716 : OAI22_X1 port map( A1 => n1727, A2 => n1862, B1 => n1692, B2 => n56,
                           ZN => n8766);
   U1717 : OAI22_X1 port map( A1 => n1728, A2 => n1862, B1 => n1692, B2 => n58,
                           ZN => n8765);
   U1718 : OAI22_X1 port map( A1 => n1729, A2 => n1862, B1 => n1692, B2 => n60,
                           ZN => n8764);
   U1719 : OAI22_X1 port map( A1 => n1725, A2 => n1862, B1 => n1692, B2 => n62,
                           ZN => n8763);
   U1720 : OAI22_X1 port map( A1 => n1768, A2 => n1862, B1 => n1692, B2 => n64,
                           ZN => n8762);
   U1721 : OAI21_X1 port map( B1 => n1769, B2 => n1862, A => n1770, ZN => n1863
                           );
   U1722 : OAI22_X1 port map( A1 => n1759, A2 => n1864, B1 => n5822, B2 => 
                           n1618, ZN => n8761);
   U1723 : OAI22_X1 port map( A1 => n1761, A2 => n1864, B1 => n5818, B2 => 
                           n1618, ZN => n8760);
   U1724 : OAI22_X1 port map( A1 => n1762, A2 => n1864, B1 => n5814, B2 => 
                           n1618, ZN => n8759);
   U1725 : OAI22_X1 port map( A1 => n1763, A2 => n1864, B1 => n5810, B2 => 
                           n1618, ZN => n8758);
   U1726 : OAI22_X1 port map( A1 => n1764, A2 => n1864, B1 => n5806, B2 => 
                           n1618, ZN => n8757);
   U1727 : OAI22_X1 port map( A1 => n1765, A2 => n1864, B1 => n5802, B2 => 
                           n1618, ZN => n8756);
   U1728 : OAI22_X1 port map( A1 => n1766, A2 => n1864, B1 => n5798, B2 => 
                           n1618, ZN => n8755);
   U1729 : OAI22_X1 port map( A1 => n1767, A2 => n1864, B1 => n5794, B2 => 
                           n1618, ZN => n8754);
   U1730 : OAI22_X1 port map( A1 => n1746, A2 => n1864, B1 => n5790, B2 => 
                           n1618, ZN => n8753);
   U1731 : OAI22_X1 port map( A1 => n1747, A2 => n1864, B1 => n5786, B2 => 
                           n1618, ZN => n8752);
   U1732 : OAI22_X1 port map( A1 => n1742, A2 => n1864, B1 => n5782, B2 => 
                           n1618, ZN => n8751);
   U1733 : OAI22_X1 port map( A1 => n1743, A2 => n1864, B1 => n5778, B2 => 
                           n1618, ZN => n8750);
   U1734 : OAI22_X1 port map( A1 => n1744, A2 => n1864, B1 => n5774, B2 => 
                           n1618, ZN => n8749);
   U1735 : OAI22_X1 port map( A1 => n1745, A2 => n1864, B1 => n5770, B2 => 
                           n1618, ZN => n8748);
   U1736 : OAI22_X1 port map( A1 => n1738, A2 => n1864, B1 => n5766, B2 => 
                           n1618, ZN => n8747);
   U1737 : OAI22_X1 port map( A1 => n1739, A2 => n1864, B1 => n5762, B2 => 
                           n1618, ZN => n8746);
   U1738 : OAI22_X1 port map( A1 => n1740, A2 => n1864, B1 => n5758, B2 => 
                           n1618, ZN => n8745);
   U1739 : OAI22_X1 port map( A1 => n1741, A2 => n1864, B1 => n5754, B2 => 
                           n1618, ZN => n8744);
   U1740 : OAI22_X1 port map( A1 => n1734, A2 => n1864, B1 => n5750, B2 => 
                           n1618, ZN => n8743);
   U1741 : OAI22_X1 port map( A1 => n1735, A2 => n1864, B1 => n5746, B2 => 
                           n1618, ZN => n8742);
   U1742 : OAI22_X1 port map( A1 => n1736, A2 => n1864, B1 => n5742, B2 => 
                           n1618, ZN => n8741);
   U1743 : OAI22_X1 port map( A1 => n1737, A2 => n1864, B1 => n5738, B2 => 
                           n1618, ZN => n8740);
   U1744 : OAI22_X1 port map( A1 => n1730, A2 => n1864, B1 => n5734, B2 => 
                           n1618, ZN => n8739);
   U1745 : OAI22_X1 port map( A1 => n1731, A2 => n1864, B1 => n5730, B2 => 
                           n1618, ZN => n8738);
   U1746 : OAI22_X1 port map( A1 => n1732, A2 => n1864, B1 => n5726, B2 => 
                           n1618, ZN => n8737);
   U1747 : OAI22_X1 port map( A1 => n1733, A2 => n1864, B1 => n5722, B2 => 
                           n1618, ZN => n8736);
   U1748 : OAI22_X1 port map( A1 => n1726, A2 => n1864, B1 => n5718, B2 => 
                           n1618, ZN => n8735);
   U1749 : OAI22_X1 port map( A1 => n1727, A2 => n1864, B1 => n5714, B2 => 
                           n1618, ZN => n8734);
   U1750 : OAI22_X1 port map( A1 => n1728, A2 => n1864, B1 => n5710, B2 => 
                           n1618, ZN => n8733);
   U1751 : OAI22_X1 port map( A1 => n1729, A2 => n1864, B1 => n5706, B2 => 
                           n1618, ZN => n8732);
   U1752 : OAI22_X1 port map( A1 => n1725, A2 => n1864, B1 => n5702, B2 => 
                           n1618, ZN => n8731);
   U1753 : OAI22_X1 port map( A1 => n1768, A2 => n1864, B1 => n5698, B2 => 
                           n1618, ZN => n8730);
   U1754 : OAI21_X1 port map( B1 => n1769, B2 => n1864, A => n1770, ZN => n1865
                           );
   U1755 : OAI22_X1 port map( A1 => n1759, A2 => n1866, B1 => n5823, B2 => 
                           n1620, ZN => n8729);
   U1756 : OAI22_X1 port map( A1 => n1761, A2 => n1866, B1 => n5819, B2 => 
                           n1620, ZN => n8728);
   U1757 : OAI22_X1 port map( A1 => n1762, A2 => n1866, B1 => n5815, B2 => 
                           n1620, ZN => n8727);
   U1758 : OAI22_X1 port map( A1 => n1763, A2 => n1866, B1 => n5811, B2 => 
                           n1620, ZN => n8726);
   U1759 : OAI22_X1 port map( A1 => n1764, A2 => n1866, B1 => n5807, B2 => 
                           n1620, ZN => n8725);
   U1760 : OAI22_X1 port map( A1 => n1765, A2 => n1866, B1 => n5803, B2 => 
                           n1620, ZN => n8724);
   U1761 : OAI22_X1 port map( A1 => n1766, A2 => n1866, B1 => n5799, B2 => 
                           n1620, ZN => n8723);
   U1762 : OAI22_X1 port map( A1 => n1767, A2 => n1866, B1 => n5795, B2 => 
                           n1620, ZN => n8722);
   U1763 : OAI22_X1 port map( A1 => n1746, A2 => n1866, B1 => n5791, B2 => 
                           n1620, ZN => n8721);
   U1764 : OAI22_X1 port map( A1 => n1747, A2 => n1866, B1 => n5787, B2 => 
                           n1620, ZN => n8720);
   U1765 : OAI22_X1 port map( A1 => n1742, A2 => n1866, B1 => n5783, B2 => 
                           n1620, ZN => n8719);
   U1766 : OAI22_X1 port map( A1 => n1743, A2 => n1866, B1 => n5779, B2 => 
                           n1620, ZN => n8718);
   U1767 : OAI22_X1 port map( A1 => n1744, A2 => n1866, B1 => n5775, B2 => 
                           n1620, ZN => n8717);
   U1768 : OAI22_X1 port map( A1 => n1745, A2 => n1866, B1 => n5771, B2 => 
                           n1620, ZN => n8716);
   U1769 : OAI22_X1 port map( A1 => n1738, A2 => n1866, B1 => n5767, B2 => 
                           n1620, ZN => n8715);
   U1770 : OAI22_X1 port map( A1 => n1739, A2 => n1866, B1 => n5763, B2 => 
                           n1620, ZN => n8714);
   U1771 : OAI22_X1 port map( A1 => n1740, A2 => n1866, B1 => n5759, B2 => 
                           n1620, ZN => n8713);
   U1772 : OAI22_X1 port map( A1 => n1741, A2 => n1866, B1 => n5755, B2 => 
                           n1620, ZN => n8712);
   U1773 : OAI22_X1 port map( A1 => n1734, A2 => n1866, B1 => n5751, B2 => 
                           n1620, ZN => n8711);
   U1774 : OAI22_X1 port map( A1 => n1735, A2 => n1866, B1 => n5747, B2 => 
                           n1620, ZN => n8710);
   U1775 : OAI22_X1 port map( A1 => n1736, A2 => n1866, B1 => n5743, B2 => 
                           n1620, ZN => n8709);
   U1776 : OAI22_X1 port map( A1 => n1737, A2 => n1866, B1 => n5739, B2 => 
                           n1620, ZN => n8708);
   U1777 : OAI22_X1 port map( A1 => n1730, A2 => n1866, B1 => n5735, B2 => 
                           n1620, ZN => n8707);
   U1778 : OAI22_X1 port map( A1 => n1731, A2 => n1866, B1 => n5731, B2 => 
                           n1620, ZN => n8706);
   U1779 : OAI22_X1 port map( A1 => n1732, A2 => n1866, B1 => n5727, B2 => 
                           n1620, ZN => n8705);
   U1780 : OAI22_X1 port map( A1 => n1733, A2 => n1866, B1 => n5723, B2 => 
                           n1620, ZN => n8704);
   U1781 : OAI22_X1 port map( A1 => n1726, A2 => n1866, B1 => n5719, B2 => 
                           n1620, ZN => n8703);
   U1782 : OAI22_X1 port map( A1 => n1727, A2 => n1866, B1 => n5715, B2 => 
                           n1620, ZN => n8702);
   U1783 : OAI22_X1 port map( A1 => n1728, A2 => n1866, B1 => n5711, B2 => 
                           n1620, ZN => n8701);
   U1784 : OAI22_X1 port map( A1 => n1729, A2 => n1866, B1 => n5707, B2 => 
                           n1620, ZN => n8700);
   U1785 : OAI22_X1 port map( A1 => n1725, A2 => n1866, B1 => n5703, B2 => 
                           n1620, ZN => n8699);
   U1786 : OAI22_X1 port map( A1 => n1768, A2 => n1866, B1 => n5699, B2 => 
                           n1620, ZN => n8698);
   U1787 : OAI21_X1 port map( B1 => n1769, B2 => n1866, A => n1770, ZN => n1867
                           );
   U1788 : OAI22_X1 port map( A1 => n1759, A2 => n1868, B1 => n1686, B2 => n937
                           , ZN => n8697);
   U1789 : OAI22_X1 port map( A1 => n1761, A2 => n1868, B1 => n1686, B2 => n938
                           , ZN => n8696);
   U1790 : OAI22_X1 port map( A1 => n1762, A2 => n1868, B1 => n1686, B2 => n939
                           , ZN => n8695);
   U1791 : OAI22_X1 port map( A1 => n1763, A2 => n1868, B1 => n1686, B2 => n940
                           , ZN => n8694);
   U1792 : OAI22_X1 port map( A1 => n1764, A2 => n1868, B1 => n1686, B2 => n941
                           , ZN => n8693);
   U1793 : OAI22_X1 port map( A1 => n1765, A2 => n1868, B1 => n1686, B2 => n942
                           , ZN => n8692);
   U1794 : OAI22_X1 port map( A1 => n1766, A2 => n1868, B1 => n1686, B2 => n943
                           , ZN => n8691);
   U1795 : OAI22_X1 port map( A1 => n1767, A2 => n1868, B1 => n1686, B2 => n944
                           , ZN => n8690);
   U1796 : OAI22_X1 port map( A1 => n1746, A2 => n1868, B1 => n1686, B2 => n945
                           , ZN => n8689);
   U1797 : OAI22_X1 port map( A1 => n1747, A2 => n1868, B1 => n1686, B2 => n946
                           , ZN => n8688);
   U1798 : OAI22_X1 port map( A1 => n1742, A2 => n1868, B1 => n1686, B2 => n947
                           , ZN => n8687);
   U1799 : OAI22_X1 port map( A1 => n1743, A2 => n1868, B1 => n1686, B2 => n948
                           , ZN => n8686);
   U1800 : OAI22_X1 port map( A1 => n1744, A2 => n1868, B1 => n1686, B2 => n949
                           , ZN => n8685);
   U1801 : OAI22_X1 port map( A1 => n1745, A2 => n1868, B1 => n1686, B2 => n950
                           , ZN => n8684);
   U1802 : OAI22_X1 port map( A1 => n1738, A2 => n1868, B1 => n1686, B2 => n951
                           , ZN => n8683);
   U1803 : OAI22_X1 port map( A1 => n1739, A2 => n1868, B1 => n1686, B2 => n952
                           , ZN => n8682);
   U1804 : OAI22_X1 port map( A1 => n1740, A2 => n1868, B1 => n1686, B2 => n953
                           , ZN => n8681);
   U1805 : OAI22_X1 port map( A1 => n1741, A2 => n1868, B1 => n1686, B2 => n954
                           , ZN => n8680);
   U1806 : OAI22_X1 port map( A1 => n1734, A2 => n1868, B1 => n1686, B2 => n955
                           , ZN => n8679);
   U1807 : OAI22_X1 port map( A1 => n1735, A2 => n1868, B1 => n1686, B2 => n956
                           , ZN => n8678);
   U1808 : OAI22_X1 port map( A1 => n1736, A2 => n1868, B1 => n1686, B2 => n957
                           , ZN => n8677);
   U1809 : OAI22_X1 port map( A1 => n1737, A2 => n1868, B1 => n1686, B2 => n958
                           , ZN => n8676);
   U1810 : OAI22_X1 port map( A1 => n1730, A2 => n1868, B1 => n1686, B2 => n959
                           , ZN => n8675);
   U1811 : OAI22_X1 port map( A1 => n1731, A2 => n1868, B1 => n1686, B2 => n960
                           , ZN => n8674);
   U1812 : OAI22_X1 port map( A1 => n1732, A2 => n1868, B1 => n1686, B2 => n961
                           , ZN => n8673);
   U1813 : OAI22_X1 port map( A1 => n1733, A2 => n1868, B1 => n1686, B2 => n962
                           , ZN => n8672);
   U1814 : OAI22_X1 port map( A1 => n1726, A2 => n1868, B1 => n1686, B2 => n963
                           , ZN => n8671);
   U1815 : OAI22_X1 port map( A1 => n1727, A2 => n1868, B1 => n1686, B2 => n964
                           , ZN => n8670);
   U1816 : OAI22_X1 port map( A1 => n1728, A2 => n1868, B1 => n1686, B2 => n965
                           , ZN => n8669);
   U1817 : OAI22_X1 port map( A1 => n1729, A2 => n1868, B1 => n1686, B2 => n966
                           , ZN => n8668);
   U1818 : OAI22_X1 port map( A1 => n1725, A2 => n1868, B1 => n1686, B2 => n967
                           , ZN => n8667);
   U1819 : OAI22_X1 port map( A1 => n1768, A2 => n1868, B1 => n1686, B2 => n968
                           , ZN => n8666);
   U1820 : OAI21_X1 port map( B1 => n1769, B2 => n1868, A => n1770, ZN => n1869
                           );
   U1821 : OAI22_X1 port map( A1 => n1759, A2 => n1870, B1 => n1688, B2 => 
                           n1289, ZN => n8665);
   U1822 : OAI22_X1 port map( A1 => n1761, A2 => n1870, B1 => n1688, B2 => 
                           n1290, ZN => n8664);
   U1823 : OAI22_X1 port map( A1 => n1762, A2 => n1870, B1 => n1688, B2 => 
                           n1291, ZN => n8663);
   U1824 : OAI22_X1 port map( A1 => n1763, A2 => n1870, B1 => n1688, B2 => 
                           n1292, ZN => n8662);
   U1825 : OAI22_X1 port map( A1 => n1764, A2 => n1870, B1 => n1688, B2 => 
                           n1293, ZN => n8661);
   U1826 : OAI22_X1 port map( A1 => n1765, A2 => n1870, B1 => n1688, B2 => 
                           n1294, ZN => n8660);
   U1827 : OAI22_X1 port map( A1 => n1766, A2 => n1870, B1 => n1688, B2 => 
                           n1295, ZN => n8659);
   U1828 : OAI22_X1 port map( A1 => n1767, A2 => n1870, B1 => n1688, B2 => 
                           n1296, ZN => n8658);
   U1829 : OAI22_X1 port map( A1 => n1746, A2 => n1870, B1 => n1688, B2 => 
                           n1297, ZN => n8657);
   U1830 : OAI22_X1 port map( A1 => n1747, A2 => n1870, B1 => n1688, B2 => 
                           n1298, ZN => n8656);
   U1831 : OAI22_X1 port map( A1 => n1742, A2 => n1870, B1 => n1688, B2 => 
                           n1299, ZN => n8655);
   U1832 : OAI22_X1 port map( A1 => n1743, A2 => n1870, B1 => n1688, B2 => 
                           n1300, ZN => n8654);
   U1833 : OAI22_X1 port map( A1 => n1744, A2 => n1870, B1 => n1688, B2 => 
                           n1301, ZN => n8653);
   U1834 : OAI22_X1 port map( A1 => n1745, A2 => n1870, B1 => n1688, B2 => 
                           n1302, ZN => n8652);
   U1835 : OAI22_X1 port map( A1 => n1738, A2 => n1870, B1 => n1688, B2 => 
                           n1303, ZN => n8651);
   U1836 : OAI22_X1 port map( A1 => n1739, A2 => n1870, B1 => n1688, B2 => 
                           n1304, ZN => n8650);
   U1837 : OAI22_X1 port map( A1 => n1740, A2 => n1870, B1 => n1688, B2 => 
                           n1305, ZN => n8649);
   U1838 : OAI22_X1 port map( A1 => n1741, A2 => n1870, B1 => n1688, B2 => 
                           n1306, ZN => n8648);
   U1839 : OAI22_X1 port map( A1 => n1734, A2 => n1870, B1 => n1688, B2 => 
                           n1307, ZN => n8647);
   U1840 : OAI22_X1 port map( A1 => n1735, A2 => n1870, B1 => n1688, B2 => 
                           n1308, ZN => n8646);
   U1841 : OAI22_X1 port map( A1 => n1736, A2 => n1870, B1 => n1688, B2 => 
                           n1309, ZN => n8645);
   U1842 : OAI22_X1 port map( A1 => n1737, A2 => n1870, B1 => n1688, B2 => 
                           n1310, ZN => n8644);
   U1843 : OAI22_X1 port map( A1 => n1730, A2 => n1870, B1 => n1688, B2 => 
                           n1311, ZN => n8643);
   U1844 : OAI22_X1 port map( A1 => n1731, A2 => n1870, B1 => n1688, B2 => 
                           n1312, ZN => n8642);
   U1845 : OAI22_X1 port map( A1 => n1732, A2 => n1870, B1 => n1688, B2 => 
                           n1313, ZN => n8641);
   U1846 : OAI22_X1 port map( A1 => n1733, A2 => n1870, B1 => n1688, B2 => 
                           n1314, ZN => n8640);
   U1847 : OAI22_X1 port map( A1 => n1726, A2 => n1870, B1 => n1688, B2 => 
                           n1315, ZN => n8639);
   U1848 : OAI22_X1 port map( A1 => n1727, A2 => n1870, B1 => n1688, B2 => 
                           n1316, ZN => n8638);
   U1849 : OAI22_X1 port map( A1 => n1728, A2 => n1870, B1 => n1688, B2 => 
                           n1317, ZN => n8637);
   U1850 : OAI22_X1 port map( A1 => n1729, A2 => n1870, B1 => n1688, B2 => 
                           n1318, ZN => n8636);
   U1851 : OAI22_X1 port map( A1 => n1725, A2 => n1870, B1 => n1688, B2 => 
                           n1319, ZN => n8635);
   U1852 : OAI22_X1 port map( A1 => n1768, A2 => n1870, B1 => n1688, B2 => 
                           n1320, ZN => n8634);
   U1853 : OAI21_X1 port map( B1 => n1769, B2 => n1870, A => n1770, ZN => n1871
                           );
   U1854 : OAI22_X1 port map( A1 => n1759, A2 => n1872, B1 => n4993, B2 => 
                           n1614, ZN => n8633);
   U1855 : OAI22_X1 port map( A1 => n1761, A2 => n1872, B1 => n4992, B2 => 
                           n1614, ZN => n8632);
   U1856 : OAI22_X1 port map( A1 => n1762, A2 => n1872, B1 => n4991, B2 => 
                           n1614, ZN => n8631);
   U1857 : OAI22_X1 port map( A1 => n1763, A2 => n1872, B1 => n4990, B2 => 
                           n1614, ZN => n8630);
   U1858 : OAI22_X1 port map( A1 => n1764, A2 => n1872, B1 => n4989, B2 => 
                           n1614, ZN => n8629);
   U1859 : OAI22_X1 port map( A1 => n1765, A2 => n1872, B1 => n4988, B2 => 
                           n1614, ZN => n8628);
   U1860 : OAI22_X1 port map( A1 => n1766, A2 => n1872, B1 => n4987, B2 => 
                           n1614, ZN => n8627);
   U1861 : OAI22_X1 port map( A1 => n1767, A2 => n1872, B1 => n4986, B2 => 
                           n1614, ZN => n8626);
   U1862 : OAI22_X1 port map( A1 => n1746, A2 => n1872, B1 => n4985, B2 => 
                           n1614, ZN => n8625);
   U1863 : OAI22_X1 port map( A1 => n1747, A2 => n1872, B1 => n4984, B2 => 
                           n1614, ZN => n8624);
   U1864 : OAI22_X1 port map( A1 => n1742, A2 => n1872, B1 => n4983, B2 => 
                           n1614, ZN => n8623);
   U1865 : OAI22_X1 port map( A1 => n1743, A2 => n1872, B1 => n4982, B2 => 
                           n1614, ZN => n8622);
   U1866 : OAI22_X1 port map( A1 => n1744, A2 => n1872, B1 => n4981, B2 => 
                           n1614, ZN => n8621);
   U1867 : OAI22_X1 port map( A1 => n1745, A2 => n1872, B1 => n4980, B2 => 
                           n1614, ZN => n8620);
   U1868 : OAI22_X1 port map( A1 => n1738, A2 => n1872, B1 => n4979, B2 => 
                           n1614, ZN => n8619);
   U1869 : OAI22_X1 port map( A1 => n1739, A2 => n1872, B1 => n4978, B2 => 
                           n1614, ZN => n8618);
   U1870 : OAI22_X1 port map( A1 => n1740, A2 => n1872, B1 => n4977, B2 => 
                           n1614, ZN => n8617);
   U1871 : OAI22_X1 port map( A1 => n1741, A2 => n1872, B1 => n4976, B2 => 
                           n1614, ZN => n8616);
   U1872 : OAI22_X1 port map( A1 => n1734, A2 => n1872, B1 => n4975, B2 => 
                           n1614, ZN => n8615);
   U1873 : OAI22_X1 port map( A1 => n1735, A2 => n1872, B1 => n4974, B2 => 
                           n1614, ZN => n8614);
   U1874 : OAI22_X1 port map( A1 => n1736, A2 => n1872, B1 => n4973, B2 => 
                           n1614, ZN => n8613);
   U1875 : OAI22_X1 port map( A1 => n1737, A2 => n1872, B1 => n4972, B2 => 
                           n1614, ZN => n8612);
   U1876 : OAI22_X1 port map( A1 => n1730, A2 => n1872, B1 => n4971, B2 => 
                           n1614, ZN => n8611);
   U1877 : OAI22_X1 port map( A1 => n1731, A2 => n1872, B1 => n4970, B2 => 
                           n1614, ZN => n8610);
   U1878 : OAI22_X1 port map( A1 => n1732, A2 => n1872, B1 => n4969, B2 => 
                           n1614, ZN => n8609);
   U1879 : OAI22_X1 port map( A1 => n1733, A2 => n1872, B1 => n4968, B2 => 
                           n1614, ZN => n8608);
   U1880 : OAI22_X1 port map( A1 => n1726, A2 => n1872, B1 => n4967, B2 => 
                           n1614, ZN => n8607);
   U1881 : OAI22_X1 port map( A1 => n1727, A2 => n1872, B1 => n4966, B2 => 
                           n1614, ZN => n8606);
   U1882 : OAI22_X1 port map( A1 => n1728, A2 => n1872, B1 => n4965, B2 => 
                           n1614, ZN => n8605);
   U1883 : OAI22_X1 port map( A1 => n1729, A2 => n1872, B1 => n4964, B2 => 
                           n1614, ZN => n8604);
   U1884 : OAI22_X1 port map( A1 => n1725, A2 => n1872, B1 => n4963, B2 => 
                           n1614, ZN => n8603);
   U1885 : OAI22_X1 port map( A1 => n1768, A2 => n1872, B1 => n4962, B2 => 
                           n1614, ZN => n8602);
   U1886 : OAI21_X1 port map( B1 => n1769, B2 => n1872, A => n1770, ZN => n1873
                           );
   U1887 : OAI22_X1 port map( A1 => n1759, A2 => n1874, B1 => n4961, B2 => 
                           n1616, ZN => n8601);
   U1888 : OAI22_X1 port map( A1 => n1761, A2 => n1874, B1 => n4960, B2 => 
                           n1616, ZN => n8600);
   U1889 : OAI22_X1 port map( A1 => n1762, A2 => n1874, B1 => n4959, B2 => 
                           n1616, ZN => n8599);
   U1890 : OAI22_X1 port map( A1 => n1763, A2 => n1874, B1 => n4958, B2 => 
                           n1616, ZN => n8598);
   U1891 : OAI22_X1 port map( A1 => n1764, A2 => n1874, B1 => n4957, B2 => 
                           n1616, ZN => n8597);
   U1892 : OAI22_X1 port map( A1 => n1765, A2 => n1874, B1 => n4956, B2 => 
                           n1616, ZN => n8596);
   U1893 : OAI22_X1 port map( A1 => n1766, A2 => n1874, B1 => n4955, B2 => 
                           n1616, ZN => n8595);
   U1894 : OAI22_X1 port map( A1 => n1767, A2 => n1874, B1 => n4954, B2 => 
                           n1616, ZN => n8594);
   U1895 : OAI22_X1 port map( A1 => n1746, A2 => n1874, B1 => n4953, B2 => 
                           n1616, ZN => n8593);
   U1896 : OAI22_X1 port map( A1 => n1747, A2 => n1874, B1 => n4952, B2 => 
                           n1616, ZN => n8592);
   U1897 : OAI22_X1 port map( A1 => n1742, A2 => n1874, B1 => n4951, B2 => 
                           n1616, ZN => n8591);
   U1898 : OAI22_X1 port map( A1 => n1743, A2 => n1874, B1 => n4950, B2 => 
                           n1616, ZN => n8590);
   U1899 : OAI22_X1 port map( A1 => n1744, A2 => n1874, B1 => n4949, B2 => 
                           n1616, ZN => n8589);
   U1900 : OAI22_X1 port map( A1 => n1745, A2 => n1874, B1 => n4948, B2 => 
                           n1616, ZN => n8588);
   U1901 : OAI22_X1 port map( A1 => n1738, A2 => n1874, B1 => n4947, B2 => 
                           n1616, ZN => n8587);
   U1902 : OAI22_X1 port map( A1 => n1739, A2 => n1874, B1 => n4946, B2 => 
                           n1616, ZN => n8586);
   U1903 : OAI22_X1 port map( A1 => n1740, A2 => n1874, B1 => n4945, B2 => 
                           n1616, ZN => n8585);
   U1904 : OAI22_X1 port map( A1 => n1741, A2 => n1874, B1 => n4944, B2 => 
                           n1616, ZN => n8584);
   U1905 : OAI22_X1 port map( A1 => n1734, A2 => n1874, B1 => n4943, B2 => 
                           n1616, ZN => n8583);
   U1906 : OAI22_X1 port map( A1 => n1735, A2 => n1874, B1 => n4942, B2 => 
                           n1616, ZN => n8582);
   U1907 : OAI22_X1 port map( A1 => n1736, A2 => n1874, B1 => n4941, B2 => 
                           n1616, ZN => n8581);
   U1908 : OAI22_X1 port map( A1 => n1737, A2 => n1874, B1 => n4940, B2 => 
                           n1616, ZN => n8580);
   U1909 : OAI22_X1 port map( A1 => n1730, A2 => n1874, B1 => n4939, B2 => 
                           n1616, ZN => n8579);
   U1910 : OAI22_X1 port map( A1 => n1731, A2 => n1874, B1 => n4938, B2 => 
                           n1616, ZN => n8578);
   U1911 : OAI22_X1 port map( A1 => n1732, A2 => n1874, B1 => n4937, B2 => 
                           n1616, ZN => n8577);
   U1912 : OAI22_X1 port map( A1 => n1733, A2 => n1874, B1 => n4936, B2 => 
                           n1616, ZN => n8576);
   U1913 : OAI22_X1 port map( A1 => n1726, A2 => n1874, B1 => n4935, B2 => 
                           n1616, ZN => n8575);
   U1914 : OAI22_X1 port map( A1 => n1727, A2 => n1874, B1 => n4934, B2 => 
                           n1616, ZN => n8574);
   U1915 : OAI22_X1 port map( A1 => n1728, A2 => n1874, B1 => n4933, B2 => 
                           n1616, ZN => n8573);
   U1916 : OAI22_X1 port map( A1 => n1729, A2 => n1874, B1 => n4932, B2 => 
                           n1616, ZN => n8572);
   U1917 : OAI22_X1 port map( A1 => n1725, A2 => n1874, B1 => n4931, B2 => 
                           n1616, ZN => n8571);
   U1918 : OAI22_X1 port map( A1 => n1768, A2 => n1874, B1 => n4930, B2 => 
                           n1616, ZN => n8570);
   U1919 : OAI21_X1 port map( B1 => n1769, B2 => n1874, A => n1770, ZN => n1875
                           );
   U1920 : OAI22_X1 port map( A1 => n1759, A2 => n1876, B1 => n4929, B2 => 
                           n1610, ZN => n8569);
   U1921 : OAI22_X1 port map( A1 => n1761, A2 => n1876, B1 => n4928, B2 => 
                           n1610, ZN => n8568);
   U1922 : OAI22_X1 port map( A1 => n1762, A2 => n1876, B1 => n4927, B2 => 
                           n1610, ZN => n8567);
   U1923 : OAI22_X1 port map( A1 => n1763, A2 => n1876, B1 => n4926, B2 => 
                           n1610, ZN => n8566);
   U1924 : OAI22_X1 port map( A1 => n1764, A2 => n1876, B1 => n4925, B2 => 
                           n1610, ZN => n8565);
   U1925 : OAI22_X1 port map( A1 => n1765, A2 => n1876, B1 => n4924, B2 => 
                           n1610, ZN => n8564);
   U1926 : OAI22_X1 port map( A1 => n1766, A2 => n1876, B1 => n4923, B2 => 
                           n1610, ZN => n8563);
   U1927 : OAI22_X1 port map( A1 => n1767, A2 => n1876, B1 => n4922, B2 => 
                           n1610, ZN => n8562);
   U1928 : OAI22_X1 port map( A1 => n1746, A2 => n1876, B1 => n4921, B2 => 
                           n1610, ZN => n8561);
   U1929 : OAI22_X1 port map( A1 => n1747, A2 => n1876, B1 => n4920, B2 => 
                           n1610, ZN => n8560);
   U1930 : OAI22_X1 port map( A1 => n1742, A2 => n1876, B1 => n4919, B2 => 
                           n1610, ZN => n8559);
   U1931 : OAI22_X1 port map( A1 => n1743, A2 => n1876, B1 => n4918, B2 => 
                           n1610, ZN => n8558);
   U1932 : OAI22_X1 port map( A1 => n1744, A2 => n1876, B1 => n4917, B2 => 
                           n1610, ZN => n8557);
   U1933 : OAI22_X1 port map( A1 => n1745, A2 => n1876, B1 => n4916, B2 => 
                           n1610, ZN => n8556);
   U1934 : OAI22_X1 port map( A1 => n1738, A2 => n1876, B1 => n4915, B2 => 
                           n1610, ZN => n8555);
   U1935 : OAI22_X1 port map( A1 => n1739, A2 => n1876, B1 => n4914, B2 => 
                           n1610, ZN => n8554);
   U1936 : OAI22_X1 port map( A1 => n1740, A2 => n1876, B1 => n4913, B2 => 
                           n1610, ZN => n8553);
   U1937 : OAI22_X1 port map( A1 => n1741, A2 => n1876, B1 => n4912, B2 => 
                           n1610, ZN => n8552);
   U1938 : OAI22_X1 port map( A1 => n1734, A2 => n1876, B1 => n4911, B2 => 
                           n1610, ZN => n8551);
   U1939 : OAI22_X1 port map( A1 => n1735, A2 => n1876, B1 => n4910, B2 => 
                           n1610, ZN => n8550);
   U1940 : OAI22_X1 port map( A1 => n1736, A2 => n1876, B1 => n4909, B2 => 
                           n1610, ZN => n8549);
   U1941 : OAI22_X1 port map( A1 => n1737, A2 => n1876, B1 => n4908, B2 => 
                           n1610, ZN => n8548);
   U1942 : OAI22_X1 port map( A1 => n1730, A2 => n1876, B1 => n4907, B2 => 
                           n1610, ZN => n8547);
   U1943 : OAI22_X1 port map( A1 => n1731, A2 => n1876, B1 => n4906, B2 => 
                           n1610, ZN => n8546);
   U1944 : OAI22_X1 port map( A1 => n1732, A2 => n1876, B1 => n4905, B2 => 
                           n1610, ZN => n8545);
   U1945 : OAI22_X1 port map( A1 => n1733, A2 => n1876, B1 => n4904, B2 => 
                           n1610, ZN => n8544);
   U1946 : OAI22_X1 port map( A1 => n1726, A2 => n1876, B1 => n4903, B2 => 
                           n1610, ZN => n8543);
   U1947 : OAI22_X1 port map( A1 => n1727, A2 => n1876, B1 => n4902, B2 => 
                           n1610, ZN => n8542);
   U1948 : OAI22_X1 port map( A1 => n1728, A2 => n1876, B1 => n4901, B2 => 
                           n1610, ZN => n8541);
   U1949 : OAI22_X1 port map( A1 => n1729, A2 => n1876, B1 => n4900, B2 => 
                           n1610, ZN => n8540);
   U1950 : OAI22_X1 port map( A1 => n1725, A2 => n1876, B1 => n4899, B2 => 
                           n1610, ZN => n8539);
   U1951 : OAI22_X1 port map( A1 => n1768, A2 => n1876, B1 => n4898, B2 => 
                           n1610, ZN => n8538);
   U1952 : OAI21_X1 port map( B1 => n1769, B2 => n1876, A => n1770, ZN => n1877
                           );
   U1953 : OAI22_X1 port map( A1 => n1759, A2 => n1878, B1 => n1682, B2 => n619
                           , ZN => n8537);
   U1954 : OAI22_X1 port map( A1 => n1761, A2 => n1878, B1 => n1682, B2 => n622
                           , ZN => n8536);
   U1955 : OAI22_X1 port map( A1 => n1762, A2 => n1878, B1 => n1682, B2 => n625
                           , ZN => n8535);
   U1956 : OAI22_X1 port map( A1 => n1763, A2 => n1878, B1 => n1682, B2 => n628
                           , ZN => n8534);
   U1957 : OAI22_X1 port map( A1 => n1764, A2 => n1878, B1 => n1682, B2 => n631
                           , ZN => n8533);
   U1958 : OAI22_X1 port map( A1 => n1765, A2 => n1878, B1 => n1682, B2 => n634
                           , ZN => n8532);
   U1959 : OAI22_X1 port map( A1 => n1766, A2 => n1878, B1 => n1682, B2 => n637
                           , ZN => n8531);
   U1960 : OAI22_X1 port map( A1 => n1767, A2 => n1878, B1 => n1682, B2 => n640
                           , ZN => n8530);
   U1961 : OAI22_X1 port map( A1 => n1746, A2 => n1878, B1 => n1682, B2 => n643
                           , ZN => n8529);
   U1962 : OAI22_X1 port map( A1 => n1747, A2 => n1878, B1 => n1682, B2 => n646
                           , ZN => n8528);
   U1963 : OAI22_X1 port map( A1 => n1742, A2 => n1878, B1 => n1682, B2 => n649
                           , ZN => n8527);
   U1964 : OAI22_X1 port map( A1 => n1743, A2 => n1878, B1 => n1682, B2 => n652
                           , ZN => n8526);
   U1965 : OAI22_X1 port map( A1 => n1744, A2 => n1878, B1 => n1682, B2 => n655
                           , ZN => n8525);
   U1966 : OAI22_X1 port map( A1 => n1745, A2 => n1878, B1 => n1682, B2 => n658
                           , ZN => n8524);
   U1967 : OAI22_X1 port map( A1 => n1738, A2 => n1878, B1 => n1682, B2 => n661
                           , ZN => n8523);
   U1968 : OAI22_X1 port map( A1 => n1739, A2 => n1878, B1 => n1682, B2 => n664
                           , ZN => n8522);
   U1969 : OAI22_X1 port map( A1 => n1740, A2 => n1878, B1 => n1682, B2 => n667
                           , ZN => n8521);
   U1970 : OAI22_X1 port map( A1 => n1741, A2 => n1878, B1 => n1682, B2 => n670
                           , ZN => n8520);
   U1971 : OAI22_X1 port map( A1 => n1734, A2 => n1878, B1 => n1682, B2 => n673
                           , ZN => n8519);
   U1972 : OAI22_X1 port map( A1 => n1735, A2 => n1878, B1 => n1682, B2 => n676
                           , ZN => n8518);
   U1973 : OAI22_X1 port map( A1 => n1736, A2 => n1878, B1 => n1682, B2 => n679
                           , ZN => n8517);
   U1974 : OAI22_X1 port map( A1 => n1737, A2 => n1878, B1 => n1682, B2 => n682
                           , ZN => n8516);
   U1975 : OAI22_X1 port map( A1 => n1730, A2 => n1878, B1 => n1682, B2 => n685
                           , ZN => n8515);
   U1976 : OAI22_X1 port map( A1 => n1731, A2 => n1878, B1 => n1682, B2 => n688
                           , ZN => n8514);
   U1977 : OAI22_X1 port map( A1 => n1732, A2 => n1878, B1 => n1682, B2 => n691
                           , ZN => n8513);
   U1978 : OAI22_X1 port map( A1 => n1733, A2 => n1878, B1 => n1682, B2 => n694
                           , ZN => n8512);
   U1979 : OAI22_X1 port map( A1 => n1726, A2 => n1878, B1 => n1682, B2 => n697
                           , ZN => n8511);
   U1980 : OAI22_X1 port map( A1 => n1727, A2 => n1878, B1 => n1682, B2 => n700
                           , ZN => n8510);
   U1981 : OAI22_X1 port map( A1 => n1728, A2 => n1878, B1 => n1682, B2 => n703
                           , ZN => n8509);
   U1982 : OAI22_X1 port map( A1 => n1729, A2 => n1878, B1 => n1682, B2 => n706
                           , ZN => n8508);
   U1983 : OAI22_X1 port map( A1 => n1725, A2 => n1878, B1 => n1682, B2 => n709
                           , ZN => n8507);
   U1984 : OAI22_X1 port map( A1 => n1768, A2 => n1878, B1 => n1682, B2 => n712
                           , ZN => n8506);
   U1985 : OAI21_X1 port map( B1 => n1769, B2 => n1878, A => n1770, ZN => n1879
                           );
   U1986 : OAI22_X1 port map( A1 => n1759, A2 => n1880, B1 => n1684, B2 => n195
                           , ZN => n8505);
   U1987 : OAI22_X1 port map( A1 => n1761, A2 => n1880, B1 => n1684, B2 => n198
                           , ZN => n8504);
   U1988 : OAI22_X1 port map( A1 => n1762, A2 => n1880, B1 => n1684, B2 => n201
                           , ZN => n8503);
   U1989 : OAI22_X1 port map( A1 => n1763, A2 => n1880, B1 => n1684, B2 => n204
                           , ZN => n8502);
   U1990 : OAI22_X1 port map( A1 => n1764, A2 => n1880, B1 => n1684, B2 => n207
                           , ZN => n8501);
   U1991 : OAI22_X1 port map( A1 => n1765, A2 => n1880, B1 => n1684, B2 => n210
                           , ZN => n8500);
   U1992 : OAI22_X1 port map( A1 => n1766, A2 => n1880, B1 => n1684, B2 => n213
                           , ZN => n8499);
   U1993 : OAI22_X1 port map( A1 => n1767, A2 => n1880, B1 => n1684, B2 => n216
                           , ZN => n8498);
   U1994 : OAI22_X1 port map( A1 => n1746, A2 => n1880, B1 => n1684, B2 => n219
                           , ZN => n8497);
   U1995 : OAI22_X1 port map( A1 => n1747, A2 => n1880, B1 => n1684, B2 => n222
                           , ZN => n8496);
   U1996 : OAI22_X1 port map( A1 => n1742, A2 => n1880, B1 => n1684, B2 => n225
                           , ZN => n8495);
   U1997 : OAI22_X1 port map( A1 => n1743, A2 => n1880, B1 => n1684, B2 => n228
                           , ZN => n8494);
   U1998 : OAI22_X1 port map( A1 => n1744, A2 => n1880, B1 => n1684, B2 => n231
                           , ZN => n8493);
   U1999 : OAI22_X1 port map( A1 => n1745, A2 => n1880, B1 => n1684, B2 => n234
                           , ZN => n8492);
   U2000 : OAI22_X1 port map( A1 => n1738, A2 => n1880, B1 => n1684, B2 => n237
                           , ZN => n8491);
   U2001 : OAI22_X1 port map( A1 => n1739, A2 => n1880, B1 => n1684, B2 => n240
                           , ZN => n8490);
   U2002 : OAI22_X1 port map( A1 => n1740, A2 => n1880, B1 => n1684, B2 => n243
                           , ZN => n8489);
   U2003 : OAI22_X1 port map( A1 => n1741, A2 => n1880, B1 => n1684, B2 => n246
                           , ZN => n8488);
   U2004 : OAI22_X1 port map( A1 => n1734, A2 => n1880, B1 => n1684, B2 => n249
                           , ZN => n8487);
   U2005 : OAI22_X1 port map( A1 => n1735, A2 => n1880, B1 => n1684, B2 => n252
                           , ZN => n8486);
   U2006 : OAI22_X1 port map( A1 => n1736, A2 => n1880, B1 => n1684, B2 => n255
                           , ZN => n8485);
   U2007 : OAI22_X1 port map( A1 => n1737, A2 => n1880, B1 => n1684, B2 => n258
                           , ZN => n8484);
   U2008 : OAI22_X1 port map( A1 => n1730, A2 => n1880, B1 => n1684, B2 => n261
                           , ZN => n8483);
   U2009 : OAI22_X1 port map( A1 => n1731, A2 => n1880, B1 => n1684, B2 => n264
                           , ZN => n8482);
   U2010 : OAI22_X1 port map( A1 => n1732, A2 => n1880, B1 => n1684, B2 => n267
                           , ZN => n8481);
   U2011 : OAI22_X1 port map( A1 => n1733, A2 => n1880, B1 => n1684, B2 => n270
                           , ZN => n8480);
   U2012 : OAI22_X1 port map( A1 => n1726, A2 => n1880, B1 => n1684, B2 => n273
                           , ZN => n8479);
   U2013 : OAI22_X1 port map( A1 => n1727, A2 => n1880, B1 => n1684, B2 => n276
                           , ZN => n8478);
   U2014 : OAI22_X1 port map( A1 => n1728, A2 => n1880, B1 => n1684, B2 => n279
                           , ZN => n8477);
   U2015 : OAI22_X1 port map( A1 => n1729, A2 => n1880, B1 => n1684, B2 => n282
                           , ZN => n8476);
   U2016 : OAI22_X1 port map( A1 => n1725, A2 => n1880, B1 => n1684, B2 => n285
                           , ZN => n8475);
   U2017 : OAI22_X1 port map( A1 => n1768, A2 => n1880, B1 => n1684, B2 => n288
                           , ZN => n8474);
   U2018 : OAI21_X1 port map( B1 => n1769, B2 => n1880, A => n1770, ZN => n1881
                           );
   U2019 : OAI22_X1 port map( A1 => n1759, A2 => n1882, B1 => n5690, B2 => 
                           n1612, ZN => n8473);
   U2020 : OAI22_X1 port map( A1 => n1761, A2 => n1882, B1 => n5680, B2 => 
                           n1612, ZN => n8472);
   U2021 : OAI22_X1 port map( A1 => n1762, A2 => n1882, B1 => n5670, B2 => 
                           n1612, ZN => n8471);
   U2022 : OAI22_X1 port map( A1 => n1763, A2 => n1882, B1 => n5660, B2 => 
                           n1612, ZN => n8470);
   U2023 : OAI22_X1 port map( A1 => n1764, A2 => n1882, B1 => n5650, B2 => 
                           n1612, ZN => n8469);
   U2024 : OAI22_X1 port map( A1 => n1765, A2 => n1882, B1 => n5640, B2 => 
                           n1612, ZN => n8468);
   U2025 : OAI22_X1 port map( A1 => n1766, A2 => n1882, B1 => n5630, B2 => 
                           n1612, ZN => n8467);
   U2026 : OAI22_X1 port map( A1 => n1767, A2 => n1882, B1 => n5620, B2 => 
                           n1612, ZN => n8466);
   U2027 : OAI22_X1 port map( A1 => n1746, A2 => n1882, B1 => n5610, B2 => 
                           n1612, ZN => n8465);
   U2028 : OAI22_X1 port map( A1 => n1747, A2 => n1882, B1 => n5600, B2 => 
                           n1612, ZN => n8464);
   U2029 : OAI22_X1 port map( A1 => n1742, A2 => n1882, B1 => n5590, B2 => 
                           n1612, ZN => n8463);
   U2030 : OAI22_X1 port map( A1 => n1743, A2 => n1882, B1 => n5580, B2 => 
                           n1612, ZN => n8462);
   U2031 : OAI22_X1 port map( A1 => n1744, A2 => n1882, B1 => n5570, B2 => 
                           n1612, ZN => n8461);
   U2032 : OAI22_X1 port map( A1 => n1745, A2 => n1882, B1 => n5560, B2 => 
                           n1612, ZN => n8460);
   U2033 : OAI22_X1 port map( A1 => n1738, A2 => n1882, B1 => n5550, B2 => 
                           n1612, ZN => n8459);
   U2034 : OAI22_X1 port map( A1 => n1739, A2 => n1882, B1 => n5540, B2 => 
                           n1612, ZN => n8458);
   U2035 : OAI22_X1 port map( A1 => n1740, A2 => n1882, B1 => n5530, B2 => 
                           n1612, ZN => n8457);
   U2036 : OAI22_X1 port map( A1 => n1741, A2 => n1882, B1 => n5520, B2 => 
                           n1612, ZN => n8456);
   U2037 : OAI22_X1 port map( A1 => n1734, A2 => n1882, B1 => n5510, B2 => 
                           n1612, ZN => n8455);
   U2038 : OAI22_X1 port map( A1 => n1735, A2 => n1882, B1 => n5500, B2 => 
                           n1612, ZN => n8454);
   U2039 : OAI22_X1 port map( A1 => n1736, A2 => n1882, B1 => n5490, B2 => 
                           n1612, ZN => n8453);
   U2040 : OAI22_X1 port map( A1 => n1737, A2 => n1882, B1 => n5480, B2 => 
                           n1612, ZN => n8452);
   U2041 : OAI22_X1 port map( A1 => n1730, A2 => n1882, B1 => n5470, B2 => 
                           n1612, ZN => n8451);
   U2042 : OAI22_X1 port map( A1 => n1731, A2 => n1882, B1 => n5460, B2 => 
                           n1612, ZN => n8450);
   U2043 : OAI22_X1 port map( A1 => n1732, A2 => n1882, B1 => n5450, B2 => 
                           n1612, ZN => n8449);
   U2044 : OAI22_X1 port map( A1 => n1733, A2 => n1882, B1 => n5440, B2 => 
                           n1612, ZN => n8448);
   U2045 : OAI22_X1 port map( A1 => n1726, A2 => n1882, B1 => n5430, B2 => 
                           n1612, ZN => n8447);
   U2046 : OAI22_X1 port map( A1 => n1727, A2 => n1882, B1 => n5420, B2 => 
                           n1612, ZN => n8446);
   U2047 : OAI22_X1 port map( A1 => n1728, A2 => n1882, B1 => n5410, B2 => 
                           n1612, ZN => n8445);
   U2048 : OAI22_X1 port map( A1 => n1729, A2 => n1882, B1 => n5400, B2 => 
                           n1612, ZN => n8444);
   U2049 : OAI22_X1 port map( A1 => n1725, A2 => n1882, B1 => n5390, B2 => 
                           n1612, ZN => n8443);
   U2050 : OAI22_X1 port map( A1 => n1768, A2 => n1882, B1 => n5380, B2 => 
                           n1612, ZN => n8442);
   U2051 : OAI21_X1 port map( B1 => n1769, B2 => n1882, A => n1770, ZN => n1883
                           );
   U2052 : OAI22_X1 port map( A1 => n1759, A2 => n1885, B1 => n5691, B2 => 
                           n1606, ZN => n8441);
   U2053 : OAI22_X1 port map( A1 => n1761, A2 => n1885, B1 => n5681, B2 => 
                           n1606, ZN => n8440);
   U2054 : OAI22_X1 port map( A1 => n1762, A2 => n1885, B1 => n5671, B2 => 
                           n1606, ZN => n8439);
   U2055 : OAI22_X1 port map( A1 => n1763, A2 => n1885, B1 => n5661, B2 => 
                           n1606, ZN => n8438);
   U2056 : OAI22_X1 port map( A1 => n1764, A2 => n1885, B1 => n5651, B2 => 
                           n1606, ZN => n8437);
   U2057 : OAI22_X1 port map( A1 => n1765, A2 => n1885, B1 => n5641, B2 => 
                           n1606, ZN => n8436);
   U2058 : OAI22_X1 port map( A1 => n1766, A2 => n1885, B1 => n5631, B2 => 
                           n1606, ZN => n8435);
   U2059 : OAI22_X1 port map( A1 => n1767, A2 => n1885, B1 => n5621, B2 => 
                           n1606, ZN => n8434);
   U2060 : OAI22_X1 port map( A1 => n1746, A2 => n1885, B1 => n5611, B2 => 
                           n1606, ZN => n8433);
   U2061 : OAI22_X1 port map( A1 => n1747, A2 => n1885, B1 => n5601, B2 => 
                           n1606, ZN => n8432);
   U2062 : OAI22_X1 port map( A1 => n1742, A2 => n1885, B1 => n5591, B2 => 
                           n1606, ZN => n8431);
   U2063 : OAI22_X1 port map( A1 => n1743, A2 => n1885, B1 => n5581, B2 => 
                           n1606, ZN => n8430);
   U2064 : OAI22_X1 port map( A1 => n1744, A2 => n1885, B1 => n5571, B2 => 
                           n1606, ZN => n8429);
   U2065 : OAI22_X1 port map( A1 => n1745, A2 => n1885, B1 => n5561, B2 => 
                           n1606, ZN => n8428);
   U2066 : OAI22_X1 port map( A1 => n1738, A2 => n1885, B1 => n5551, B2 => 
                           n1606, ZN => n8427);
   U2067 : OAI22_X1 port map( A1 => n1739, A2 => n1885, B1 => n5541, B2 => 
                           n1606, ZN => n8426);
   U2068 : OAI22_X1 port map( A1 => n1740, A2 => n1885, B1 => n5531, B2 => 
                           n1606, ZN => n8425);
   U2069 : OAI22_X1 port map( A1 => n1741, A2 => n1885, B1 => n5521, B2 => 
                           n1606, ZN => n8424);
   U2070 : OAI22_X1 port map( A1 => n1734, A2 => n1885, B1 => n5511, B2 => 
                           n1606, ZN => n8423);
   U2071 : OAI22_X1 port map( A1 => n1735, A2 => n1885, B1 => n5501, B2 => 
                           n1606, ZN => n8422);
   U2072 : OAI22_X1 port map( A1 => n1736, A2 => n1885, B1 => n5491, B2 => 
                           n1606, ZN => n8421);
   U2073 : OAI22_X1 port map( A1 => n1737, A2 => n1885, B1 => n5481, B2 => 
                           n1606, ZN => n8420);
   U2074 : OAI22_X1 port map( A1 => n1730, A2 => n1885, B1 => n5471, B2 => 
                           n1606, ZN => n8419);
   U2075 : OAI22_X1 port map( A1 => n1731, A2 => n1885, B1 => n5461, B2 => 
                           n1606, ZN => n8418);
   U2076 : OAI22_X1 port map( A1 => n1732, A2 => n1885, B1 => n5451, B2 => 
                           n1606, ZN => n8417);
   U2077 : OAI22_X1 port map( A1 => n1733, A2 => n1885, B1 => n5441, B2 => 
                           n1606, ZN => n8416);
   U2078 : OAI22_X1 port map( A1 => n1726, A2 => n1885, B1 => n5431, B2 => 
                           n1606, ZN => n8415);
   U2079 : OAI22_X1 port map( A1 => n1727, A2 => n1885, B1 => n5421, B2 => 
                           n1606, ZN => n8414);
   U2080 : OAI22_X1 port map( A1 => n1728, A2 => n1885, B1 => n5411, B2 => 
                           n1606, ZN => n8413);
   U2081 : OAI22_X1 port map( A1 => n1729, A2 => n1885, B1 => n5401, B2 => 
                           n1606, ZN => n8412);
   U2082 : OAI22_X1 port map( A1 => n1725, A2 => n1885, B1 => n5391, B2 => 
                           n1606, ZN => n8411);
   U2083 : OAI22_X1 port map( A1 => n1768, A2 => n1885, B1 => n5381, B2 => 
                           n1606, ZN => n8410);
   U2084 : OAI21_X1 port map( B1 => n1769, B2 => n1885, A => n1770, ZN => n1886
                           );
   U2085 : OAI22_X1 port map( A1 => n1759, A2 => n1888, B1 => n1678, B2 => n969
                           , ZN => n8409);
   U2086 : OAI22_X1 port map( A1 => n1761, A2 => n1888, B1 => n1678, B2 => n970
                           , ZN => n8408);
   U2087 : OAI22_X1 port map( A1 => n1762, A2 => n1888, B1 => n1678, B2 => n971
                           , ZN => n8407);
   U2088 : OAI22_X1 port map( A1 => n1763, A2 => n1888, B1 => n1678, B2 => n972
                           , ZN => n8406);
   U2089 : OAI22_X1 port map( A1 => n1764, A2 => n1888, B1 => n1678, B2 => n973
                           , ZN => n8405);
   U2090 : OAI22_X1 port map( A1 => n1765, A2 => n1888, B1 => n1678, B2 => n974
                           , ZN => n8404);
   U2091 : OAI22_X1 port map( A1 => n1766, A2 => n1888, B1 => n1678, B2 => n975
                           , ZN => n8403);
   U2092 : OAI22_X1 port map( A1 => n1767, A2 => n1888, B1 => n1678, B2 => n976
                           , ZN => n8402);
   U2093 : OAI22_X1 port map( A1 => n1746, A2 => n1888, B1 => n1678, B2 => n977
                           , ZN => n8401);
   U2094 : OAI22_X1 port map( A1 => n1747, A2 => n1888, B1 => n1678, B2 => n978
                           , ZN => n8400);
   U2095 : OAI22_X1 port map( A1 => n1742, A2 => n1888, B1 => n1678, B2 => n979
                           , ZN => n8399);
   U2096 : OAI22_X1 port map( A1 => n1743, A2 => n1888, B1 => n1678, B2 => n980
                           , ZN => n8398);
   U2097 : OAI22_X1 port map( A1 => n1744, A2 => n1888, B1 => n1678, B2 => n981
                           , ZN => n8397);
   U2098 : OAI22_X1 port map( A1 => n1745, A2 => n1888, B1 => n1678, B2 => n982
                           , ZN => n8396);
   U2099 : OAI22_X1 port map( A1 => n1738, A2 => n1888, B1 => n1678, B2 => n983
                           , ZN => n8395);
   U2100 : OAI22_X1 port map( A1 => n1739, A2 => n1888, B1 => n1678, B2 => n984
                           , ZN => n8394);
   U2101 : OAI22_X1 port map( A1 => n1740, A2 => n1888, B1 => n1678, B2 => n985
                           , ZN => n8393);
   U2102 : OAI22_X1 port map( A1 => n1741, A2 => n1888, B1 => n1678, B2 => n986
                           , ZN => n8392);
   U2103 : OAI22_X1 port map( A1 => n1734, A2 => n1888, B1 => n1678, B2 => n987
                           , ZN => n8391);
   U2104 : OAI22_X1 port map( A1 => n1735, A2 => n1888, B1 => n1678, B2 => n988
                           , ZN => n8390);
   U2105 : OAI22_X1 port map( A1 => n1736, A2 => n1888, B1 => n1678, B2 => n989
                           , ZN => n8389);
   U2106 : OAI22_X1 port map( A1 => n1737, A2 => n1888, B1 => n1678, B2 => n990
                           , ZN => n8388);
   U2107 : OAI22_X1 port map( A1 => n1730, A2 => n1888, B1 => n1678, B2 => n991
                           , ZN => n8387);
   U2108 : OAI22_X1 port map( A1 => n1731, A2 => n1888, B1 => n1678, B2 => n992
                           , ZN => n8386);
   U2109 : OAI22_X1 port map( A1 => n1732, A2 => n1888, B1 => n1678, B2 => n993
                           , ZN => n8385);
   U2110 : OAI22_X1 port map( A1 => n1733, A2 => n1888, B1 => n1678, B2 => n994
                           , ZN => n8384);
   U2111 : OAI22_X1 port map( A1 => n1726, A2 => n1888, B1 => n1678, B2 => n995
                           , ZN => n8383);
   U2112 : OAI22_X1 port map( A1 => n1727, A2 => n1888, B1 => n1678, B2 => n996
                           , ZN => n8382);
   U2113 : OAI22_X1 port map( A1 => n1728, A2 => n1888, B1 => n1678, B2 => n997
                           , ZN => n8381);
   U2114 : OAI22_X1 port map( A1 => n1729, A2 => n1888, B1 => n1678, B2 => n998
                           , ZN => n8380);
   U2115 : OAI22_X1 port map( A1 => n1725, A2 => n1888, B1 => n1678, B2 => n999
                           , ZN => n8379);
   U2116 : OAI22_X1 port map( A1 => n1768, A2 => n1888, B1 => n1678, B2 => 
                           n1000, ZN => n8378);
   U2117 : OAI21_X1 port map( B1 => n1769, B2 => n1888, A => n1770, ZN => n1889
                           );
   U2118 : OAI22_X1 port map( A1 => n1759, A2 => n1890, B1 => n1680, B2 => 
                           n1321, ZN => n8377);
   U2119 : OAI22_X1 port map( A1 => n1761, A2 => n1890, B1 => n1680, B2 => 
                           n1322, ZN => n8376);
   U2120 : OAI22_X1 port map( A1 => n1762, A2 => n1890, B1 => n1680, B2 => 
                           n1323, ZN => n8375);
   U2121 : OAI22_X1 port map( A1 => n1763, A2 => n1890, B1 => n1680, B2 => 
                           n1324, ZN => n8374);
   U2122 : OAI22_X1 port map( A1 => n1764, A2 => n1890, B1 => n1680, B2 => 
                           n1325, ZN => n8373);
   U2123 : OAI22_X1 port map( A1 => n1765, A2 => n1890, B1 => n1680, B2 => 
                           n1326, ZN => n8372);
   U2124 : OAI22_X1 port map( A1 => n1766, A2 => n1890, B1 => n1680, B2 => 
                           n1327, ZN => n8371);
   U2125 : OAI22_X1 port map( A1 => n1767, A2 => n1890, B1 => n1680, B2 => 
                           n1328, ZN => n8370);
   U2126 : OAI22_X1 port map( A1 => n1746, A2 => n1890, B1 => n1680, B2 => 
                           n1329, ZN => n8369);
   U2127 : OAI22_X1 port map( A1 => n1747, A2 => n1890, B1 => n1680, B2 => 
                           n1330, ZN => n8368);
   U2128 : OAI22_X1 port map( A1 => n1742, A2 => n1890, B1 => n1680, B2 => 
                           n1331, ZN => n8367);
   U2129 : OAI22_X1 port map( A1 => n1743, A2 => n1890, B1 => n1680, B2 => 
                           n1332, ZN => n8366);
   U2130 : OAI22_X1 port map( A1 => n1744, A2 => n1890, B1 => n1680, B2 => 
                           n1333, ZN => n8365);
   U2131 : OAI22_X1 port map( A1 => n1745, A2 => n1890, B1 => n1680, B2 => 
                           n1334, ZN => n8364);
   U2132 : OAI22_X1 port map( A1 => n1738, A2 => n1890, B1 => n1680, B2 => 
                           n1335, ZN => n8363);
   U2133 : OAI22_X1 port map( A1 => n1739, A2 => n1890, B1 => n1680, B2 => 
                           n1336, ZN => n8362);
   U2134 : OAI22_X1 port map( A1 => n1740, A2 => n1890, B1 => n1680, B2 => 
                           n1337, ZN => n8361);
   U2135 : OAI22_X1 port map( A1 => n1741, A2 => n1890, B1 => n1680, B2 => 
                           n1338, ZN => n8360);
   U2136 : OAI22_X1 port map( A1 => n1734, A2 => n1890, B1 => n1680, B2 => 
                           n1339, ZN => n8359);
   U2137 : OAI22_X1 port map( A1 => n1735, A2 => n1890, B1 => n1680, B2 => 
                           n1340, ZN => n8358);
   U2138 : OAI22_X1 port map( A1 => n1736, A2 => n1890, B1 => n1680, B2 => 
                           n1341, ZN => n8357);
   U2139 : OAI22_X1 port map( A1 => n1737, A2 => n1890, B1 => n1680, B2 => 
                           n1342, ZN => n8356);
   U2140 : OAI22_X1 port map( A1 => n1730, A2 => n1890, B1 => n1680, B2 => 
                           n1343, ZN => n8355);
   U2141 : OAI22_X1 port map( A1 => n1731, A2 => n1890, B1 => n1680, B2 => 
                           n1344, ZN => n8354);
   U2142 : OAI22_X1 port map( A1 => n1732, A2 => n1890, B1 => n1680, B2 => 
                           n1345, ZN => n8353);
   U2143 : OAI22_X1 port map( A1 => n1733, A2 => n1890, B1 => n1680, B2 => 
                           n1346, ZN => n8352);
   U2144 : OAI22_X1 port map( A1 => n1726, A2 => n1890, B1 => n1680, B2 => 
                           n1347, ZN => n8351);
   U2145 : OAI22_X1 port map( A1 => n1727, A2 => n1890, B1 => n1680, B2 => 
                           n1348, ZN => n8350);
   U2146 : OAI22_X1 port map( A1 => n1728, A2 => n1890, B1 => n1680, B2 => 
                           n1349, ZN => n8349);
   U2147 : OAI22_X1 port map( A1 => n1729, A2 => n1890, B1 => n1680, B2 => 
                           n1350, ZN => n8348);
   U2148 : OAI22_X1 port map( A1 => n1725, A2 => n1890, B1 => n1680, B2 => 
                           n1351, ZN => n8347);
   U2149 : OAI22_X1 port map( A1 => n1768, A2 => n1890, B1 => n1680, B2 => 
                           n1352, ZN => n8346);
   U2150 : OAI21_X1 port map( B1 => n1769, B2 => n1890, A => n1770, ZN => n1891
                           );
   U2151 : OAI22_X1 port map( A1 => n1759, A2 => n1892, B1 => n4897, B2 => 
                           n1608, ZN => n8345);
   U2152 : OAI22_X1 port map( A1 => n1761, A2 => n1892, B1 => n4896, B2 => 
                           n1608, ZN => n8344);
   U2153 : OAI22_X1 port map( A1 => n1762, A2 => n1892, B1 => n4895, B2 => 
                           n1608, ZN => n8343);
   U2154 : OAI22_X1 port map( A1 => n1763, A2 => n1892, B1 => n4894, B2 => 
                           n1608, ZN => n8342);
   U2155 : OAI22_X1 port map( A1 => n1764, A2 => n1892, B1 => n4893, B2 => 
                           n1608, ZN => n8341);
   U2156 : OAI22_X1 port map( A1 => n1765, A2 => n1892, B1 => n4892, B2 => 
                           n1608, ZN => n8340);
   U2157 : OAI22_X1 port map( A1 => n1766, A2 => n1892, B1 => n4891, B2 => 
                           n1608, ZN => n8339);
   U2158 : OAI22_X1 port map( A1 => n1767, A2 => n1892, B1 => n4890, B2 => 
                           n1608, ZN => n8338);
   U2159 : OAI22_X1 port map( A1 => n1746, A2 => n1892, B1 => n4889, B2 => 
                           n1608, ZN => n8337);
   U2160 : OAI22_X1 port map( A1 => n1747, A2 => n1892, B1 => n4888, B2 => 
                           n1608, ZN => n8336);
   U2161 : OAI22_X1 port map( A1 => n1742, A2 => n1892, B1 => n4887, B2 => 
                           n1608, ZN => n8335);
   U2162 : OAI22_X1 port map( A1 => n1743, A2 => n1892, B1 => n4886, B2 => 
                           n1608, ZN => n8334);
   U2163 : OAI22_X1 port map( A1 => n1744, A2 => n1892, B1 => n4885, B2 => 
                           n1608, ZN => n8333);
   U2164 : OAI22_X1 port map( A1 => n1745, A2 => n1892, B1 => n4884, B2 => 
                           n1608, ZN => n8332);
   U2165 : OAI22_X1 port map( A1 => n1738, A2 => n1892, B1 => n4883, B2 => 
                           n1608, ZN => n8331);
   U2166 : OAI22_X1 port map( A1 => n1739, A2 => n1892, B1 => n4882, B2 => 
                           n1608, ZN => n8330);
   U2167 : OAI22_X1 port map( A1 => n1740, A2 => n1892, B1 => n4881, B2 => 
                           n1608, ZN => n8329);
   U2168 : OAI22_X1 port map( A1 => n1741, A2 => n1892, B1 => n4880, B2 => 
                           n1608, ZN => n8328);
   U2169 : OAI22_X1 port map( A1 => n1734, A2 => n1892, B1 => n4879, B2 => 
                           n1608, ZN => n8327);
   U2170 : OAI22_X1 port map( A1 => n1735, A2 => n1892, B1 => n4878, B2 => 
                           n1608, ZN => n8326);
   U2171 : OAI22_X1 port map( A1 => n1736, A2 => n1892, B1 => n4877, B2 => 
                           n1608, ZN => n8325);
   U2172 : OAI22_X1 port map( A1 => n1737, A2 => n1892, B1 => n4876, B2 => 
                           n1608, ZN => n8324);
   U2173 : OAI22_X1 port map( A1 => n1730, A2 => n1892, B1 => n4875, B2 => 
                           n1608, ZN => n8323);
   U2174 : OAI22_X1 port map( A1 => n1731, A2 => n1892, B1 => n4874, B2 => 
                           n1608, ZN => n8322);
   U2175 : OAI22_X1 port map( A1 => n1732, A2 => n1892, B1 => n4873, B2 => 
                           n1608, ZN => n8321);
   U2176 : OAI22_X1 port map( A1 => n1733, A2 => n1892, B1 => n4872, B2 => 
                           n1608, ZN => n8320);
   U2177 : OAI22_X1 port map( A1 => n1726, A2 => n1892, B1 => n4871, B2 => 
                           n1608, ZN => n8319);
   U2178 : OAI22_X1 port map( A1 => n1727, A2 => n1892, B1 => n4870, B2 => 
                           n1608, ZN => n8318);
   U2179 : OAI22_X1 port map( A1 => n1728, A2 => n1892, B1 => n4869, B2 => 
                           n1608, ZN => n8317);
   U2180 : OAI22_X1 port map( A1 => n1729, A2 => n1892, B1 => n4868, B2 => 
                           n1608, ZN => n8316);
   U2181 : OAI22_X1 port map( A1 => n1725, A2 => n1892, B1 => n4867, B2 => 
                           n1608, ZN => n8315);
   U2182 : OAI22_X1 port map( A1 => n1768, A2 => n1892, B1 => n4866, B2 => 
                           n1608, ZN => n8314);
   U2183 : OAI21_X1 port map( B1 => n1769, B2 => n1892, A => n1770, ZN => n1893
                           );
   U2184 : OAI22_X1 port map( A1 => n1759, A2 => n1894, B1 => n4865, B2 => 
                           n1602, ZN => n8313);
   U2185 : OAI22_X1 port map( A1 => n1761, A2 => n1894, B1 => n4864, B2 => 
                           n1602, ZN => n8312);
   U2186 : OAI22_X1 port map( A1 => n1762, A2 => n1894, B1 => n4863, B2 => 
                           n1602, ZN => n8311);
   U2187 : OAI22_X1 port map( A1 => n1763, A2 => n1894, B1 => n4862, B2 => 
                           n1602, ZN => n8310);
   U2188 : OAI22_X1 port map( A1 => n1764, A2 => n1894, B1 => n4861, B2 => 
                           n1602, ZN => n8309);
   U2189 : OAI22_X1 port map( A1 => n1765, A2 => n1894, B1 => n4860, B2 => 
                           n1602, ZN => n8308);
   U2190 : OAI22_X1 port map( A1 => n1766, A2 => n1894, B1 => n4859, B2 => 
                           n1602, ZN => n8307);
   U2191 : OAI22_X1 port map( A1 => n1767, A2 => n1894, B1 => n4858, B2 => 
                           n1602, ZN => n8306);
   U2192 : OAI22_X1 port map( A1 => n1746, A2 => n1894, B1 => n4857, B2 => 
                           n1602, ZN => n8305);
   U2193 : OAI22_X1 port map( A1 => n1747, A2 => n1894, B1 => n4856, B2 => 
                           n1602, ZN => n8304);
   U2194 : OAI22_X1 port map( A1 => n1742, A2 => n1894, B1 => n4855, B2 => 
                           n1602, ZN => n8303);
   U2195 : OAI22_X1 port map( A1 => n1743, A2 => n1894, B1 => n4854, B2 => 
                           n1602, ZN => n8302);
   U2196 : OAI22_X1 port map( A1 => n1744, A2 => n1894, B1 => n4853, B2 => 
                           n1602, ZN => n8301);
   U2197 : OAI22_X1 port map( A1 => n1745, A2 => n1894, B1 => n4852, B2 => 
                           n1602, ZN => n8300);
   U2198 : OAI22_X1 port map( A1 => n1738, A2 => n1894, B1 => n4851, B2 => 
                           n1602, ZN => n8299);
   U2199 : OAI22_X1 port map( A1 => n1739, A2 => n1894, B1 => n4850, B2 => 
                           n1602, ZN => n8298);
   U2200 : OAI22_X1 port map( A1 => n1740, A2 => n1894, B1 => n4849, B2 => 
                           n1602, ZN => n8297);
   U2201 : OAI22_X1 port map( A1 => n1741, A2 => n1894, B1 => n4848, B2 => 
                           n1602, ZN => n8296);
   U2202 : OAI22_X1 port map( A1 => n1734, A2 => n1894, B1 => n4847, B2 => 
                           n1602, ZN => n8295);
   U2203 : OAI22_X1 port map( A1 => n1735, A2 => n1894, B1 => n4846, B2 => 
                           n1602, ZN => n8294);
   U2204 : OAI22_X1 port map( A1 => n1736, A2 => n1894, B1 => n4845, B2 => 
                           n1602, ZN => n8293);
   U2205 : OAI22_X1 port map( A1 => n1737, A2 => n1894, B1 => n4844, B2 => 
                           n1602, ZN => n8292);
   U2206 : OAI22_X1 port map( A1 => n1730, A2 => n1894, B1 => n4843, B2 => 
                           n1602, ZN => n8291);
   U2207 : OAI22_X1 port map( A1 => n1731, A2 => n1894, B1 => n4842, B2 => 
                           n1602, ZN => n8290);
   U2208 : OAI22_X1 port map( A1 => n1732, A2 => n1894, B1 => n4841, B2 => 
                           n1602, ZN => n8289);
   U2209 : OAI22_X1 port map( A1 => n1733, A2 => n1894, B1 => n4840, B2 => 
                           n1602, ZN => n8288);
   U2210 : OAI22_X1 port map( A1 => n1726, A2 => n1894, B1 => n4839, B2 => 
                           n1602, ZN => n8287);
   U2211 : OAI22_X1 port map( A1 => n1727, A2 => n1894, B1 => n4838, B2 => 
                           n1602, ZN => n8286);
   U2212 : OAI22_X1 port map( A1 => n1728, A2 => n1894, B1 => n4837, B2 => 
                           n1602, ZN => n8285);
   U2213 : OAI22_X1 port map( A1 => n1729, A2 => n1894, B1 => n4836, B2 => 
                           n1602, ZN => n8284);
   U2214 : OAI22_X1 port map( A1 => n1725, A2 => n1894, B1 => n4835, B2 => 
                           n1602, ZN => n8283);
   U2215 : OAI22_X1 port map( A1 => n1768, A2 => n1894, B1 => n4834, B2 => 
                           n1602, ZN => n8282);
   U2216 : OAI21_X1 port map( B1 => n1769, B2 => n1894, A => n1770, ZN => n1895
                           );
   U2217 : OAI22_X1 port map( A1 => n1759, A2 => n1896, B1 => n4833, B2 => 
                           n1604, ZN => n8281);
   U2218 : OAI22_X1 port map( A1 => n1761, A2 => n1896, B1 => n4832, B2 => 
                           n1604, ZN => n8280);
   U2219 : OAI22_X1 port map( A1 => n1762, A2 => n1896, B1 => n4831, B2 => 
                           n1604, ZN => n8279);
   U2220 : OAI22_X1 port map( A1 => n1763, A2 => n1896, B1 => n4830, B2 => 
                           n1604, ZN => n8278);
   U2221 : OAI22_X1 port map( A1 => n1764, A2 => n1896, B1 => n4829, B2 => 
                           n1604, ZN => n8277);
   U2222 : OAI22_X1 port map( A1 => n1765, A2 => n1896, B1 => n4828, B2 => 
                           n1604, ZN => n8276);
   U2223 : OAI22_X1 port map( A1 => n1766, A2 => n1896, B1 => n4827, B2 => 
                           n1604, ZN => n8275);
   U2224 : OAI22_X1 port map( A1 => n1767, A2 => n1896, B1 => n4826, B2 => 
                           n1604, ZN => n8274);
   U2225 : OAI22_X1 port map( A1 => n1746, A2 => n1896, B1 => n4825, B2 => 
                           n1604, ZN => n8273);
   U2226 : OAI22_X1 port map( A1 => n1747, A2 => n1896, B1 => n4824, B2 => 
                           n1604, ZN => n8272);
   U2227 : OAI22_X1 port map( A1 => n1742, A2 => n1896, B1 => n4823, B2 => 
                           n1604, ZN => n8271);
   U2228 : OAI22_X1 port map( A1 => n1743, A2 => n1896, B1 => n4822, B2 => 
                           n1604, ZN => n8270);
   U2229 : OAI22_X1 port map( A1 => n1744, A2 => n1896, B1 => n4821, B2 => 
                           n1604, ZN => n8269);
   U2230 : OAI22_X1 port map( A1 => n1745, A2 => n1896, B1 => n4820, B2 => 
                           n1604, ZN => n8268);
   U2231 : OAI22_X1 port map( A1 => n1738, A2 => n1896, B1 => n4819, B2 => 
                           n1604, ZN => n8267);
   U2232 : OAI22_X1 port map( A1 => n1739, A2 => n1896, B1 => n4818, B2 => 
                           n1604, ZN => n8266);
   U2233 : OAI22_X1 port map( A1 => n1740, A2 => n1896, B1 => n4817, B2 => 
                           n1604, ZN => n8265);
   U2234 : OAI22_X1 port map( A1 => n1741, A2 => n1896, B1 => n4816, B2 => 
                           n1604, ZN => n8264);
   U2235 : OAI22_X1 port map( A1 => n1734, A2 => n1896, B1 => n4815, B2 => 
                           n1604, ZN => n8263);
   U2236 : OAI22_X1 port map( A1 => n1735, A2 => n1896, B1 => n4814, B2 => 
                           n1604, ZN => n8262);
   U2237 : OAI22_X1 port map( A1 => n1736, A2 => n1896, B1 => n4813, B2 => 
                           n1604, ZN => n8261);
   U2238 : OAI22_X1 port map( A1 => n1737, A2 => n1896, B1 => n4812, B2 => 
                           n1604, ZN => n8260);
   U2239 : OAI22_X1 port map( A1 => n1730, A2 => n1896, B1 => n4811, B2 => 
                           n1604, ZN => n8259);
   U2240 : OAI22_X1 port map( A1 => n1731, A2 => n1896, B1 => n4810, B2 => 
                           n1604, ZN => n8258);
   U2241 : OAI22_X1 port map( A1 => n1732, A2 => n1896, B1 => n4809, B2 => 
                           n1604, ZN => n8257);
   U2242 : OAI22_X1 port map( A1 => n1733, A2 => n1896, B1 => n4808, B2 => 
                           n1604, ZN => n8256);
   U2243 : OAI22_X1 port map( A1 => n1726, A2 => n1896, B1 => n4807, B2 => 
                           n1604, ZN => n8255);
   U2244 : OAI22_X1 port map( A1 => n1727, A2 => n1896, B1 => n4806, B2 => 
                           n1604, ZN => n8254);
   U2245 : OAI22_X1 port map( A1 => n1728, A2 => n1896, B1 => n4805, B2 => 
                           n1604, ZN => n8253);
   U2246 : OAI22_X1 port map( A1 => n1729, A2 => n1896, B1 => n4804, B2 => 
                           n1604, ZN => n8252);
   U2247 : OAI22_X1 port map( A1 => n1725, A2 => n1896, B1 => n4803, B2 => 
                           n1604, ZN => n8251);
   U2248 : OAI22_X1 port map( A1 => n1768, A2 => n1896, B1 => n4802, B2 => 
                           n1604, ZN => n8250);
   U2249 : OAI21_X1 port map( B1 => n1769, B2 => n1896, A => n1770, ZN => n1897
                           );
   U2250 : OAI22_X1 port map( A1 => n1759, A2 => n1898, B1 => n5688, B2 => 
                           n1598, ZN => n8249);
   U2251 : OAI22_X1 port map( A1 => n1761, A2 => n1898, B1 => n5678, B2 => 
                           n1598, ZN => n8248);
   U2252 : OAI22_X1 port map( A1 => n1762, A2 => n1898, B1 => n5668, B2 => 
                           n1598, ZN => n8247);
   U2253 : OAI22_X1 port map( A1 => n1763, A2 => n1898, B1 => n5658, B2 => 
                           n1598, ZN => n8246);
   U2254 : OAI22_X1 port map( A1 => n1764, A2 => n1898, B1 => n5648, B2 => 
                           n1598, ZN => n8245);
   U2255 : OAI22_X1 port map( A1 => n1765, A2 => n1898, B1 => n5638, B2 => 
                           n1598, ZN => n8244);
   U2256 : OAI22_X1 port map( A1 => n1766, A2 => n1898, B1 => n5628, B2 => 
                           n1598, ZN => n8243);
   U2257 : OAI22_X1 port map( A1 => n1767, A2 => n1898, B1 => n5618, B2 => 
                           n1598, ZN => n8242);
   U2258 : OAI22_X1 port map( A1 => n1746, A2 => n1898, B1 => n5608, B2 => 
                           n1598, ZN => n8241);
   U2259 : OAI22_X1 port map( A1 => n1747, A2 => n1898, B1 => n5598, B2 => 
                           n1598, ZN => n8240);
   U2260 : OAI22_X1 port map( A1 => n1742, A2 => n1898, B1 => n5588, B2 => 
                           n1598, ZN => n8239);
   U2261 : OAI22_X1 port map( A1 => n1743, A2 => n1898, B1 => n5578, B2 => 
                           n1598, ZN => n8238);
   U2262 : OAI22_X1 port map( A1 => n1744, A2 => n1898, B1 => n5568, B2 => 
                           n1598, ZN => n8237);
   U2263 : OAI22_X1 port map( A1 => n1745, A2 => n1898, B1 => n5558, B2 => 
                           n1598, ZN => n8236);
   U2264 : OAI22_X1 port map( A1 => n1738, A2 => n1898, B1 => n5548, B2 => 
                           n1598, ZN => n8235);
   U2265 : OAI22_X1 port map( A1 => n1739, A2 => n1898, B1 => n5538, B2 => 
                           n1598, ZN => n8234);
   U2266 : OAI22_X1 port map( A1 => n1740, A2 => n1898, B1 => n5528, B2 => 
                           n1598, ZN => n8233);
   U2267 : OAI22_X1 port map( A1 => n1741, A2 => n1898, B1 => n5518, B2 => 
                           n1598, ZN => n8232);
   U2268 : OAI22_X1 port map( A1 => n1734, A2 => n1898, B1 => n5508, B2 => 
                           n1598, ZN => n8231);
   U2269 : OAI22_X1 port map( A1 => n1735, A2 => n1898, B1 => n5498, B2 => 
                           n1598, ZN => n8230);
   U2270 : OAI22_X1 port map( A1 => n1736, A2 => n1898, B1 => n5488, B2 => 
                           n1598, ZN => n8229);
   U2271 : OAI22_X1 port map( A1 => n1737, A2 => n1898, B1 => n5478, B2 => 
                           n1598, ZN => n8228);
   U2272 : OAI22_X1 port map( A1 => n1730, A2 => n1898, B1 => n5468, B2 => 
                           n1598, ZN => n8227);
   U2273 : OAI22_X1 port map( A1 => n1731, A2 => n1898, B1 => n5458, B2 => 
                           n1598, ZN => n8226);
   U2274 : OAI22_X1 port map( A1 => n1732, A2 => n1898, B1 => n5448, B2 => 
                           n1598, ZN => n8225);
   U2275 : OAI22_X1 port map( A1 => n1733, A2 => n1898, B1 => n5438, B2 => 
                           n1598, ZN => n8224);
   U2276 : OAI22_X1 port map( A1 => n1726, A2 => n1898, B1 => n5428, B2 => 
                           n1598, ZN => n8223);
   U2277 : OAI22_X1 port map( A1 => n1727, A2 => n1898, B1 => n5418, B2 => 
                           n1598, ZN => n8222);
   U2278 : OAI22_X1 port map( A1 => n1728, A2 => n1898, B1 => n5408, B2 => 
                           n1598, ZN => n8221);
   U2279 : OAI22_X1 port map( A1 => n1729, A2 => n1898, B1 => n5398, B2 => 
                           n1598, ZN => n8220);
   U2280 : OAI22_X1 port map( A1 => n1725, A2 => n1898, B1 => n5388, B2 => 
                           n1598, ZN => n8219);
   U2281 : OAI22_X1 port map( A1 => n1768, A2 => n1898, B1 => n5378, B2 => 
                           n1598, ZN => n8218);
   U2282 : OAI21_X1 port map( B1 => n1769, B2 => n1898, A => n1770, ZN => n1899
                           );
   U2283 : OAI22_X1 port map( A1 => n1759, A2 => n1900, B1 => n5689, B2 => 
                           n1600, ZN => n8217);
   U2284 : OAI22_X1 port map( A1 => n1761, A2 => n1900, B1 => n5679, B2 => 
                           n1600, ZN => n8216);
   U2285 : OAI22_X1 port map( A1 => n1762, A2 => n1900, B1 => n5669, B2 => 
                           n1600, ZN => n8215);
   U2286 : OAI22_X1 port map( A1 => n1763, A2 => n1900, B1 => n5659, B2 => 
                           n1600, ZN => n8214);
   U2287 : OAI22_X1 port map( A1 => n1764, A2 => n1900, B1 => n5649, B2 => 
                           n1600, ZN => n8213);
   U2288 : OAI22_X1 port map( A1 => n1765, A2 => n1900, B1 => n5639, B2 => 
                           n1600, ZN => n8212);
   U2289 : OAI22_X1 port map( A1 => n1766, A2 => n1900, B1 => n5629, B2 => 
                           n1600, ZN => n8211);
   U2290 : OAI22_X1 port map( A1 => n1767, A2 => n1900, B1 => n5619, B2 => 
                           n1600, ZN => n8210);
   U2291 : OAI22_X1 port map( A1 => n1746, A2 => n1900, B1 => n5609, B2 => 
                           n1600, ZN => n8209);
   U2292 : OAI22_X1 port map( A1 => n1747, A2 => n1900, B1 => n5599, B2 => 
                           n1600, ZN => n8208);
   U2293 : OAI22_X1 port map( A1 => n1742, A2 => n1900, B1 => n5589, B2 => 
                           n1600, ZN => n8207);
   U2294 : OAI22_X1 port map( A1 => n1743, A2 => n1900, B1 => n5579, B2 => 
                           n1600, ZN => n8206);
   U2295 : OAI22_X1 port map( A1 => n1744, A2 => n1900, B1 => n5569, B2 => 
                           n1600, ZN => n8205);
   U2296 : OAI22_X1 port map( A1 => n1745, A2 => n1900, B1 => n5559, B2 => 
                           n1600, ZN => n8204);
   U2297 : OAI22_X1 port map( A1 => n1738, A2 => n1900, B1 => n5549, B2 => 
                           n1600, ZN => n8203);
   U2298 : OAI22_X1 port map( A1 => n1739, A2 => n1900, B1 => n5539, B2 => 
                           n1600, ZN => n8202);
   U2299 : OAI22_X1 port map( A1 => n1740, A2 => n1900, B1 => n5529, B2 => 
                           n1600, ZN => n8201);
   U2300 : OAI22_X1 port map( A1 => n1741, A2 => n1900, B1 => n5519, B2 => 
                           n1600, ZN => n8200);
   U2301 : OAI22_X1 port map( A1 => n1734, A2 => n1900, B1 => n5509, B2 => 
                           n1600, ZN => n8199);
   U2302 : OAI22_X1 port map( A1 => n1735, A2 => n1900, B1 => n5499, B2 => 
                           n1600, ZN => n8198);
   U2303 : OAI22_X1 port map( A1 => n1736, A2 => n1900, B1 => n5489, B2 => 
                           n1600, ZN => n8197);
   U2304 : OAI22_X1 port map( A1 => n1737, A2 => n1900, B1 => n5479, B2 => 
                           n1600, ZN => n8196);
   U2305 : OAI22_X1 port map( A1 => n1730, A2 => n1900, B1 => n5469, B2 => 
                           n1600, ZN => n8195);
   U2306 : OAI22_X1 port map( A1 => n1731, A2 => n1900, B1 => n5459, B2 => 
                           n1600, ZN => n8194);
   U2307 : OAI22_X1 port map( A1 => n1732, A2 => n1900, B1 => n5449, B2 => 
                           n1600, ZN => n8193);
   U2308 : OAI22_X1 port map( A1 => n1733, A2 => n1900, B1 => n5439, B2 => 
                           n1600, ZN => n8192);
   U2309 : OAI22_X1 port map( A1 => n1726, A2 => n1900, B1 => n5429, B2 => 
                           n1600, ZN => n8191);
   U2310 : OAI22_X1 port map( A1 => n1727, A2 => n1900, B1 => n5419, B2 => 
                           n1600, ZN => n8190);
   U2311 : OAI22_X1 port map( A1 => n1728, A2 => n1900, B1 => n5409, B2 => 
                           n1600, ZN => n8189);
   U2312 : OAI22_X1 port map( A1 => n1729, A2 => n1900, B1 => n5399, B2 => 
                           n1600, ZN => n8188);
   U2313 : OAI22_X1 port map( A1 => n1725, A2 => n1900, B1 => n5389, B2 => 
                           n1600, ZN => n8187);
   U2314 : OAI22_X1 port map( A1 => n1768, A2 => n1900, B1 => n5379, B2 => 
                           n1600, ZN => n8186);
   U2315 : OAI21_X1 port map( B1 => n1769, B2 => n1900, A => n1770, ZN => n1901
                           );
   U2316 : OAI22_X1 port map( A1 => n1759, A2 => n1902, B1 => n1674, B2 => 
                           n1097, ZN => n8185);
   U2317 : OAI22_X1 port map( A1 => n1761, A2 => n1902, B1 => n1674, B2 => 
                           n1098, ZN => n8184);
   U2318 : OAI22_X1 port map( A1 => n1762, A2 => n1902, B1 => n1674, B2 => 
                           n1099, ZN => n8183);
   U2319 : OAI22_X1 port map( A1 => n1763, A2 => n1902, B1 => n1674, B2 => 
                           n1100, ZN => n8182);
   U2320 : OAI22_X1 port map( A1 => n1764, A2 => n1902, B1 => n1674, B2 => 
                           n1101, ZN => n8181);
   U2321 : OAI22_X1 port map( A1 => n1765, A2 => n1902, B1 => n1674, B2 => 
                           n1102, ZN => n8180);
   U2322 : OAI22_X1 port map( A1 => n1766, A2 => n1902, B1 => n1674, B2 => 
                           n1103, ZN => n8179);
   U2323 : OAI22_X1 port map( A1 => n1767, A2 => n1902, B1 => n1674, B2 => 
                           n1104, ZN => n8178);
   U2324 : OAI22_X1 port map( A1 => n1746, A2 => n1902, B1 => n1674, B2 => 
                           n1105, ZN => n8177);
   U2325 : OAI22_X1 port map( A1 => n1747, A2 => n1902, B1 => n1674, B2 => 
                           n1106, ZN => n8176);
   U2326 : OAI22_X1 port map( A1 => n1742, A2 => n1902, B1 => n1674, B2 => 
                           n1107, ZN => n8175);
   U2327 : OAI22_X1 port map( A1 => n1743, A2 => n1902, B1 => n1674, B2 => 
                           n1108, ZN => n8174);
   U2328 : OAI22_X1 port map( A1 => n1744, A2 => n1902, B1 => n1674, B2 => 
                           n1109, ZN => n8173);
   U2329 : OAI22_X1 port map( A1 => n1745, A2 => n1902, B1 => n1674, B2 => 
                           n1110, ZN => n8172);
   U2330 : OAI22_X1 port map( A1 => n1738, A2 => n1902, B1 => n1674, B2 => 
                           n1111, ZN => n8171);
   U2331 : OAI22_X1 port map( A1 => n1739, A2 => n1902, B1 => n1674, B2 => 
                           n1112, ZN => n8170);
   U2332 : OAI22_X1 port map( A1 => n1740, A2 => n1902, B1 => n1674, B2 => 
                           n1113, ZN => n8169);
   U2333 : OAI22_X1 port map( A1 => n1741, A2 => n1902, B1 => n1674, B2 => 
                           n1114, ZN => n8168);
   U2334 : OAI22_X1 port map( A1 => n1734, A2 => n1902, B1 => n1674, B2 => 
                           n1115, ZN => n8167);
   U2335 : OAI22_X1 port map( A1 => n1735, A2 => n1902, B1 => n1674, B2 => 
                           n1116, ZN => n8166);
   U2336 : OAI22_X1 port map( A1 => n1736, A2 => n1902, B1 => n1674, B2 => 
                           n1117, ZN => n8165);
   U2337 : OAI22_X1 port map( A1 => n1737, A2 => n1902, B1 => n1674, B2 => 
                           n1118, ZN => n8164);
   U2338 : OAI22_X1 port map( A1 => n1730, A2 => n1902, B1 => n1674, B2 => 
                           n1119, ZN => n8163);
   U2339 : OAI22_X1 port map( A1 => n1731, A2 => n1902, B1 => n1674, B2 => 
                           n1120, ZN => n8162);
   U2340 : OAI22_X1 port map( A1 => n1732, A2 => n1902, B1 => n1674, B2 => 
                           n1121, ZN => n8161);
   U2341 : OAI22_X1 port map( A1 => n1733, A2 => n1902, B1 => n1674, B2 => 
                           n1122, ZN => n8160);
   U2342 : OAI22_X1 port map( A1 => n1726, A2 => n1902, B1 => n1674, B2 => 
                           n1123, ZN => n8159);
   U2343 : OAI22_X1 port map( A1 => n1727, A2 => n1902, B1 => n1674, B2 => 
                           n1124, ZN => n8158);
   U2344 : OAI22_X1 port map( A1 => n1728, A2 => n1902, B1 => n1674, B2 => 
                           n1125, ZN => n8157);
   U2345 : OAI22_X1 port map( A1 => n1729, A2 => n1902, B1 => n1674, B2 => 
                           n1126, ZN => n8156);
   U2346 : OAI22_X1 port map( A1 => n1725, A2 => n1902, B1 => n1674, B2 => 
                           n1127, ZN => n8155);
   U2347 : OAI22_X1 port map( A1 => n1768, A2 => n1902, B1 => n1674, B2 => 
                           n1128, ZN => n8154);
   U2348 : OAI21_X1 port map( B1 => n1769, B2 => n1902, A => n1770, ZN => n1903
                           );
   U2349 : AND2_X1 port map( A1 => n1904, A2 => n1905, ZN => n1796);
   U2350 : OAI22_X1 port map( A1 => n1759, A2 => n1906, B1 => n1676, B2 => 
                           n1129, ZN => n8153);
   U2351 : OAI22_X1 port map( A1 => n1761, A2 => n1906, B1 => n1676, B2 => 
                           n1130, ZN => n8152);
   U2352 : OAI22_X1 port map( A1 => n1762, A2 => n1906, B1 => n1676, B2 => 
                           n1131, ZN => n8151);
   U2353 : OAI22_X1 port map( A1 => n1763, A2 => n1906, B1 => n1676, B2 => 
                           n1132, ZN => n8150);
   U2354 : OAI22_X1 port map( A1 => n1764, A2 => n1906, B1 => n1676, B2 => 
                           n1133, ZN => n8149);
   U2355 : OAI22_X1 port map( A1 => n1765, A2 => n1906, B1 => n1676, B2 => 
                           n1134, ZN => n8148);
   U2356 : OAI22_X1 port map( A1 => n1766, A2 => n1906, B1 => n1676, B2 => 
                           n1135, ZN => n8147);
   U2357 : OAI22_X1 port map( A1 => n1767, A2 => n1906, B1 => n1676, B2 => 
                           n1136, ZN => n8146);
   U2358 : OAI22_X1 port map( A1 => n1746, A2 => n1906, B1 => n1676, B2 => 
                           n1137, ZN => n8145);
   U2359 : OAI22_X1 port map( A1 => n1747, A2 => n1906, B1 => n1676, B2 => 
                           n1138, ZN => n8144);
   U2360 : OAI22_X1 port map( A1 => n1742, A2 => n1906, B1 => n1676, B2 => 
                           n1139, ZN => n8143);
   U2361 : OAI22_X1 port map( A1 => n1743, A2 => n1906, B1 => n1676, B2 => 
                           n1140, ZN => n8142);
   U2362 : OAI22_X1 port map( A1 => n1744, A2 => n1906, B1 => n1676, B2 => 
                           n1141, ZN => n8141);
   U2363 : OAI22_X1 port map( A1 => n1745, A2 => n1906, B1 => n1676, B2 => 
                           n1142, ZN => n8140);
   U2364 : OAI22_X1 port map( A1 => n1738, A2 => n1906, B1 => n1676, B2 => 
                           n1143, ZN => n8139);
   U2365 : OAI22_X1 port map( A1 => n1739, A2 => n1906, B1 => n1676, B2 => 
                           n1144, ZN => n8138);
   U2366 : OAI22_X1 port map( A1 => n1740, A2 => n1906, B1 => n1676, B2 => 
                           n1145, ZN => n8137);
   U2367 : OAI22_X1 port map( A1 => n1741, A2 => n1906, B1 => n1676, B2 => 
                           n1146, ZN => n8136);
   U2368 : OAI22_X1 port map( A1 => n1734, A2 => n1906, B1 => n1676, B2 => 
                           n1147, ZN => n8135);
   U2369 : OAI22_X1 port map( A1 => n1735, A2 => n1906, B1 => n1676, B2 => 
                           n1148, ZN => n8134);
   U2370 : OAI22_X1 port map( A1 => n1736, A2 => n1906, B1 => n1676, B2 => 
                           n1149, ZN => n8133);
   U2371 : OAI22_X1 port map( A1 => n1737, A2 => n1906, B1 => n1676, B2 => 
                           n1150, ZN => n8132);
   U2372 : OAI22_X1 port map( A1 => n1730, A2 => n1906, B1 => n1676, B2 => 
                           n1151, ZN => n8131);
   U2373 : OAI22_X1 port map( A1 => n1731, A2 => n1906, B1 => n1676, B2 => 
                           n1152, ZN => n8130);
   U2374 : OAI22_X1 port map( A1 => n1732, A2 => n1906, B1 => n1676, B2 => 
                           n1153, ZN => n8129);
   U2375 : OAI22_X1 port map( A1 => n1733, A2 => n1906, B1 => n1676, B2 => 
                           n1154, ZN => n8128);
   U2376 : OAI22_X1 port map( A1 => n1726, A2 => n1906, B1 => n1676, B2 => 
                           n1155, ZN => n8127);
   U2377 : OAI22_X1 port map( A1 => n1727, A2 => n1906, B1 => n1676, B2 => 
                           n1156, ZN => n8126);
   U2378 : OAI22_X1 port map( A1 => n1728, A2 => n1906, B1 => n1676, B2 => 
                           n1157, ZN => n8125);
   U2379 : OAI22_X1 port map( A1 => n1729, A2 => n1906, B1 => n1676, B2 => 
                           n1158, ZN => n8124);
   U2380 : OAI22_X1 port map( A1 => n1725, A2 => n1906, B1 => n1676, B2 => 
                           n1159, ZN => n8123);
   U2381 : OAI22_X1 port map( A1 => n1768, A2 => n1906, B1 => n1676, B2 => 
                           n1160, ZN => n8122);
   U2382 : OAI21_X1 port map( B1 => n1769, B2 => n1906, A => n1770, ZN => n1907
                           );
   U2383 : AND2_X1 port map( A1 => n1904, A2 => n1908, ZN => n1799);
   U2384 : OAI22_X1 port map( A1 => n1759, A2 => n1909, B1 => n1670, B2 => 
                           n1001, ZN => n8121);
   U2385 : OAI22_X1 port map( A1 => n1761, A2 => n1909, B1 => n1670, B2 => 
                           n1002, ZN => n8120);
   U2386 : OAI22_X1 port map( A1 => n1762, A2 => n1909, B1 => n1670, B2 => 
                           n1003, ZN => n8119);
   U2387 : OAI22_X1 port map( A1 => n1763, A2 => n1909, B1 => n1670, B2 => 
                           n1004, ZN => n8118);
   U2388 : OAI22_X1 port map( A1 => n1764, A2 => n1909, B1 => n1670, B2 => 
                           n1005, ZN => n8117);
   U2389 : OAI22_X1 port map( A1 => n1765, A2 => n1909, B1 => n1670, B2 => 
                           n1006, ZN => n8116);
   U2390 : OAI22_X1 port map( A1 => n1766, A2 => n1909, B1 => n1670, B2 => 
                           n1007, ZN => n8115);
   U2391 : OAI22_X1 port map( A1 => n1767, A2 => n1909, B1 => n1670, B2 => 
                           n1008, ZN => n8114);
   U2392 : OAI22_X1 port map( A1 => n1746, A2 => n1909, B1 => n1670, B2 => 
                           n1009, ZN => n8113);
   U2393 : OAI22_X1 port map( A1 => n1747, A2 => n1909, B1 => n1670, B2 => 
                           n1010, ZN => n8112);
   U2394 : OAI22_X1 port map( A1 => n1742, A2 => n1909, B1 => n1670, B2 => 
                           n1011, ZN => n8111);
   U2395 : OAI22_X1 port map( A1 => n1743, A2 => n1909, B1 => n1670, B2 => 
                           n1012, ZN => n8110);
   U2396 : OAI22_X1 port map( A1 => n1744, A2 => n1909, B1 => n1670, B2 => 
                           n1013, ZN => n8109);
   U2397 : OAI22_X1 port map( A1 => n1745, A2 => n1909, B1 => n1670, B2 => 
                           n1014, ZN => n8108);
   U2398 : OAI22_X1 port map( A1 => n1738, A2 => n1909, B1 => n1670, B2 => 
                           n1015, ZN => n8107);
   U2399 : OAI22_X1 port map( A1 => n1739, A2 => n1909, B1 => n1670, B2 => 
                           n1016, ZN => n8106);
   U2400 : OAI22_X1 port map( A1 => n1740, A2 => n1909, B1 => n1670, B2 => 
                           n1017, ZN => n8105);
   U2401 : OAI22_X1 port map( A1 => n1741, A2 => n1909, B1 => n1670, B2 => 
                           n1018, ZN => n8104);
   U2402 : OAI22_X1 port map( A1 => n1734, A2 => n1909, B1 => n1670, B2 => 
                           n1019, ZN => n8103);
   U2403 : OAI22_X1 port map( A1 => n1735, A2 => n1909, B1 => n1670, B2 => 
                           n1020, ZN => n8102);
   U2404 : OAI22_X1 port map( A1 => n1736, A2 => n1909, B1 => n1670, B2 => 
                           n1021, ZN => n8101);
   U2405 : OAI22_X1 port map( A1 => n1737, A2 => n1909, B1 => n1670, B2 => 
                           n1022, ZN => n8100);
   U2406 : OAI22_X1 port map( A1 => n1730, A2 => n1909, B1 => n1670, B2 => 
                           n1023, ZN => n8099);
   U2407 : OAI22_X1 port map( A1 => n1731, A2 => n1909, B1 => n1670, B2 => 
                           n1024, ZN => n8098);
   U2408 : OAI22_X1 port map( A1 => n1732, A2 => n1909, B1 => n1670, B2 => 
                           n1025, ZN => n8097);
   U2409 : OAI22_X1 port map( A1 => n1733, A2 => n1909, B1 => n1670, B2 => 
                           n1026, ZN => n8096);
   U2410 : OAI22_X1 port map( A1 => n1726, A2 => n1909, B1 => n1670, B2 => 
                           n1027, ZN => n8095);
   U2411 : OAI22_X1 port map( A1 => n1727, A2 => n1909, B1 => n1670, B2 => 
                           n1028, ZN => n8094);
   U2412 : OAI22_X1 port map( A1 => n1728, A2 => n1909, B1 => n1670, B2 => 
                           n1029, ZN => n8093);
   U2413 : OAI22_X1 port map( A1 => n1729, A2 => n1909, B1 => n1670, B2 => 
                           n1030, ZN => n8092);
   U2414 : OAI22_X1 port map( A1 => n1725, A2 => n1909, B1 => n1670, B2 => 
                           n1031, ZN => n8091);
   U2415 : OAI22_X1 port map( A1 => n1768, A2 => n1909, B1 => n1670, B2 => 
                           n1032, ZN => n8090);
   U2416 : OAI21_X1 port map( B1 => n1769, B2 => n1909, A => n1770, ZN => n1910
                           );
   U2417 : AND2_X1 port map( A1 => n1904, A2 => n1911, ZN => n1802);
   U2418 : OAI22_X1 port map( A1 => n1759, A2 => n1912, B1 => n1672, B2 => 
                           n1353, ZN => n8089);
   U2419 : OAI22_X1 port map( A1 => n1761, A2 => n1912, B1 => n1672, B2 => 
                           n1354, ZN => n8088);
   U2420 : OAI22_X1 port map( A1 => n1762, A2 => n1912, B1 => n1672, B2 => 
                           n1355, ZN => n8087);
   U2421 : OAI22_X1 port map( A1 => n1763, A2 => n1912, B1 => n1672, B2 => 
                           n1356, ZN => n8086);
   U2422 : OAI22_X1 port map( A1 => n1764, A2 => n1912, B1 => n1672, B2 => 
                           n1357, ZN => n8085);
   U2423 : OAI22_X1 port map( A1 => n1765, A2 => n1912, B1 => n1672, B2 => 
                           n1358, ZN => n8084);
   U2424 : OAI22_X1 port map( A1 => n1766, A2 => n1912, B1 => n1672, B2 => 
                           n1359, ZN => n8083);
   U2425 : OAI22_X1 port map( A1 => n1767, A2 => n1912, B1 => n1672, B2 => 
                           n1360, ZN => n8082);
   U2426 : OAI22_X1 port map( A1 => n1746, A2 => n1912, B1 => n1672, B2 => 
                           n1361, ZN => n8081);
   U2427 : OAI22_X1 port map( A1 => n1747, A2 => n1912, B1 => n1672, B2 => 
                           n1362, ZN => n8080);
   U2428 : OAI22_X1 port map( A1 => n1742, A2 => n1912, B1 => n1672, B2 => 
                           n1363, ZN => n8079);
   U2429 : OAI22_X1 port map( A1 => n1743, A2 => n1912, B1 => n1672, B2 => 
                           n1364, ZN => n8078);
   U2430 : OAI22_X1 port map( A1 => n1744, A2 => n1912, B1 => n1672, B2 => 
                           n1365, ZN => n8077);
   U2431 : OAI22_X1 port map( A1 => n1745, A2 => n1912, B1 => n1672, B2 => 
                           n1366, ZN => n8076);
   U2432 : OAI22_X1 port map( A1 => n1738, A2 => n1912, B1 => n1672, B2 => 
                           n1367, ZN => n8075);
   U2433 : OAI22_X1 port map( A1 => n1739, A2 => n1912, B1 => n1672, B2 => 
                           n1368, ZN => n8074);
   U2434 : OAI22_X1 port map( A1 => n1740, A2 => n1912, B1 => n1672, B2 => 
                           n1369, ZN => n8073);
   U2435 : OAI22_X1 port map( A1 => n1741, A2 => n1912, B1 => n1672, B2 => 
                           n1370, ZN => n8072);
   U2436 : OAI22_X1 port map( A1 => n1734, A2 => n1912, B1 => n1672, B2 => 
                           n1371, ZN => n8071);
   U2437 : OAI22_X1 port map( A1 => n1735, A2 => n1912, B1 => n1672, B2 => 
                           n1372, ZN => n8070);
   U2438 : OAI22_X1 port map( A1 => n1736, A2 => n1912, B1 => n1672, B2 => 
                           n1373, ZN => n8069);
   U2439 : OAI22_X1 port map( A1 => n1737, A2 => n1912, B1 => n1672, B2 => 
                           n1374, ZN => n8068);
   U2440 : OAI22_X1 port map( A1 => n1730, A2 => n1912, B1 => n1672, B2 => 
                           n1375, ZN => n8067);
   U2441 : OAI22_X1 port map( A1 => n1731, A2 => n1912, B1 => n1672, B2 => 
                           n1376, ZN => n8066);
   U2442 : OAI22_X1 port map( A1 => n1732, A2 => n1912, B1 => n1672, B2 => 
                           n1377, ZN => n8065);
   U2443 : OAI22_X1 port map( A1 => n1733, A2 => n1912, B1 => n1672, B2 => 
                           n1378, ZN => n8064);
   U2444 : OAI22_X1 port map( A1 => n1726, A2 => n1912, B1 => n1672, B2 => 
                           n1379, ZN => n8063);
   U2445 : OAI22_X1 port map( A1 => n1727, A2 => n1912, B1 => n1672, B2 => 
                           n1380, ZN => n8062);
   U2446 : OAI22_X1 port map( A1 => n1728, A2 => n1912, B1 => n1672, B2 => 
                           n1381, ZN => n8061);
   U2447 : OAI22_X1 port map( A1 => n1729, A2 => n1912, B1 => n1672, B2 => 
                           n1382, ZN => n8060);
   U2448 : OAI22_X1 port map( A1 => n1725, A2 => n1912, B1 => n1672, B2 => 
                           n1383, ZN => n8059);
   U2449 : OAI22_X1 port map( A1 => n1768, A2 => n1912, B1 => n1672, B2 => 
                           n1384, ZN => n8058);
   U2450 : OAI21_X1 port map( B1 => n1769, B2 => n1912, A => n1770, ZN => n1913
                           );
   U2451 : AND2_X1 port map( A1 => n1904, A2 => n1914, ZN => n1805);
   U2452 : AND2_X1 port map( A1 => ADD_WR(3), A2 => n1915, ZN => n1904);
   U2453 : OAI22_X1 port map( A1 => n1759, A2 => n1916, B1 => n4801, B2 => 
                           n1594, ZN => n8057);
   U2454 : OAI22_X1 port map( A1 => n1761, A2 => n1916, B1 => n4800, B2 => 
                           n1594, ZN => n8056);
   U2455 : OAI22_X1 port map( A1 => n1762, A2 => n1916, B1 => n4799, B2 => 
                           n1594, ZN => n8055);
   U2456 : OAI22_X1 port map( A1 => n1763, A2 => n1916, B1 => n4798, B2 => 
                           n1594, ZN => n8054);
   U2457 : OAI22_X1 port map( A1 => n1764, A2 => n1916, B1 => n4797, B2 => 
                           n1594, ZN => n8053);
   U2458 : OAI22_X1 port map( A1 => n1765, A2 => n1916, B1 => n4796, B2 => 
                           n1594, ZN => n8052);
   U2459 : OAI22_X1 port map( A1 => n1766, A2 => n1916, B1 => n4795, B2 => 
                           n1594, ZN => n8051);
   U2460 : OAI22_X1 port map( A1 => n1767, A2 => n1916, B1 => n4794, B2 => 
                           n1594, ZN => n8050);
   U2461 : OAI22_X1 port map( A1 => n1746, A2 => n1916, B1 => n4793, B2 => 
                           n1594, ZN => n8049);
   U2462 : OAI22_X1 port map( A1 => n1747, A2 => n1916, B1 => n4792, B2 => 
                           n1594, ZN => n8048);
   U2463 : OAI22_X1 port map( A1 => n1742, A2 => n1916, B1 => n4791, B2 => 
                           n1594, ZN => n8047);
   U2464 : OAI22_X1 port map( A1 => n1743, A2 => n1916, B1 => n4790, B2 => 
                           n1594, ZN => n8046);
   U2465 : OAI22_X1 port map( A1 => n1744, A2 => n1916, B1 => n4789, B2 => 
                           n1594, ZN => n8045);
   U2466 : OAI22_X1 port map( A1 => n1745, A2 => n1916, B1 => n4788, B2 => 
                           n1594, ZN => n8044);
   U2467 : OAI22_X1 port map( A1 => n1738, A2 => n1916, B1 => n4787, B2 => 
                           n1594, ZN => n8043);
   U2468 : OAI22_X1 port map( A1 => n1739, A2 => n1916, B1 => n4786, B2 => 
                           n1594, ZN => n8042);
   U2469 : OAI22_X1 port map( A1 => n1740, A2 => n1916, B1 => n4785, B2 => 
                           n1594, ZN => n8041);
   U2470 : OAI22_X1 port map( A1 => n1741, A2 => n1916, B1 => n4784, B2 => 
                           n1594, ZN => n8040);
   U2471 : OAI22_X1 port map( A1 => n1734, A2 => n1916, B1 => n4783, B2 => 
                           n1594, ZN => n8039);
   U2472 : OAI22_X1 port map( A1 => n1735, A2 => n1916, B1 => n4782, B2 => 
                           n1594, ZN => n8038);
   U2473 : OAI22_X1 port map( A1 => n1736, A2 => n1916, B1 => n4781, B2 => 
                           n1594, ZN => n8037);
   U2474 : OAI22_X1 port map( A1 => n1737, A2 => n1916, B1 => n4780, B2 => 
                           n1594, ZN => n8036);
   U2475 : OAI22_X1 port map( A1 => n1730, A2 => n1916, B1 => n4779, B2 => 
                           n1594, ZN => n8035);
   U2476 : OAI22_X1 port map( A1 => n1731, A2 => n1916, B1 => n4778, B2 => 
                           n1594, ZN => n8034);
   U2477 : OAI22_X1 port map( A1 => n1732, A2 => n1916, B1 => n4777, B2 => 
                           n1594, ZN => n8033);
   U2478 : OAI22_X1 port map( A1 => n1733, A2 => n1916, B1 => n4776, B2 => 
                           n1594, ZN => n8032);
   U2479 : OAI22_X1 port map( A1 => n1726, A2 => n1916, B1 => n4775, B2 => 
                           n1594, ZN => n8031);
   U2480 : OAI22_X1 port map( A1 => n1727, A2 => n1916, B1 => n4774, B2 => 
                           n1594, ZN => n8030);
   U2481 : OAI22_X1 port map( A1 => n1728, A2 => n1916, B1 => n4773, B2 => 
                           n1594, ZN => n8029);
   U2482 : OAI22_X1 port map( A1 => n1729, A2 => n1916, B1 => n4772, B2 => 
                           n1594, ZN => n8028);
   U2483 : OAI22_X1 port map( A1 => n1725, A2 => n1916, B1 => n4771, B2 => 
                           n1594, ZN => n8027);
   U2484 : OAI22_X1 port map( A1 => n1768, A2 => n1916, B1 => n4770, B2 => 
                           n1594, ZN => n8026);
   U2485 : OAI21_X1 port map( B1 => n1769, B2 => n1916, A => n1770, ZN => n1917
                           );
   U2486 : AND2_X1 port map( A1 => n1918, A2 => n1905, ZN => n1808);
   U2487 : OAI22_X1 port map( A1 => n1759, A2 => n1919, B1 => n4769, B2 => 
                           n1596, ZN => n8025);
   U2488 : OAI22_X1 port map( A1 => n1761, A2 => n1919, B1 => n4768, B2 => 
                           n1596, ZN => n8024);
   U2489 : OAI22_X1 port map( A1 => n1762, A2 => n1919, B1 => n4767, B2 => 
                           n1596, ZN => n8023);
   U2490 : OAI22_X1 port map( A1 => n1763, A2 => n1919, B1 => n4766, B2 => 
                           n1596, ZN => n8022);
   U2491 : OAI22_X1 port map( A1 => n1764, A2 => n1919, B1 => n4765, B2 => 
                           n1596, ZN => n8021);
   U2492 : OAI22_X1 port map( A1 => n1765, A2 => n1919, B1 => n4764, B2 => 
                           n1596, ZN => n8020);
   U2493 : OAI22_X1 port map( A1 => n1766, A2 => n1919, B1 => n4763, B2 => 
                           n1596, ZN => n8019);
   U2494 : OAI22_X1 port map( A1 => n1767, A2 => n1919, B1 => n4762, B2 => 
                           n1596, ZN => n8018);
   U2495 : OAI22_X1 port map( A1 => n1746, A2 => n1919, B1 => n4761, B2 => 
                           n1596, ZN => n8017);
   U2496 : OAI22_X1 port map( A1 => n1747, A2 => n1919, B1 => n4760, B2 => 
                           n1596, ZN => n8016);
   U2497 : OAI22_X1 port map( A1 => n1742, A2 => n1919, B1 => n4759, B2 => 
                           n1596, ZN => n8015);
   U2498 : OAI22_X1 port map( A1 => n1743, A2 => n1919, B1 => n4758, B2 => 
                           n1596, ZN => n8014);
   U2499 : OAI22_X1 port map( A1 => n1744, A2 => n1919, B1 => n4757, B2 => 
                           n1596, ZN => n8013);
   U2500 : OAI22_X1 port map( A1 => n1745, A2 => n1919, B1 => n4756, B2 => 
                           n1596, ZN => n8012);
   U2501 : OAI22_X1 port map( A1 => n1738, A2 => n1919, B1 => n4755, B2 => 
                           n1596, ZN => n8011);
   U2502 : OAI22_X1 port map( A1 => n1739, A2 => n1919, B1 => n4754, B2 => 
                           n1596, ZN => n8010);
   U2503 : OAI22_X1 port map( A1 => n1740, A2 => n1919, B1 => n4753, B2 => 
                           n1596, ZN => n8009);
   U2504 : OAI22_X1 port map( A1 => n1741, A2 => n1919, B1 => n4752, B2 => 
                           n1596, ZN => n8008);
   U2505 : OAI22_X1 port map( A1 => n1734, A2 => n1919, B1 => n4751, B2 => 
                           n1596, ZN => n8007);
   U2506 : OAI22_X1 port map( A1 => n1735, A2 => n1919, B1 => n4750, B2 => 
                           n1596, ZN => n8006);
   U2507 : OAI22_X1 port map( A1 => n1736, A2 => n1919, B1 => n4749, B2 => 
                           n1596, ZN => n8005);
   U2508 : OAI22_X1 port map( A1 => n1737, A2 => n1919, B1 => n4748, B2 => 
                           n1596, ZN => n8004);
   U2509 : OAI22_X1 port map( A1 => n1730, A2 => n1919, B1 => n4747, B2 => 
                           n1596, ZN => n8003);
   U2510 : OAI22_X1 port map( A1 => n1731, A2 => n1919, B1 => n4746, B2 => 
                           n1596, ZN => n8002);
   U2511 : OAI22_X1 port map( A1 => n1732, A2 => n1919, B1 => n4745, B2 => 
                           n1596, ZN => n8001);
   U2512 : OAI22_X1 port map( A1 => n1733, A2 => n1919, B1 => n4744, B2 => 
                           n1596, ZN => n8000);
   U2513 : OAI22_X1 port map( A1 => n1726, A2 => n1919, B1 => n4743, B2 => 
                           n1596, ZN => n7999);
   U2514 : OAI22_X1 port map( A1 => n1727, A2 => n1919, B1 => n4742, B2 => 
                           n1596, ZN => n7998);
   U2515 : OAI22_X1 port map( A1 => n1728, A2 => n1919, B1 => n4741, B2 => 
                           n1596, ZN => n7997);
   U2516 : OAI22_X1 port map( A1 => n1729, A2 => n1919, B1 => n4740, B2 => 
                           n1596, ZN => n7996);
   U2517 : OAI22_X1 port map( A1 => n1725, A2 => n1919, B1 => n4739, B2 => 
                           n1596, ZN => n7995);
   U2518 : OAI22_X1 port map( A1 => n1768, A2 => n1919, B1 => n4738, B2 => 
                           n1596, ZN => n7994);
   U2519 : OAI21_X1 port map( B1 => n1769, B2 => n1919, A => n1770, ZN => n1920
                           );
   U2520 : AND2_X1 port map( A1 => n1918, A2 => n1908, ZN => n1811);
   U2521 : OAI22_X1 port map( A1 => n1759, A2 => n1921, B1 => n4737, B2 => 
                           n1590, ZN => n7993);
   U2522 : OAI22_X1 port map( A1 => n1761, A2 => n1921, B1 => n4736, B2 => 
                           n1590, ZN => n7992);
   U2523 : OAI22_X1 port map( A1 => n1762, A2 => n1921, B1 => n4735, B2 => 
                           n1590, ZN => n7991);
   U2524 : OAI22_X1 port map( A1 => n1763, A2 => n1921, B1 => n4734, B2 => 
                           n1590, ZN => n7990);
   U2525 : OAI22_X1 port map( A1 => n1764, A2 => n1921, B1 => n4733, B2 => 
                           n1590, ZN => n7989);
   U2526 : OAI22_X1 port map( A1 => n1765, A2 => n1921, B1 => n4732, B2 => 
                           n1590, ZN => n7988);
   U2527 : OAI22_X1 port map( A1 => n1766, A2 => n1921, B1 => n4731, B2 => 
                           n1590, ZN => n7987);
   U2528 : OAI22_X1 port map( A1 => n1767, A2 => n1921, B1 => n4730, B2 => 
                           n1590, ZN => n7986);
   U2529 : OAI22_X1 port map( A1 => n1746, A2 => n1921, B1 => n4729, B2 => 
                           n1590, ZN => n7985);
   U2530 : OAI22_X1 port map( A1 => n1747, A2 => n1921, B1 => n4728, B2 => 
                           n1590, ZN => n7984);
   U2531 : OAI22_X1 port map( A1 => n1742, A2 => n1921, B1 => n4727, B2 => 
                           n1590, ZN => n7983);
   U2532 : OAI22_X1 port map( A1 => n1743, A2 => n1921, B1 => n4726, B2 => 
                           n1590, ZN => n7982);
   U2533 : OAI22_X1 port map( A1 => n1744, A2 => n1921, B1 => n4725, B2 => 
                           n1590, ZN => n7981);
   U2534 : OAI22_X1 port map( A1 => n1745, A2 => n1921, B1 => n4724, B2 => 
                           n1590, ZN => n7980);
   U2535 : OAI22_X1 port map( A1 => n1738, A2 => n1921, B1 => n4723, B2 => 
                           n1590, ZN => n7979);
   U2536 : OAI22_X1 port map( A1 => n1739, A2 => n1921, B1 => n4722, B2 => 
                           n1590, ZN => n7978);
   U2537 : OAI22_X1 port map( A1 => n1740, A2 => n1921, B1 => n4721, B2 => 
                           n1590, ZN => n7977);
   U2538 : OAI22_X1 port map( A1 => n1741, A2 => n1921, B1 => n4720, B2 => 
                           n1590, ZN => n7976);
   U2539 : OAI22_X1 port map( A1 => n1734, A2 => n1921, B1 => n4719, B2 => 
                           n1590, ZN => n7975);
   U2540 : OAI22_X1 port map( A1 => n1735, A2 => n1921, B1 => n4718, B2 => 
                           n1590, ZN => n7974);
   U2541 : OAI22_X1 port map( A1 => n1736, A2 => n1921, B1 => n4717, B2 => 
                           n1590, ZN => n7973);
   U2542 : OAI22_X1 port map( A1 => n1737, A2 => n1921, B1 => n4716, B2 => 
                           n1590, ZN => n7972);
   U2543 : OAI22_X1 port map( A1 => n1730, A2 => n1921, B1 => n4715, B2 => 
                           n1590, ZN => n7971);
   U2544 : OAI22_X1 port map( A1 => n1731, A2 => n1921, B1 => n4714, B2 => 
                           n1590, ZN => n7970);
   U2545 : OAI22_X1 port map( A1 => n1732, A2 => n1921, B1 => n4713, B2 => 
                           n1590, ZN => n7969);
   U2546 : OAI22_X1 port map( A1 => n1733, A2 => n1921, B1 => n4712, B2 => 
                           n1590, ZN => n7968);
   U2547 : OAI22_X1 port map( A1 => n1726, A2 => n1921, B1 => n4711, B2 => 
                           n1590, ZN => n7967);
   U2548 : OAI22_X1 port map( A1 => n1727, A2 => n1921, B1 => n4710, B2 => 
                           n1590, ZN => n7966);
   U2549 : OAI22_X1 port map( A1 => n1728, A2 => n1921, B1 => n4709, B2 => 
                           n1590, ZN => n7965);
   U2550 : OAI22_X1 port map( A1 => n1729, A2 => n1921, B1 => n4708, B2 => 
                           n1590, ZN => n7964);
   U2551 : OAI22_X1 port map( A1 => n1725, A2 => n1921, B1 => n4707, B2 => 
                           n1590, ZN => n7963);
   U2552 : OAI22_X1 port map( A1 => n1768, A2 => n1921, B1 => n4706, B2 => 
                           n1590, ZN => n7962);
   U2553 : OAI21_X1 port map( B1 => n1769, B2 => n1921, A => n1770, ZN => n1922
                           );
   U2554 : AND2_X1 port map( A1 => n1918, A2 => n1911, ZN => n1814);
   U2555 : OAI22_X1 port map( A1 => n1759, A2 => n1923, B1 => n1666, B2 => 
                           n1033, ZN => n7961);
   U2556 : OAI22_X1 port map( A1 => n1761, A2 => n1923, B1 => n1666, B2 => 
                           n1034, ZN => n7960);
   U2557 : OAI22_X1 port map( A1 => n1762, A2 => n1923, B1 => n1666, B2 => 
                           n1035, ZN => n7959);
   U2558 : OAI22_X1 port map( A1 => n1763, A2 => n1923, B1 => n1666, B2 => 
                           n1036, ZN => n7958);
   U2559 : OAI22_X1 port map( A1 => n1764, A2 => n1923, B1 => n1666, B2 => 
                           n1037, ZN => n7957);
   U2560 : OAI22_X1 port map( A1 => n1765, A2 => n1923, B1 => n1666, B2 => 
                           n1038, ZN => n7956);
   U2561 : OAI22_X1 port map( A1 => n1766, A2 => n1923, B1 => n1666, B2 => 
                           n1039, ZN => n7955);
   U2562 : OAI22_X1 port map( A1 => n1767, A2 => n1923, B1 => n1666, B2 => 
                           n1040, ZN => n7954);
   U2563 : OAI22_X1 port map( A1 => n1746, A2 => n1923, B1 => n1666, B2 => 
                           n1041, ZN => n7953);
   U2564 : OAI22_X1 port map( A1 => n1747, A2 => n1923, B1 => n1666, B2 => 
                           n1042, ZN => n7952);
   U2565 : OAI22_X1 port map( A1 => n1742, A2 => n1923, B1 => n1666, B2 => 
                           n1043, ZN => n7951);
   U2566 : OAI22_X1 port map( A1 => n1743, A2 => n1923, B1 => n1666, B2 => 
                           n1044, ZN => n7950);
   U2567 : OAI22_X1 port map( A1 => n1744, A2 => n1923, B1 => n1666, B2 => 
                           n1045, ZN => n7949);
   U2568 : OAI22_X1 port map( A1 => n1745, A2 => n1923, B1 => n1666, B2 => 
                           n1046, ZN => n7948);
   U2569 : OAI22_X1 port map( A1 => n1738, A2 => n1923, B1 => n1666, B2 => 
                           n1047, ZN => n7947);
   U2570 : OAI22_X1 port map( A1 => n1739, A2 => n1923, B1 => n1666, B2 => 
                           n1048, ZN => n7946);
   U2571 : OAI22_X1 port map( A1 => n1740, A2 => n1923, B1 => n1666, B2 => 
                           n1049, ZN => n7945);
   U2572 : OAI22_X1 port map( A1 => n1741, A2 => n1923, B1 => n1666, B2 => 
                           n1050, ZN => n7944);
   U2573 : OAI22_X1 port map( A1 => n1734, A2 => n1923, B1 => n1666, B2 => 
                           n1051, ZN => n7943);
   U2574 : OAI22_X1 port map( A1 => n1735, A2 => n1923, B1 => n1666, B2 => 
                           n1052, ZN => n7942);
   U2575 : OAI22_X1 port map( A1 => n1736, A2 => n1923, B1 => n1666, B2 => 
                           n1053, ZN => n7941);
   U2576 : OAI22_X1 port map( A1 => n1737, A2 => n1923, B1 => n1666, B2 => 
                           n1054, ZN => n7940);
   U2577 : OAI22_X1 port map( A1 => n1730, A2 => n1923, B1 => n1666, B2 => 
                           n1055, ZN => n7939);
   U2578 : OAI22_X1 port map( A1 => n1731, A2 => n1923, B1 => n1666, B2 => 
                           n1056, ZN => n7938);
   U2579 : OAI22_X1 port map( A1 => n1732, A2 => n1923, B1 => n1666, B2 => 
                           n1057, ZN => n7937);
   U2580 : OAI22_X1 port map( A1 => n1733, A2 => n1923, B1 => n1666, B2 => 
                           n1058, ZN => n7936);
   U2581 : OAI22_X1 port map( A1 => n1726, A2 => n1923, B1 => n1666, B2 => 
                           n1059, ZN => n7935);
   U2582 : OAI22_X1 port map( A1 => n1727, A2 => n1923, B1 => n1666, B2 => 
                           n1060, ZN => n7934);
   U2583 : OAI22_X1 port map( A1 => n1728, A2 => n1923, B1 => n1666, B2 => 
                           n1061, ZN => n7933);
   U2584 : OAI22_X1 port map( A1 => n1729, A2 => n1923, B1 => n1666, B2 => 
                           n1062, ZN => n7932);
   U2585 : OAI22_X1 port map( A1 => n1725, A2 => n1923, B1 => n1666, B2 => 
                           n1063, ZN => n7931);
   U2586 : OAI22_X1 port map( A1 => n1768, A2 => n1923, B1 => n1666, B2 => 
                           n1064, ZN => n7930);
   U2587 : OAI21_X1 port map( B1 => n1769, B2 => n1923, A => n1770, ZN => n1924
                           );
   U2588 : AND2_X1 port map( A1 => n1918, A2 => n1914, ZN => n1816);
   U2589 : AND2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n1918);
   U2590 : OAI22_X1 port map( A1 => n1759, A2 => n1925, B1 => n1668, B2 => 
                           n1385, ZN => n7929);
   U2591 : OAI22_X1 port map( A1 => n1761, A2 => n1925, B1 => n1668, B2 => 
                           n1386, ZN => n7928);
   U2592 : OAI22_X1 port map( A1 => n1762, A2 => n1925, B1 => n1668, B2 => 
                           n1387, ZN => n7927);
   U2593 : OAI22_X1 port map( A1 => n1763, A2 => n1925, B1 => n1668, B2 => 
                           n1388, ZN => n7926);
   U2594 : OAI22_X1 port map( A1 => n1764, A2 => n1925, B1 => n1668, B2 => 
                           n1389, ZN => n7925);
   U2595 : OAI22_X1 port map( A1 => n1765, A2 => n1925, B1 => n1668, B2 => 
                           n1390, ZN => n7924);
   U2596 : OAI22_X1 port map( A1 => n1766, A2 => n1925, B1 => n1668, B2 => 
                           n1391, ZN => n7923);
   U2597 : OAI22_X1 port map( A1 => n1767, A2 => n1925, B1 => n1668, B2 => 
                           n1392, ZN => n7922);
   U2598 : OAI22_X1 port map( A1 => n1746, A2 => n1925, B1 => n1668, B2 => 
                           n1393, ZN => n7921);
   U2599 : OAI22_X1 port map( A1 => n1747, A2 => n1925, B1 => n1668, B2 => 
                           n1394, ZN => n7920);
   U2600 : OAI22_X1 port map( A1 => n1742, A2 => n1925, B1 => n1668, B2 => 
                           n1395, ZN => n7919);
   U2601 : OAI22_X1 port map( A1 => n1743, A2 => n1925, B1 => n1668, B2 => 
                           n1396, ZN => n7918);
   U2602 : OAI22_X1 port map( A1 => n1744, A2 => n1925, B1 => n1668, B2 => 
                           n1397, ZN => n7917);
   U2603 : OAI22_X1 port map( A1 => n1745, A2 => n1925, B1 => n1668, B2 => 
                           n1398, ZN => n7916);
   U2604 : OAI22_X1 port map( A1 => n1738, A2 => n1925, B1 => n1668, B2 => 
                           n1399, ZN => n7915);
   U2605 : OAI22_X1 port map( A1 => n1739, A2 => n1925, B1 => n1668, B2 => 
                           n1400, ZN => n7914);
   U2606 : OAI22_X1 port map( A1 => n1740, A2 => n1925, B1 => n1668, B2 => 
                           n1401, ZN => n7913);
   U2607 : OAI22_X1 port map( A1 => n1741, A2 => n1925, B1 => n1668, B2 => 
                           n1402, ZN => n7912);
   U2608 : OAI22_X1 port map( A1 => n1734, A2 => n1925, B1 => n1668, B2 => 
                           n1403, ZN => n7911);
   U2609 : OAI22_X1 port map( A1 => n1735, A2 => n1925, B1 => n1668, B2 => 
                           n1404, ZN => n7910);
   U2610 : OAI22_X1 port map( A1 => n1736, A2 => n1925, B1 => n1668, B2 => 
                           n1405, ZN => n7909);
   U2611 : OAI22_X1 port map( A1 => n1737, A2 => n1925, B1 => n1668, B2 => 
                           n1406, ZN => n7908);
   U2612 : OAI22_X1 port map( A1 => n1730, A2 => n1925, B1 => n1668, B2 => 
                           n1407, ZN => n7907);
   U2613 : OAI22_X1 port map( A1 => n1731, A2 => n1925, B1 => n1668, B2 => 
                           n1408, ZN => n7906);
   U2614 : OAI22_X1 port map( A1 => n1732, A2 => n1925, B1 => n1668, B2 => 
                           n1409, ZN => n7905);
   U2615 : OAI22_X1 port map( A1 => n1733, A2 => n1925, B1 => n1668, B2 => 
                           n1410, ZN => n7904);
   U2616 : OAI22_X1 port map( A1 => n1726, A2 => n1925, B1 => n1668, B2 => 
                           n1411, ZN => n7903);
   U2617 : OAI22_X1 port map( A1 => n1727, A2 => n1925, B1 => n1668, B2 => 
                           n1412, ZN => n7902);
   U2618 : OAI22_X1 port map( A1 => n1728, A2 => n1925, B1 => n1668, B2 => 
                           n1413, ZN => n7901);
   U2619 : OAI22_X1 port map( A1 => n1729, A2 => n1925, B1 => n1668, B2 => 
                           n1414, ZN => n7900);
   U2620 : OAI22_X1 port map( A1 => n1725, A2 => n1925, B1 => n1668, B2 => 
                           n1415, ZN => n7899);
   U2621 : OAI22_X1 port map( A1 => n1768, A2 => n1925, B1 => n1668, B2 => 
                           n1416, ZN => n7898);
   U2622 : OAI21_X1 port map( B1 => n1769, B2 => n1925, A => n1770, ZN => n1926
                           );
   U2623 : AND2_X1 port map( A1 => n1928, A2 => n1905, ZN => n1771);
   U2624 : OAI22_X1 port map( A1 => n1759, A2 => n1929, B1 => n4705, B2 => 
                           n1592, ZN => n7897);
   U2625 : OAI22_X1 port map( A1 => n1761, A2 => n1929, B1 => n4704, B2 => 
                           n1592, ZN => n7896);
   U2626 : OAI22_X1 port map( A1 => n1762, A2 => n1929, B1 => n4703, B2 => 
                           n1592, ZN => n7895);
   U2627 : OAI22_X1 port map( A1 => n1763, A2 => n1929, B1 => n4702, B2 => 
                           n1592, ZN => n7894);
   U2628 : OAI22_X1 port map( A1 => n1764, A2 => n1929, B1 => n4701, B2 => 
                           n1592, ZN => n7893);
   U2629 : OAI22_X1 port map( A1 => n1765, A2 => n1929, B1 => n4700, B2 => 
                           n1592, ZN => n7892);
   U2630 : OAI22_X1 port map( A1 => n1766, A2 => n1929, B1 => n4699, B2 => 
                           n1592, ZN => n7891);
   U2631 : OAI22_X1 port map( A1 => n1767, A2 => n1929, B1 => n4698, B2 => 
                           n1592, ZN => n7890);
   U2632 : OAI22_X1 port map( A1 => n1746, A2 => n1929, B1 => n4697, B2 => 
                           n1592, ZN => n7889);
   U2633 : OAI22_X1 port map( A1 => n1747, A2 => n1929, B1 => n4696, B2 => 
                           n1592, ZN => n7888);
   U2634 : OAI22_X1 port map( A1 => n1742, A2 => n1929, B1 => n4695, B2 => 
                           n1592, ZN => n7887);
   U2635 : OAI22_X1 port map( A1 => n1743, A2 => n1929, B1 => n4694, B2 => 
                           n1592, ZN => n7886);
   U2636 : OAI22_X1 port map( A1 => n1744, A2 => n1929, B1 => n4693, B2 => 
                           n1592, ZN => n7885);
   U2637 : OAI22_X1 port map( A1 => n1745, A2 => n1929, B1 => n4692, B2 => 
                           n1592, ZN => n7884);
   U2638 : OAI22_X1 port map( A1 => n1738, A2 => n1929, B1 => n4691, B2 => 
                           n1592, ZN => n7883);
   U2639 : OAI22_X1 port map( A1 => n1739, A2 => n1929, B1 => n4690, B2 => 
                           n1592, ZN => n7882);
   U2640 : OAI22_X1 port map( A1 => n1740, A2 => n1929, B1 => n4689, B2 => 
                           n1592, ZN => n7881);
   U2641 : OAI22_X1 port map( A1 => n1741, A2 => n1929, B1 => n4688, B2 => 
                           n1592, ZN => n7880);
   U2642 : OAI22_X1 port map( A1 => n1734, A2 => n1929, B1 => n4687, B2 => 
                           n1592, ZN => n7879);
   U2643 : OAI22_X1 port map( A1 => n1735, A2 => n1929, B1 => n4686, B2 => 
                           n1592, ZN => n7878);
   U2644 : OAI22_X1 port map( A1 => n1736, A2 => n1929, B1 => n4685, B2 => 
                           n1592, ZN => n7877);
   U2645 : OAI22_X1 port map( A1 => n1737, A2 => n1929, B1 => n4684, B2 => 
                           n1592, ZN => n7876);
   U2646 : OAI22_X1 port map( A1 => n1730, A2 => n1929, B1 => n4683, B2 => 
                           n1592, ZN => n7875);
   U2647 : OAI22_X1 port map( A1 => n1731, A2 => n1929, B1 => n4682, B2 => 
                           n1592, ZN => n7874);
   U2648 : OAI22_X1 port map( A1 => n1732, A2 => n1929, B1 => n4681, B2 => 
                           n1592, ZN => n7873);
   U2649 : OAI22_X1 port map( A1 => n1733, A2 => n1929, B1 => n4680, B2 => 
                           n1592, ZN => n7872);
   U2650 : OAI22_X1 port map( A1 => n1726, A2 => n1929, B1 => n4679, B2 => 
                           n1592, ZN => n7871);
   U2651 : OAI22_X1 port map( A1 => n1727, A2 => n1929, B1 => n4678, B2 => 
                           n1592, ZN => n7870);
   U2652 : OAI22_X1 port map( A1 => n1728, A2 => n1929, B1 => n4677, B2 => 
                           n1592, ZN => n7869);
   U2653 : OAI22_X1 port map( A1 => n1729, A2 => n1929, B1 => n4676, B2 => 
                           n1592, ZN => n7868);
   U2654 : OAI22_X1 port map( A1 => n1725, A2 => n1929, B1 => n4675, B2 => 
                           n1592, ZN => n7867);
   U2655 : OAI22_X1 port map( A1 => n1768, A2 => n1929, B1 => n4674, B2 => 
                           n1592, ZN => n7866);
   U2656 : OAI21_X1 port map( B1 => n1769, B2 => n1929, A => n1770, ZN => n1930
                           );
   U2657 : AND2_X1 port map( A1 => n1908, A2 => n1928, ZN => n1775);
   U2658 : OAI22_X1 port map( A1 => n1759, A2 => n1931, B1 => n4673, B2 => 
                           n1586, ZN => n7865);
   U2659 : OAI22_X1 port map( A1 => n1761, A2 => n1931, B1 => n4672, B2 => 
                           n1586, ZN => n7864);
   U2660 : OAI22_X1 port map( A1 => n1762, A2 => n1931, B1 => n4671, B2 => 
                           n1586, ZN => n7863);
   U2661 : OAI22_X1 port map( A1 => n1763, A2 => n1931, B1 => n4670, B2 => 
                           n1586, ZN => n7862);
   U2662 : OAI22_X1 port map( A1 => n1764, A2 => n1931, B1 => n4669, B2 => 
                           n1586, ZN => n7861);
   U2663 : OAI22_X1 port map( A1 => n1765, A2 => n1931, B1 => n4668, B2 => 
                           n1586, ZN => n7860);
   U2664 : OAI22_X1 port map( A1 => n1766, A2 => n1931, B1 => n4667, B2 => 
                           n1586, ZN => n7859);
   U2665 : OAI22_X1 port map( A1 => n1767, A2 => n1931, B1 => n4666, B2 => 
                           n1586, ZN => n7858);
   U2666 : OAI22_X1 port map( A1 => n1746, A2 => n1931, B1 => n4665, B2 => 
                           n1586, ZN => n7857);
   U2667 : OAI22_X1 port map( A1 => n1747, A2 => n1931, B1 => n4664, B2 => 
                           n1586, ZN => n7856);
   U2668 : OAI22_X1 port map( A1 => n1742, A2 => n1931, B1 => n4663, B2 => 
                           n1586, ZN => n7855);
   U2669 : OAI22_X1 port map( A1 => n1743, A2 => n1931, B1 => n4662, B2 => 
                           n1586, ZN => n7854);
   U2670 : OAI22_X1 port map( A1 => n1744, A2 => n1931, B1 => n4661, B2 => 
                           n1586, ZN => n7853);
   U2671 : OAI22_X1 port map( A1 => n1745, A2 => n1931, B1 => n4660, B2 => 
                           n1586, ZN => n7852);
   U2672 : OAI22_X1 port map( A1 => n1738, A2 => n1931, B1 => n4659, B2 => 
                           n1586, ZN => n7851);
   U2673 : OAI22_X1 port map( A1 => n1739, A2 => n1931, B1 => n4658, B2 => 
                           n1586, ZN => n7850);
   U2674 : OAI22_X1 port map( A1 => n1740, A2 => n1931, B1 => n4657, B2 => 
                           n1586, ZN => n7849);
   U2675 : OAI22_X1 port map( A1 => n1741, A2 => n1931, B1 => n4656, B2 => 
                           n1586, ZN => n7848);
   U2676 : OAI22_X1 port map( A1 => n1734, A2 => n1931, B1 => n4655, B2 => 
                           n1586, ZN => n7847);
   U2677 : OAI22_X1 port map( A1 => n1735, A2 => n1931, B1 => n4654, B2 => 
                           n1586, ZN => n7846);
   U2678 : OAI22_X1 port map( A1 => n1736, A2 => n1931, B1 => n4653, B2 => 
                           n1586, ZN => n7845);
   U2679 : OAI22_X1 port map( A1 => n1737, A2 => n1931, B1 => n4652, B2 => 
                           n1586, ZN => n7844);
   U2680 : OAI22_X1 port map( A1 => n1730, A2 => n1931, B1 => n4651, B2 => 
                           n1586, ZN => n7843);
   U2681 : OAI22_X1 port map( A1 => n1731, A2 => n1931, B1 => n4650, B2 => 
                           n1586, ZN => n7842);
   U2682 : OAI22_X1 port map( A1 => n1732, A2 => n1931, B1 => n4649, B2 => 
                           n1586, ZN => n7841);
   U2683 : OAI22_X1 port map( A1 => n1733, A2 => n1931, B1 => n4648, B2 => 
                           n1586, ZN => n7840);
   U2684 : OAI22_X1 port map( A1 => n1726, A2 => n1931, B1 => n4647, B2 => 
                           n1586, ZN => n7839);
   U2685 : OAI22_X1 port map( A1 => n1727, A2 => n1931, B1 => n4646, B2 => 
                           n1586, ZN => n7838);
   U2686 : OAI22_X1 port map( A1 => n1728, A2 => n1931, B1 => n4645, B2 => 
                           n1586, ZN => n7837);
   U2687 : OAI22_X1 port map( A1 => n1729, A2 => n1931, B1 => n4644, B2 => 
                           n1586, ZN => n7836);
   U2688 : OAI22_X1 port map( A1 => n1725, A2 => n1931, B1 => n4643, B2 => 
                           n1586, ZN => n7835);
   U2689 : OAI22_X1 port map( A1 => n1768, A2 => n1931, B1 => n4642, B2 => 
                           n1586, ZN => n7834);
   U2690 : OAI21_X1 port map( B1 => n1769, B2 => n1931, A => n1770, ZN => n1932
                           );
   U2691 : AND2_X1 port map( A1 => n1911, A2 => n1928, ZN => n1778);
   U2692 : OAI22_X1 port map( A1 => n1759, A2 => n1933, B1 => n1662, B2 => 
                           n1065, ZN => n7833);
   U2693 : OAI22_X1 port map( A1 => n1761, A2 => n1933, B1 => n1662, B2 => 
                           n1066, ZN => n7832);
   U2694 : OAI22_X1 port map( A1 => n1762, A2 => n1933, B1 => n1662, B2 => 
                           n1067, ZN => n7831);
   U2695 : OAI22_X1 port map( A1 => n1763, A2 => n1933, B1 => n1662, B2 => 
                           n1068, ZN => n7830);
   U2696 : OAI22_X1 port map( A1 => n1764, A2 => n1933, B1 => n1662, B2 => 
                           n1069, ZN => n7829);
   U2697 : OAI22_X1 port map( A1 => n1765, A2 => n1933, B1 => n1662, B2 => 
                           n1070, ZN => n7828);
   U2698 : OAI22_X1 port map( A1 => n1766, A2 => n1933, B1 => n1662, B2 => 
                           n1071, ZN => n7827);
   U2699 : OAI22_X1 port map( A1 => n1767, A2 => n1933, B1 => n1662, B2 => 
                           n1072, ZN => n7826);
   U2700 : OAI22_X1 port map( A1 => n1746, A2 => n1933, B1 => n1662, B2 => 
                           n1073, ZN => n7825);
   U2701 : OAI22_X1 port map( A1 => n1747, A2 => n1933, B1 => n1662, B2 => 
                           n1074, ZN => n7824);
   U2702 : OAI22_X1 port map( A1 => n1742, A2 => n1933, B1 => n1662, B2 => 
                           n1075, ZN => n7823);
   U2703 : OAI22_X1 port map( A1 => n1743, A2 => n1933, B1 => n1662, B2 => 
                           n1076, ZN => n7822);
   U2704 : OAI22_X1 port map( A1 => n1744, A2 => n1933, B1 => n1662, B2 => 
                           n1077, ZN => n7821);
   U2705 : OAI22_X1 port map( A1 => n1745, A2 => n1933, B1 => n1662, B2 => 
                           n1078, ZN => n7820);
   U2706 : OAI22_X1 port map( A1 => n1738, A2 => n1933, B1 => n1662, B2 => 
                           n1079, ZN => n7819);
   U2707 : OAI22_X1 port map( A1 => n1739, A2 => n1933, B1 => n1662, B2 => 
                           n1080, ZN => n7818);
   U2708 : OAI22_X1 port map( A1 => n1740, A2 => n1933, B1 => n1662, B2 => 
                           n1081, ZN => n7817);
   U2709 : OAI22_X1 port map( A1 => n1741, A2 => n1933, B1 => n1662, B2 => 
                           n1082, ZN => n7816);
   U2710 : OAI22_X1 port map( A1 => n1734, A2 => n1933, B1 => n1662, B2 => 
                           n1083, ZN => n7815);
   U2711 : OAI22_X1 port map( A1 => n1735, A2 => n1933, B1 => n1662, B2 => 
                           n1084, ZN => n7814);
   U2712 : OAI22_X1 port map( A1 => n1736, A2 => n1933, B1 => n1662, B2 => 
                           n1085, ZN => n7813);
   U2713 : OAI22_X1 port map( A1 => n1737, A2 => n1933, B1 => n1662, B2 => 
                           n1086, ZN => n7812);
   U2714 : OAI22_X1 port map( A1 => n1730, A2 => n1933, B1 => n1662, B2 => 
                           n1087, ZN => n7811);
   U2715 : OAI22_X1 port map( A1 => n1731, A2 => n1933, B1 => n1662, B2 => 
                           n1088, ZN => n7810);
   U2716 : OAI22_X1 port map( A1 => n1732, A2 => n1933, B1 => n1662, B2 => 
                           n1089, ZN => n7809);
   U2717 : OAI22_X1 port map( A1 => n1733, A2 => n1933, B1 => n1662, B2 => 
                           n1090, ZN => n7808);
   U2718 : OAI22_X1 port map( A1 => n1726, A2 => n1933, B1 => n1662, B2 => 
                           n1091, ZN => n7807);
   U2719 : OAI22_X1 port map( A1 => n1727, A2 => n1933, B1 => n1662, B2 => 
                           n1092, ZN => n7806);
   U2720 : OAI22_X1 port map( A1 => n1728, A2 => n1933, B1 => n1662, B2 => 
                           n1093, ZN => n7805);
   U2721 : OAI22_X1 port map( A1 => n1729, A2 => n1933, B1 => n1662, B2 => 
                           n1094, ZN => n7804);
   U2722 : OAI22_X1 port map( A1 => n1725, A2 => n1933, B1 => n1662, B2 => 
                           n1095, ZN => n7803);
   U2723 : OAI22_X1 port map( A1 => n1768, A2 => n1933, B1 => n1662, B2 => 
                           n1096, ZN => n7802);
   U2724 : OAI21_X1 port map( B1 => n1769, B2 => n1933, A => n1770, ZN => n1934
                           );
   U2725 : AND2_X1 port map( A1 => n1914, A2 => n1928, ZN => n1781);
   U2726 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(3), ZN => n1928);
   U2727 : OAI22_X1 port map( A1 => n1759, A2 => n1935, B1 => n1664, B2 => 
                           n1417, ZN => n7801);
   U2728 : OAI22_X1 port map( A1 => n1761, A2 => n1935, B1 => n1664, B2 => 
                           n1418, ZN => n7800);
   U2729 : OAI22_X1 port map( A1 => n1762, A2 => n1935, B1 => n1664, B2 => 
                           n1419, ZN => n7799);
   U2730 : OAI22_X1 port map( A1 => n1763, A2 => n1935, B1 => n1664, B2 => 
                           n1420, ZN => n7798);
   U2731 : OAI22_X1 port map( A1 => n1764, A2 => n1935, B1 => n1664, B2 => 
                           n1421, ZN => n7797);
   U2732 : OAI22_X1 port map( A1 => n1765, A2 => n1935, B1 => n1664, B2 => 
                           n1422, ZN => n7796);
   U2733 : OAI22_X1 port map( A1 => n1766, A2 => n1935, B1 => n1664, B2 => 
                           n1423, ZN => n7795);
   U2734 : OAI22_X1 port map( A1 => n1767, A2 => n1935, B1 => n1664, B2 => 
                           n1424, ZN => n7794);
   U2735 : OAI22_X1 port map( A1 => n1746, A2 => n1935, B1 => n1664, B2 => 
                           n1425, ZN => n7793);
   U2736 : OAI22_X1 port map( A1 => n1747, A2 => n1935, B1 => n1664, B2 => 
                           n1426, ZN => n7792);
   U2737 : OAI22_X1 port map( A1 => n1742, A2 => n1935, B1 => n1664, B2 => 
                           n1427, ZN => n7791);
   U2738 : OAI22_X1 port map( A1 => n1743, A2 => n1935, B1 => n1664, B2 => 
                           n1428, ZN => n7790);
   U2739 : OAI22_X1 port map( A1 => n1744, A2 => n1935, B1 => n1664, B2 => 
                           n1429, ZN => n7789);
   U2740 : OAI22_X1 port map( A1 => n1745, A2 => n1935, B1 => n1664, B2 => 
                           n1430, ZN => n7788);
   U2741 : OAI22_X1 port map( A1 => n1738, A2 => n1935, B1 => n1664, B2 => 
                           n1431, ZN => n7787);
   U2742 : OAI22_X1 port map( A1 => n1739, A2 => n1935, B1 => n1664, B2 => 
                           n1432, ZN => n7786);
   U2743 : OAI22_X1 port map( A1 => n1740, A2 => n1935, B1 => n1664, B2 => 
                           n1433, ZN => n7785);
   U2744 : OAI22_X1 port map( A1 => n1741, A2 => n1935, B1 => n1664, B2 => 
                           n1434, ZN => n7784);
   U2745 : OAI22_X1 port map( A1 => n1734, A2 => n1935, B1 => n1664, B2 => 
                           n1435, ZN => n7783);
   U2746 : OAI22_X1 port map( A1 => n1735, A2 => n1935, B1 => n1664, B2 => 
                           n1436, ZN => n7782);
   U2747 : OAI22_X1 port map( A1 => n1736, A2 => n1935, B1 => n1664, B2 => 
                           n1437, ZN => n7781);
   U2748 : OAI22_X1 port map( A1 => n1737, A2 => n1935, B1 => n1664, B2 => 
                           n1438, ZN => n7780);
   U2749 : OAI22_X1 port map( A1 => n1730, A2 => n1935, B1 => n1664, B2 => 
                           n1439, ZN => n7779);
   U2750 : OAI22_X1 port map( A1 => n1731, A2 => n1935, B1 => n1664, B2 => 
                           n1440, ZN => n7778);
   U2751 : OAI22_X1 port map( A1 => n1732, A2 => n1935, B1 => n1664, B2 => 
                           n1441, ZN => n7777);
   U2752 : OAI22_X1 port map( A1 => n1733, A2 => n1935, B1 => n1664, B2 => 
                           n1442, ZN => n7776);
   U2753 : OAI22_X1 port map( A1 => n1726, A2 => n1935, B1 => n1664, B2 => 
                           n1443, ZN => n7775);
   U2754 : OAI22_X1 port map( A1 => n1727, A2 => n1935, B1 => n1664, B2 => 
                           n1444, ZN => n7774);
   U2755 : OAI22_X1 port map( A1 => n1728, A2 => n1935, B1 => n1664, B2 => 
                           n1445, ZN => n7773);
   U2756 : OAI22_X1 port map( A1 => n1729, A2 => n1935, B1 => n1664, B2 => 
                           n1446, ZN => n7772);
   U2757 : OAI22_X1 port map( A1 => n1725, A2 => n1935, B1 => n1664, B2 => 
                           n1447, ZN => n7771);
   U2758 : OAI22_X1 port map( A1 => n1768, A2 => n1935, B1 => n1664, B2 => 
                           n1448, ZN => n7770);
   U2759 : OAI21_X1 port map( B1 => n1769, B2 => n1935, A => n1770, ZN => n1936
                           );
   U2760 : AND2_X1 port map( A1 => n1937, A2 => n1905, ZN => n1784);
   U2761 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n1905);
   U2762 : OAI22_X1 port map( A1 => n1759, A2 => n1938, B1 => n4641, B2 => 
                           n1588, ZN => n7769);
   U2763 : OAI22_X1 port map( A1 => n1761, A2 => n1938, B1 => n4640, B2 => 
                           n1588, ZN => n7768);
   U2764 : OAI22_X1 port map( A1 => n1762, A2 => n1938, B1 => n4639, B2 => 
                           n1588, ZN => n7767);
   U2765 : OAI22_X1 port map( A1 => n1763, A2 => n1938, B1 => n4638, B2 => 
                           n1588, ZN => n7766);
   U2766 : OAI22_X1 port map( A1 => n1764, A2 => n1938, B1 => n4637, B2 => 
                           n1588, ZN => n7765);
   U2767 : OAI22_X1 port map( A1 => n1765, A2 => n1938, B1 => n4636, B2 => 
                           n1588, ZN => n7764);
   U2768 : OAI22_X1 port map( A1 => n1766, A2 => n1938, B1 => n4635, B2 => 
                           n1588, ZN => n7763);
   U2769 : OAI22_X1 port map( A1 => n1767, A2 => n1938, B1 => n4634, B2 => 
                           n1588, ZN => n7762);
   U2770 : OAI22_X1 port map( A1 => n1746, A2 => n1938, B1 => n4633, B2 => 
                           n1588, ZN => n7761);
   U2771 : OAI22_X1 port map( A1 => n1747, A2 => n1938, B1 => n4632, B2 => 
                           n1588, ZN => n7760);
   U2772 : OAI22_X1 port map( A1 => n1742, A2 => n1938, B1 => n4631, B2 => 
                           n1588, ZN => n7759);
   U2773 : OAI22_X1 port map( A1 => n1743, A2 => n1938, B1 => n4630, B2 => 
                           n1588, ZN => n7758);
   U2774 : OAI22_X1 port map( A1 => n1744, A2 => n1938, B1 => n4629, B2 => 
                           n1588, ZN => n7757);
   U2775 : OAI22_X1 port map( A1 => n1745, A2 => n1938, B1 => n4628, B2 => 
                           n1588, ZN => n7756);
   U2776 : OAI22_X1 port map( A1 => n1738, A2 => n1938, B1 => n4627, B2 => 
                           n1588, ZN => n7755);
   U2777 : OAI22_X1 port map( A1 => n1739, A2 => n1938, B1 => n4626, B2 => 
                           n1588, ZN => n7754);
   U2778 : OAI22_X1 port map( A1 => n1740, A2 => n1938, B1 => n4625, B2 => 
                           n1588, ZN => n7753);
   U2779 : OAI22_X1 port map( A1 => n1741, A2 => n1938, B1 => n4624, B2 => 
                           n1588, ZN => n7752);
   U2780 : OAI22_X1 port map( A1 => n1734, A2 => n1938, B1 => n4623, B2 => 
                           n1588, ZN => n7751);
   U2781 : OAI22_X1 port map( A1 => n1735, A2 => n1938, B1 => n4622, B2 => 
                           n1588, ZN => n7750);
   U2782 : OAI22_X1 port map( A1 => n1736, A2 => n1938, B1 => n4621, B2 => 
                           n1588, ZN => n7749);
   U2783 : OAI22_X1 port map( A1 => n1737, A2 => n1938, B1 => n4620, B2 => 
                           n1588, ZN => n7748);
   U2784 : OAI22_X1 port map( A1 => n1730, A2 => n1938, B1 => n4619, B2 => 
                           n1588, ZN => n7747);
   U2785 : OAI22_X1 port map( A1 => n1731, A2 => n1938, B1 => n4618, B2 => 
                           n1588, ZN => n7746);
   U2786 : OAI22_X1 port map( A1 => n1732, A2 => n1938, B1 => n4617, B2 => 
                           n1588, ZN => n7745);
   U2787 : OAI22_X1 port map( A1 => n1733, A2 => n1938, B1 => n4616, B2 => 
                           n1588, ZN => n7744);
   U2788 : OAI22_X1 port map( A1 => n1726, A2 => n1938, B1 => n4615, B2 => 
                           n1588, ZN => n7743);
   U2789 : OAI22_X1 port map( A1 => n1727, A2 => n1938, B1 => n4614, B2 => 
                           n1588, ZN => n7742);
   U2790 : OAI22_X1 port map( A1 => n1728, A2 => n1938, B1 => n4613, B2 => 
                           n1588, ZN => n7741);
   U2791 : OAI22_X1 port map( A1 => n1729, A2 => n1938, B1 => n4612, B2 => 
                           n1588, ZN => n7740);
   U2792 : OAI22_X1 port map( A1 => n1725, A2 => n1938, B1 => n4611, B2 => 
                           n1588, ZN => n7739);
   U2793 : OAI22_X1 port map( A1 => n1768, A2 => n1938, B1 => n4610, B2 => 
                           n1588, ZN => n7738);
   U2794 : OAI21_X1 port map( B1 => n1769, B2 => n1938, A => n1770, ZN => n1939
                           );
   U2795 : AND2_X1 port map( A1 => n1937, A2 => n1908, ZN => n1787);
   U2796 : NOR2_X1 port map( A1 => n1940, A2 => ADD_WR(1), ZN => n1908);
   U2797 : OAI22_X1 port map( A1 => n1759, A2 => n1941, B1 => n4609, B2 => 
                           n1582, ZN => n7737);
   U2798 : OAI22_X1 port map( A1 => n1761, A2 => n1941, B1 => n4608, B2 => 
                           n1582, ZN => n7736);
   U2799 : OAI22_X1 port map( A1 => n1762, A2 => n1941, B1 => n4607, B2 => 
                           n1582, ZN => n7735);
   U2800 : OAI22_X1 port map( A1 => n1763, A2 => n1941, B1 => n4606, B2 => 
                           n1582, ZN => n7734);
   U2801 : OAI22_X1 port map( A1 => n1764, A2 => n1941, B1 => n4605, B2 => 
                           n1582, ZN => n7733);
   U2802 : OAI22_X1 port map( A1 => n1765, A2 => n1941, B1 => n4604, B2 => 
                           n1582, ZN => n7732);
   U2803 : OAI22_X1 port map( A1 => n1766, A2 => n1941, B1 => n4603, B2 => 
                           n1582, ZN => n7731);
   U2804 : OAI22_X1 port map( A1 => n1767, A2 => n1941, B1 => n4602, B2 => 
                           n1582, ZN => n7730);
   U2805 : OAI22_X1 port map( A1 => n1746, A2 => n1941, B1 => n4601, B2 => 
                           n1582, ZN => n7729);
   U2806 : OAI22_X1 port map( A1 => n1747, A2 => n1941, B1 => n4600, B2 => 
                           n1582, ZN => n7728);
   U2807 : OAI22_X1 port map( A1 => n1742, A2 => n1941, B1 => n4599, B2 => 
                           n1582, ZN => n7727);
   U2808 : OAI22_X1 port map( A1 => n1743, A2 => n1941, B1 => n4598, B2 => 
                           n1582, ZN => n7726);
   U2809 : OAI22_X1 port map( A1 => n1744, A2 => n1941, B1 => n4597, B2 => 
                           n1582, ZN => n7725);
   U2810 : OAI22_X1 port map( A1 => n1745, A2 => n1941, B1 => n4596, B2 => 
                           n1582, ZN => n7724);
   U2811 : OAI22_X1 port map( A1 => n1738, A2 => n1941, B1 => n4595, B2 => 
                           n1582, ZN => n7723);
   U2812 : OAI22_X1 port map( A1 => n1739, A2 => n1941, B1 => n4594, B2 => 
                           n1582, ZN => n7722);
   U2813 : OAI22_X1 port map( A1 => n1740, A2 => n1941, B1 => n4593, B2 => 
                           n1582, ZN => n7721);
   U2814 : OAI22_X1 port map( A1 => n1741, A2 => n1941, B1 => n4592, B2 => 
                           n1582, ZN => n7720);
   U2815 : OAI22_X1 port map( A1 => n1734, A2 => n1941, B1 => n4591, B2 => 
                           n1582, ZN => n7719);
   U2816 : OAI22_X1 port map( A1 => n1735, A2 => n1941, B1 => n4590, B2 => 
                           n1582, ZN => n7718);
   U2817 : OAI22_X1 port map( A1 => n1736, A2 => n1941, B1 => n4589, B2 => 
                           n1582, ZN => n7717);
   U2818 : OAI22_X1 port map( A1 => n1737, A2 => n1941, B1 => n4588, B2 => 
                           n1582, ZN => n7716);
   U2819 : OAI22_X1 port map( A1 => n1730, A2 => n1941, B1 => n4587, B2 => 
                           n1582, ZN => n7715);
   U2820 : OAI22_X1 port map( A1 => n1731, A2 => n1941, B1 => n4586, B2 => 
                           n1582, ZN => n7714);
   U2821 : OAI22_X1 port map( A1 => n1732, A2 => n1941, B1 => n4585, B2 => 
                           n1582, ZN => n7713);
   U2822 : OAI22_X1 port map( A1 => n1733, A2 => n1941, B1 => n4584, B2 => 
                           n1582, ZN => n7712);
   U2823 : OAI22_X1 port map( A1 => n1726, A2 => n1941, B1 => n4583, B2 => 
                           n1582, ZN => n7711);
   U2824 : OAI22_X1 port map( A1 => n1727, A2 => n1941, B1 => n4582, B2 => 
                           n1582, ZN => n7710);
   U2825 : OAI22_X1 port map( A1 => n1728, A2 => n1941, B1 => n4581, B2 => 
                           n1582, ZN => n7709);
   U2826 : OAI22_X1 port map( A1 => n1729, A2 => n1941, B1 => n4580, B2 => 
                           n1582, ZN => n7708);
   U2827 : OAI22_X1 port map( A1 => n1725, A2 => n1941, B1 => n4579, B2 => 
                           n1582, ZN => n7707);
   U2828 : OAI22_X1 port map( A1 => n1768, A2 => n1941, B1 => n4578, B2 => 
                           n1582, ZN => n7706);
   U2829 : OAI21_X1 port map( B1 => n1769, B2 => n1941, A => n1770, ZN => n1942
                           );
   U2830 : AND2_X1 port map( A1 => n1937, A2 => n1911, ZN => n1790);
   U2831 : NOR2_X1 port map( A1 => n1943, A2 => ADD_WR(0), ZN => n1911);
   U2832 : OAI22_X1 port map( A1 => n4577, A2 => n1584, B1 => n1759, B2 => 
                           n1945, ZN => n7705);
   U2833 : OAI22_X1 port map( A1 => n4576, A2 => n1584, B1 => n1761, B2 => 
                           n1945, ZN => n7704);
   U2834 : OAI22_X1 port map( A1 => n4575, A2 => n1584, B1 => n1762, B2 => 
                           n1945, ZN => n7703);
   U2835 : OAI22_X1 port map( A1 => n4574, A2 => n1584, B1 => n1763, B2 => 
                           n1945, ZN => n7702);
   U2836 : OAI22_X1 port map( A1 => n4573, A2 => n1584, B1 => n1764, B2 => 
                           n1945, ZN => n7701);
   U2837 : OAI22_X1 port map( A1 => n4572, A2 => n1584, B1 => n1765, B2 => 
                           n1945, ZN => n7700);
   U2838 : OAI22_X1 port map( A1 => n4571, A2 => n1584, B1 => n1766, B2 => 
                           n1945, ZN => n7699);
   U2839 : OAI22_X1 port map( A1 => n4570, A2 => n1584, B1 => n1767, B2 => 
                           n1945, ZN => n7698);
   U2840 : OAI22_X1 port map( A1 => n4569, A2 => n1584, B1 => n1746, B2 => 
                           n1945, ZN => n7697);
   U2841 : OAI22_X1 port map( A1 => n4568, A2 => n1584, B1 => n1747, B2 => 
                           n1945, ZN => n7696);
   U2842 : OAI22_X1 port map( A1 => n4567, A2 => n1584, B1 => n1742, B2 => 
                           n1945, ZN => n7695);
   U2843 : OAI22_X1 port map( A1 => n4566, A2 => n1584, B1 => n1743, B2 => 
                           n1945, ZN => n7694);
   U2844 : OAI22_X1 port map( A1 => n4565, A2 => n1584, B1 => n1744, B2 => 
                           n1945, ZN => n7693);
   U2845 : OAI22_X1 port map( A1 => n4564, A2 => n1584, B1 => n1745, B2 => 
                           n1945, ZN => n7692);
   U2846 : OAI22_X1 port map( A1 => n4563, A2 => n1584, B1 => n1738, B2 => 
                           n1945, ZN => n7691);
   U2847 : OAI22_X1 port map( A1 => n4562, A2 => n1584, B1 => n1739, B2 => 
                           n1945, ZN => n7690);
   U2848 : OAI22_X1 port map( A1 => n4561, A2 => n1584, B1 => n1740, B2 => 
                           n1945, ZN => n7689);
   U2849 : OAI22_X1 port map( A1 => n4560, A2 => n1584, B1 => n1741, B2 => 
                           n1945, ZN => n7688);
   U2850 : OAI22_X1 port map( A1 => n4559, A2 => n1584, B1 => n1734, B2 => 
                           n1945, ZN => n7687);
   U2851 : OAI22_X1 port map( A1 => n4558, A2 => n1584, B1 => n1735, B2 => 
                           n1945, ZN => n7686);
   U2852 : OAI22_X1 port map( A1 => n4557, A2 => n1584, B1 => n1736, B2 => 
                           n1945, ZN => n7685);
   U2853 : OAI22_X1 port map( A1 => n4556, A2 => n1584, B1 => n1737, B2 => 
                           n1945, ZN => n7684);
   U2854 : OAI22_X1 port map( A1 => n4555, A2 => n1584, B1 => n1730, B2 => 
                           n1945, ZN => n7683);
   U2855 : OAI22_X1 port map( A1 => n4554, A2 => n1584, B1 => n1731, B2 => 
                           n1945, ZN => n7682);
   U2856 : OAI22_X1 port map( A1 => n4553, A2 => n1584, B1 => n1732, B2 => 
                           n1945, ZN => n7681);
   U2857 : OAI22_X1 port map( A1 => n4552, A2 => n1584, B1 => n1733, B2 => 
                           n1945, ZN => n7680);
   U2858 : OAI22_X1 port map( A1 => n4551, A2 => n1584, B1 => n1726, B2 => 
                           n1945, ZN => n7679);
   U2859 : OAI22_X1 port map( A1 => n4550, A2 => n1584, B1 => n1727, B2 => 
                           n1945, ZN => n7678);
   U2860 : OAI22_X1 port map( A1 => n4549, A2 => n1584, B1 => n1728, B2 => 
                           n1945, ZN => n7677);
   U2861 : OAI22_X1 port map( A1 => n4548, A2 => n1584, B1 => n1729, B2 => 
                           n1945, ZN => n7676);
   U2862 : OAI22_X1 port map( A1 => n4547, A2 => n1584, B1 => n1725, B2 => 
                           n1945, ZN => n7675);
   U2863 : OAI22_X1 port map( A1 => n1768, A2 => n1945, B1 => n4546, B2 => 
                           n1584, ZN => n7674);
   U2864 : OAI21_X1 port map( B1 => n1769, B2 => n1945, A => n1770, ZN => n1944
                           );
   U2865 : AND2_X1 port map( A1 => n1937, A2 => n1914, ZN => n1793);
   U2866 : NOR2_X1 port map( A1 => n1943, A2 => n1940, ZN => n1914);
   U2867 : INV_X1 port map( A => ADD_WR(0), ZN => n1940);
   U2868 : NOR2_X1 port map( A1 => n1915, A2 => ADD_WR(3), ZN => n1937);
   U2869 : AND3_X1 port map( A1 => n1850, A2 => n1884, A3 => ADD_WR(6), ZN => 
                           n1927);
   U2870 : INV_X1 port map( A => ADD_WR(5), ZN => n1884);
   U2871 : INV_X1 port map( A => ADD_WR(4), ZN => n1850);
   U2872 : OAI222_X1 port map( A1 => n1947, A2 => n1948, B1 => n1949, B2 => 
                           n1950, C1 => n1951, C2 => n1449, ZN => n7673);
   U2873 : NOR4_X1 port map( A1 => n1952, A2 => n1953, A3 => n1954, A4 => n1955
                           , ZN => n1949);
   U2874 : NAND4_X1 port map( A1 => n1956, A2 => n1957, A3 => n1958, A4 => 
                           n1959, ZN => n1955);
   U2875 : AOI221_X1 port map( B1 => n1960, B2 => n6433, C1 => n1961, C2 => 
                           n6465, A => n1962, ZN => n1959);
   U2876 : OAI222_X1 port map( A1 => n5281, A2 => n1963, B1 => n5249, B2 => 
                           n1964, C1 => n5217, C2 => n1965, ZN => n1962);
   U2877 : AOI221_X1 port map( B1 => n1966, B2 => n6497, C1 => n1967, C2 => 
                           n6529, A => n1968, ZN => n1958);
   U2878 : OAI22_X1 port map( A1 => n5694, A2 => n1969, B1 => n5695, B2 => 
                           n1970, ZN => n1968);
   U2879 : AOI221_X1 port map( B1 => n1971, B2 => n6561, C1 => n1972, C2 => 
                           n6593, A => n1973, ZN => n1957);
   U2880 : OAI222_X1 port map( A1 => n5377, A2 => n1974, B1 => n5345, B2 => 
                           n1578, C1 => n5313, C2 => n1975, ZN => n1973);
   U2881 : AOI221_X1 port map( B1 => n1976, B2 => n6625, C1 => n1977, C2 => 
                           n6657, A => n1978, ZN => n1956);
   U2882 : OAI22_X1 port map( A1 => n5696, A2 => n1756, B1 => n5697, B2 => 
                           n1980, ZN => n1978);
   U2883 : NAND4_X1 port map( A1 => n1981, A2 => n1982, A3 => n1983, A4 => 
                           n1984, ZN => n1954);
   U2884 : AOI221_X1 port map( B1 => n1985, B2 => n6305, C1 => n1986, C2 => 
                           n6337, A => n1987, ZN => n1984);
   U2885 : OAI222_X1 port map( A1 => n5089, A2 => n1988, B1 => n5057, B2 => 
                           n1989, C1 => n5025, C2 => n416, ZN => n1987);
   U2886 : AOI221_X1 port map( B1 => n1990, B2 => n161, C1 => n1991, C2 => n521
                           , A => n1992, ZN => n1983);
   U2887 : OAI22_X1 port map( A1 => n65, A2 => n1993, B1 => n425, B2 => n1994, 
                           ZN => n1992);
   U2888 : AOI221_X1 port map( B1 => n1995, B2 => n6369, C1 => n1996, C2 => 
                           n6401, A => n1997, ZN => n1982);
   U2889 : OAI222_X1 port map( A1 => n5185, A2 => n1998, B1 => n5153, B2 => 
                           n1999, C1 => n5121, C2 => n417, ZN => n1997);
   U2890 : AOI221_X1 port map( B1 => n2000, B2 => n553, C1 => n2001, C2 => n97,
                           A => n2002, ZN => n1981);
   U2891 : OAI22_X1 port map( A1 => n1, A2 => n412, B1 => n457, B2 => n2003, ZN
                           => n2002);
   U2892 : NAND4_X1 port map( A1 => n2004, A2 => n2005, A3 => n2006, A4 => 
                           n2007, ZN => n1953);
   U2893 : AOI221_X1 port map( B1 => n2008, B2 => n6113, C1 => n2009, C2 => 
                           n6145, A => n2010, ZN => n2007);
   U2894 : OAI222_X1 port map( A1 => n4897, A2 => n2011, B1 => n4865, B2 => 
                           n2012, C1 => n4833, C2 => n418, ZN => n2010);
   U2895 : AOI221_X1 port map( B1 => n2013, B2 => n6177, C1 => n2014, C2 => 
                           n6209, A => n2015, ZN => n2006);
   U2896 : OAI22_X1 port map( A1 => n5690, A2 => n2016, B1 => n5691, B2 => 
                           n2017, ZN => n2015);
   U2897 : AOI221_X1 port map( B1 => n1751, B2 => n6241, C1 => n2019, C2 => 
                           n6273, A => n2020, ZN => n2005);
   U2898 : OAI222_X1 port map( A1 => n4993, A2 => n2021, B1 => n4961, B2 => 
                           n2022, C1 => n4929, C2 => n419, ZN => n2020);
   U2899 : AOI221_X1 port map( B1 => n2023, B2 => n554, C1 => n2024, C2 => n98,
                           A => n2025, ZN => n2004);
   U2900 : OAI22_X1 port map( A1 => n2, A2 => n2026, B1 => n458, B2 => n2027, 
                           ZN => n2025);
   U2901 : NAND4_X1 port map( A1 => n2028, A2 => n2029, A3 => n2030, A4 => 
                           n2031, ZN => n1952);
   U2902 : AOI221_X1 port map( B1 => n2032, B2 => n5857, C1 => n2033, C2 => 
                           n5889, A => n2034, ZN => n2031);
   U2903 : OAI222_X1 port map( A1 => n4641, A2 => n2035, B1 => n4609, B2 => 
                           n2036, C1 => n4577, C2 => n1577, ZN => n2034);
   U2904 : AOI221_X1 port map( B1 => n2037, B2 => n5921, C1 => n2038, C2 => 
                           n5953, A => n2039, ZN => n2030);
   U2905 : OAI22_X1 port map( A1 => n4705, A2 => n2040, B1 => n4673, B2 => 
                           n2041, ZN => n2039);
   U2906 : AOI221_X1 port map( B1 => n1752, B2 => n5985, C1 => n2043, C2 => 
                           n6017, A => n2044, ZN => n2029);
   U2907 : OAI222_X1 port map( A1 => n4801, A2 => n411, B1 => n4769, B2 => 
                           n2045, C1 => n4737, C2 => n2046, ZN => n2044);
   U2908 : AOI221_X1 port map( B1 => n1749, B2 => n6049, C1 => n2048, C2 => 
                           n6081, A => n2049, ZN => n2028);
   U2909 : OAI22_X1 port map( A1 => n5688, A2 => n2050, B1 => n5689, B2 => 
                           n2051, ZN => n2049);
   U2910 : OAI21_X1 port map( B1 => n1951, B2 => n1513, A => ENABLE, ZN => 
                           n7672);
   U2911 : OAI222_X1 port map( A1 => n2052, A2 => n1948, B1 => n2053, B2 => 
                           n1950, C1 => n1951, C2 => n1450, ZN => n7671);
   U2912 : NOR4_X1 port map( A1 => n2054, A2 => n2055, A3 => n2056, A4 => n2057
                           , ZN => n2053);
   U2913 : NAND4_X1 port map( A1 => n2058, A2 => n2059, A3 => n2060, A4 => 
                           n2061, ZN => n2057);
   U2914 : AOI221_X1 port map( B1 => n1960, B2 => n6432, C1 => n1961, C2 => 
                           n6464, A => n2062, ZN => n2061);
   U2915 : OAI222_X1 port map( A1 => n5280, A2 => n1963, B1 => n5248, B2 => 
                           n1964, C1 => n5216, C2 => n1965, ZN => n2062);
   U2916 : AOI221_X1 port map( B1 => n1966, B2 => n6496, C1 => n1967, C2 => 
                           n6528, A => n2063, ZN => n2060);
   U2917 : OAI22_X1 port map( A1 => n5684, A2 => n1969, B1 => n5685, B2 => 
                           n1970, ZN => n2063);
   U2918 : AOI221_X1 port map( B1 => n1971, B2 => n6560, C1 => n1972, C2 => 
                           n6592, A => n2064, ZN => n2059);
   U2919 : OAI222_X1 port map( A1 => n5376, A2 => n1974, B1 => n5344, B2 => 
                           n1578, C1 => n5312, C2 => n1975, ZN => n2064);
   U2920 : AOI221_X1 port map( B1 => n1976, B2 => n6624, C1 => n1977, C2 => 
                           n6656, A => n2065, ZN => n2058);
   U2921 : OAI22_X1 port map( A1 => n5686, A2 => n1756, B1 => n5687, B2 => 
                           n1980, ZN => n2065);
   U2922 : NAND4_X1 port map( A1 => n2066, A2 => n2067, A3 => n2068, A4 => 
                           n2069, ZN => n2056);
   U2923 : AOI221_X1 port map( B1 => n1985, B2 => n6304, C1 => n1986, C2 => 
                           n6336, A => n2070, ZN => n2069);
   U2924 : OAI222_X1 port map( A1 => n5088, A2 => n1988, B1 => n5056, B2 => 
                           n1989, C1 => n5024, C2 => n416, ZN => n2070);
   U2925 : AOI221_X1 port map( B1 => n1990, B2 => n162, C1 => n1991, C2 => n522
                           , A => n2071, ZN => n2068);
   U2926 : OAI22_X1 port map( A1 => n66, A2 => n1993, B1 => n426, B2 => n1994, 
                           ZN => n2071);
   U2927 : AOI221_X1 port map( B1 => n1995, B2 => n6368, C1 => n1996, C2 => 
                           n6400, A => n2072, ZN => n2067);
   U2928 : OAI222_X1 port map( A1 => n5184, A2 => n1998, B1 => n5152, B2 => 
                           n1999, C1 => n5120, C2 => n417, ZN => n2072);
   U2929 : AOI221_X1 port map( B1 => n2000, B2 => n555, C1 => n2001, C2 => n99,
                           A => n2073, ZN => n2066);
   U2930 : OAI22_X1 port map( A1 => n3, A2 => n412, B1 => n459, B2 => n2003, ZN
                           => n2073);
   U2931 : NAND4_X1 port map( A1 => n2074, A2 => n2075, A3 => n2076, A4 => 
                           n2077, ZN => n2055);
   U2932 : AOI221_X1 port map( B1 => n2008, B2 => n6112, C1 => n2009, C2 => 
                           n6144, A => n2078, ZN => n2077);
   U2933 : OAI222_X1 port map( A1 => n4896, A2 => n2011, B1 => n4864, B2 => 
                           n2012, C1 => n4832, C2 => n418, ZN => n2078);
   U2934 : AOI221_X1 port map( B1 => n2013, B2 => n6176, C1 => n2014, C2 => 
                           n6208, A => n2079, ZN => n2076);
   U2935 : OAI22_X1 port map( A1 => n5680, A2 => n2016, B1 => n5681, B2 => 
                           n2017, ZN => n2079);
   U2936 : AOI221_X1 port map( B1 => n1751, B2 => n6240, C1 => n2019, C2 => 
                           n6272, A => n2080, ZN => n2075);
   U2937 : OAI222_X1 port map( A1 => n4992, A2 => n2021, B1 => n4960, B2 => 
                           n2022, C1 => n4928, C2 => n419, ZN => n2080);
   U2938 : AOI221_X1 port map( B1 => n2023, B2 => n556, C1 => n2024, C2 => n100
                           , A => n2081, ZN => n2074);
   U2939 : OAI22_X1 port map( A1 => n4, A2 => n2026, B1 => n460, B2 => n2027, 
                           ZN => n2081);
   U2940 : NAND4_X1 port map( A1 => n2082, A2 => n2083, A3 => n2084, A4 => 
                           n2085, ZN => n2054);
   U2941 : AOI221_X1 port map( B1 => n2032, B2 => n5856, C1 => n2033, C2 => 
                           n5888, A => n2086, ZN => n2085);
   U2942 : OAI222_X1 port map( A1 => n4640, A2 => n2035, B1 => n4608, B2 => 
                           n2036, C1 => n4576, C2 => n1577, ZN => n2086);
   U2943 : AOI221_X1 port map( B1 => n2037, B2 => n5920, C1 => n2038, C2 => 
                           n5952, A => n2087, ZN => n2084);
   U2944 : OAI22_X1 port map( A1 => n4704, A2 => n2040, B1 => n4672, B2 => 
                           n2041, ZN => n2087);
   U2945 : AOI221_X1 port map( B1 => n1752, B2 => n5984, C1 => n2043, C2 => 
                           n6016, A => n2088, ZN => n2083);
   U2946 : OAI222_X1 port map( A1 => n4800, A2 => n411, B1 => n4768, B2 => 
                           n2045, C1 => n4736, C2 => n2046, ZN => n2088);
   U2947 : AOI221_X1 port map( B1 => n1749, B2 => n6048, C1 => n2048, C2 => 
                           n6080, A => n2089, ZN => n2082);
   U2948 : OAI22_X1 port map( A1 => n5678, A2 => n2050, B1 => n5679, B2 => 
                           n2051, ZN => n2089);
   U2949 : OAI21_X1 port map( B1 => n1951, B2 => n1514, A => ENABLE, ZN => 
                           n7670);
   U2950 : OAI222_X1 port map( A1 => n2090, A2 => n1948, B1 => n2091, B2 => 
                           n1950, C1 => n1951, C2 => n1451, ZN => n7669);
   U2951 : NOR4_X1 port map( A1 => n2092, A2 => n2093, A3 => n2094, A4 => n2095
                           , ZN => n2091);
   U2952 : NAND4_X1 port map( A1 => n2096, A2 => n2097, A3 => n2098, A4 => 
                           n2099, ZN => n2095);
   U2953 : AOI221_X1 port map( B1 => n1960, B2 => n6431, C1 => n1961, C2 => 
                           n6463, A => n2100, ZN => n2099);
   U2954 : OAI222_X1 port map( A1 => n5279, A2 => n1963, B1 => n5247, B2 => 
                           n1964, C1 => n5215, C2 => n1965, ZN => n2100);
   U2955 : AOI221_X1 port map( B1 => n1966, B2 => n6495, C1 => n1967, C2 => 
                           n6527, A => n2101, ZN => n2098);
   U2956 : OAI22_X1 port map( A1 => n5674, A2 => n1969, B1 => n5675, B2 => 
                           n1970, ZN => n2101);
   U2957 : AOI221_X1 port map( B1 => n1971, B2 => n6559, C1 => n1972, C2 => 
                           n6591, A => n2102, ZN => n2097);
   U2958 : OAI222_X1 port map( A1 => n5375, A2 => n1974, B1 => n5343, B2 => 
                           n1578, C1 => n5311, C2 => n1975, ZN => n2102);
   U2959 : AOI221_X1 port map( B1 => n1976, B2 => n6623, C1 => n1977, C2 => 
                           n6655, A => n2103, ZN => n2096);
   U2960 : OAI22_X1 port map( A1 => n5676, A2 => n1756, B1 => n5677, B2 => 
                           n1980, ZN => n2103);
   U2961 : NAND4_X1 port map( A1 => n2104, A2 => n2105, A3 => n2106, A4 => 
                           n2107, ZN => n2094);
   U2962 : AOI221_X1 port map( B1 => n1985, B2 => n6303, C1 => n1986, C2 => 
                           n6335, A => n2108, ZN => n2107);
   U2963 : OAI222_X1 port map( A1 => n5087, A2 => n1988, B1 => n5055, B2 => 
                           n1989, C1 => n5023, C2 => n416, ZN => n2108);
   U2964 : AOI221_X1 port map( B1 => n1990, B2 => n163, C1 => n1991, C2 => n523
                           , A => n2109, ZN => n2106);
   U2965 : OAI22_X1 port map( A1 => n67, A2 => n1993, B1 => n427, B2 => n1994, 
                           ZN => n2109);
   U2966 : AOI221_X1 port map( B1 => n1995, B2 => n6367, C1 => n1996, C2 => 
                           n6399, A => n2110, ZN => n2105);
   U2967 : OAI222_X1 port map( A1 => n5183, A2 => n1998, B1 => n5151, B2 => 
                           n1999, C1 => n5119, C2 => n417, ZN => n2110);
   U2968 : AOI221_X1 port map( B1 => n2000, B2 => n557, C1 => n2001, C2 => n101
                           , A => n2111, ZN => n2104);
   U2969 : OAI22_X1 port map( A1 => n5, A2 => n412, B1 => n461, B2 => n2003, ZN
                           => n2111);
   U2970 : NAND4_X1 port map( A1 => n2112, A2 => n2113, A3 => n2114, A4 => 
                           n2115, ZN => n2093);
   U2971 : AOI221_X1 port map( B1 => n2008, B2 => n6111, C1 => n2009, C2 => 
                           n6143, A => n2116, ZN => n2115);
   U2972 : OAI222_X1 port map( A1 => n4895, A2 => n2011, B1 => n4863, B2 => 
                           n2012, C1 => n4831, C2 => n418, ZN => n2116);
   U2973 : AOI221_X1 port map( B1 => n2013, B2 => n6175, C1 => n2014, C2 => 
                           n6207, A => n2117, ZN => n2114);
   U2974 : OAI22_X1 port map( A1 => n5670, A2 => n2016, B1 => n5671, B2 => 
                           n2017, ZN => n2117);
   U2975 : AOI221_X1 port map( B1 => n1751, B2 => n6239, C1 => n2019, C2 => 
                           n6271, A => n2118, ZN => n2113);
   U2976 : OAI222_X1 port map( A1 => n4991, A2 => n2021, B1 => n4959, B2 => 
                           n2022, C1 => n4927, C2 => n419, ZN => n2118);
   U2977 : AOI221_X1 port map( B1 => n2023, B2 => n558, C1 => n2024, C2 => n102
                           , A => n2119, ZN => n2112);
   U2978 : OAI22_X1 port map( A1 => n6, A2 => n2026, B1 => n462, B2 => n2027, 
                           ZN => n2119);
   U2979 : NAND4_X1 port map( A1 => n2120, A2 => n2121, A3 => n2122, A4 => 
                           n2123, ZN => n2092);
   U2980 : AOI221_X1 port map( B1 => n2032, B2 => n5855, C1 => n2033, C2 => 
                           n5887, A => n2124, ZN => n2123);
   U2981 : OAI222_X1 port map( A1 => n4639, A2 => n2035, B1 => n4607, B2 => 
                           n2036, C1 => n4575, C2 => n1577, ZN => n2124);
   U2982 : AOI221_X1 port map( B1 => n2037, B2 => n5919, C1 => n2038, C2 => 
                           n5951, A => n2125, ZN => n2122);
   U2983 : OAI22_X1 port map( A1 => n4703, A2 => n2040, B1 => n4671, B2 => 
                           n2041, ZN => n2125);
   U2984 : AOI221_X1 port map( B1 => n1752, B2 => n5983, C1 => n2043, C2 => 
                           n6015, A => n2126, ZN => n2121);
   U2985 : OAI222_X1 port map( A1 => n4799, A2 => n411, B1 => n4767, B2 => 
                           n2045, C1 => n4735, C2 => n2046, ZN => n2126);
   U2986 : AOI221_X1 port map( B1 => n1749, B2 => n6047, C1 => n2048, C2 => 
                           n6079, A => n2127, ZN => n2120);
   U2987 : OAI22_X1 port map( A1 => n5668, A2 => n2050, B1 => n5669, B2 => 
                           n2051, ZN => n2127);
   U2988 : OAI21_X1 port map( B1 => n1951, B2 => n1515, A => ENABLE, ZN => 
                           n7668);
   U2989 : OAI222_X1 port map( A1 => n2128, A2 => n1948, B1 => n2129, B2 => 
                           n1950, C1 => n1951, C2 => n1452, ZN => n7667);
   U2990 : NOR4_X1 port map( A1 => n2130, A2 => n2131, A3 => n2132, A4 => n2133
                           , ZN => n2129);
   U2991 : NAND4_X1 port map( A1 => n2134, A2 => n2135, A3 => n2136, A4 => 
                           n2137, ZN => n2133);
   U2992 : AOI221_X1 port map( B1 => n1960, B2 => n6430, C1 => n1961, C2 => 
                           n6462, A => n2138, ZN => n2137);
   U2993 : OAI222_X1 port map( A1 => n5278, A2 => n1963, B1 => n5246, B2 => 
                           n1964, C1 => n5214, C2 => n1965, ZN => n2138);
   U2994 : AOI221_X1 port map( B1 => n1966, B2 => n6494, C1 => n1967, C2 => 
                           n6526, A => n2139, ZN => n2136);
   U2995 : OAI22_X1 port map( A1 => n5664, A2 => n1969, B1 => n5665, B2 => 
                           n1970, ZN => n2139);
   U2996 : AOI221_X1 port map( B1 => n1971, B2 => n6558, C1 => n1972, C2 => 
                           n6590, A => n2140, ZN => n2135);
   U2997 : OAI222_X1 port map( A1 => n5374, A2 => n1974, B1 => n5342, B2 => 
                           n1578, C1 => n5310, C2 => n1975, ZN => n2140);
   U2998 : AOI221_X1 port map( B1 => n1976, B2 => n6622, C1 => n1977, C2 => 
                           n6654, A => n2141, ZN => n2134);
   U2999 : OAI22_X1 port map( A1 => n5666, A2 => n1756, B1 => n5667, B2 => 
                           n1980, ZN => n2141);
   U3000 : NAND4_X1 port map( A1 => n2142, A2 => n2143, A3 => n2144, A4 => 
                           n2145, ZN => n2132);
   U3001 : AOI221_X1 port map( B1 => n1985, B2 => n6302, C1 => n1986, C2 => 
                           n6334, A => n2146, ZN => n2145);
   U3002 : OAI222_X1 port map( A1 => n5086, A2 => n1988, B1 => n5054, B2 => 
                           n1989, C1 => n5022, C2 => n416, ZN => n2146);
   U3003 : AOI221_X1 port map( B1 => n1990, B2 => n164, C1 => n1991, C2 => n524
                           , A => n2147, ZN => n2144);
   U3004 : OAI22_X1 port map( A1 => n68, A2 => n1993, B1 => n428, B2 => n1994, 
                           ZN => n2147);
   U3005 : AOI221_X1 port map( B1 => n1995, B2 => n6366, C1 => n1996, C2 => 
                           n6398, A => n2148, ZN => n2143);
   U3006 : OAI222_X1 port map( A1 => n5182, A2 => n1998, B1 => n5150, B2 => 
                           n1999, C1 => n5118, C2 => n417, ZN => n2148);
   U3007 : AOI221_X1 port map( B1 => n2000, B2 => n559, C1 => n2001, C2 => n103
                           , A => n2149, ZN => n2142);
   U3008 : OAI22_X1 port map( A1 => n7, A2 => n412, B1 => n463, B2 => n2003, ZN
                           => n2149);
   U3009 : NAND4_X1 port map( A1 => n2150, A2 => n2151, A3 => n2152, A4 => 
                           n2153, ZN => n2131);
   U3010 : AOI221_X1 port map( B1 => n2008, B2 => n6110, C1 => n2009, C2 => 
                           n6142, A => n2154, ZN => n2153);
   U3011 : OAI222_X1 port map( A1 => n4894, A2 => n2011, B1 => n4862, B2 => 
                           n2012, C1 => n4830, C2 => n418, ZN => n2154);
   U3012 : AOI221_X1 port map( B1 => n2013, B2 => n6174, C1 => n2014, C2 => 
                           n6206, A => n2155, ZN => n2152);
   U3013 : OAI22_X1 port map( A1 => n5660, A2 => n2016, B1 => n5661, B2 => 
                           n2017, ZN => n2155);
   U3014 : AOI221_X1 port map( B1 => n1751, B2 => n6238, C1 => n2019, C2 => 
                           n6270, A => n2156, ZN => n2151);
   U3015 : OAI222_X1 port map( A1 => n4990, A2 => n2021, B1 => n4958, B2 => 
                           n2022, C1 => n4926, C2 => n419, ZN => n2156);
   U3016 : AOI221_X1 port map( B1 => n2023, B2 => n560, C1 => n2024, C2 => n104
                           , A => n2157, ZN => n2150);
   U3017 : OAI22_X1 port map( A1 => n8, A2 => n2026, B1 => n464, B2 => n2027, 
                           ZN => n2157);
   U3018 : NAND4_X1 port map( A1 => n2158, A2 => n2159, A3 => n2160, A4 => 
                           n2161, ZN => n2130);
   U3019 : AOI221_X1 port map( B1 => n2032, B2 => n5854, C1 => n2033, C2 => 
                           n5886, A => n2162, ZN => n2161);
   U3020 : OAI222_X1 port map( A1 => n4638, A2 => n2035, B1 => n4606, B2 => 
                           n2036, C1 => n4574, C2 => n1577, ZN => n2162);
   U3021 : AOI221_X1 port map( B1 => n2037, B2 => n5918, C1 => n2038, C2 => 
                           n5950, A => n2163, ZN => n2160);
   U3022 : OAI22_X1 port map( A1 => n4702, A2 => n2040, B1 => n4670, B2 => 
                           n2041, ZN => n2163);
   U3023 : AOI221_X1 port map( B1 => n1752, B2 => n5982, C1 => n2043, C2 => 
                           n6014, A => n2164, ZN => n2159);
   U3024 : OAI222_X1 port map( A1 => n4798, A2 => n411, B1 => n4766, B2 => 
                           n2045, C1 => n4734, C2 => n2046, ZN => n2164);
   U3025 : AOI221_X1 port map( B1 => n1749, B2 => n6046, C1 => n2048, C2 => 
                           n6078, A => n2165, ZN => n2158);
   U3026 : OAI22_X1 port map( A1 => n5658, A2 => n2050, B1 => n5659, B2 => 
                           n2051, ZN => n2165);
   U3027 : OAI21_X1 port map( B1 => n1951, B2 => n1516, A => ENABLE, ZN => 
                           n7666);
   U3028 : OAI222_X1 port map( A1 => n2166, A2 => n1948, B1 => n2167, B2 => 
                           n1950, C1 => n1951, C2 => n1453, ZN => n7665);
   U3029 : NOR4_X1 port map( A1 => n2168, A2 => n2169, A3 => n2170, A4 => n2171
                           , ZN => n2167);
   U3030 : NAND4_X1 port map( A1 => n2172, A2 => n2173, A3 => n2174, A4 => 
                           n2175, ZN => n2171);
   U3031 : AOI221_X1 port map( B1 => n1960, B2 => n6429, C1 => n1961, C2 => 
                           n6461, A => n2176, ZN => n2175);
   U3032 : OAI222_X1 port map( A1 => n5277, A2 => n1963, B1 => n5245, B2 => 
                           n1964, C1 => n5213, C2 => n1965, ZN => n2176);
   U3033 : AOI221_X1 port map( B1 => n1966, B2 => n6493, C1 => n1967, C2 => 
                           n6525, A => n2177, ZN => n2174);
   U3034 : OAI22_X1 port map( A1 => n5654, A2 => n1969, B1 => n5655, B2 => 
                           n1970, ZN => n2177);
   U3035 : AOI221_X1 port map( B1 => n1971, B2 => n6557, C1 => n1972, C2 => 
                           n6589, A => n2178, ZN => n2173);
   U3036 : OAI222_X1 port map( A1 => n5373, A2 => n1974, B1 => n5341, B2 => 
                           n1578, C1 => n5309, C2 => n1975, ZN => n2178);
   U3037 : AOI221_X1 port map( B1 => n1976, B2 => n6621, C1 => n1977, C2 => 
                           n6653, A => n2179, ZN => n2172);
   U3038 : OAI22_X1 port map( A1 => n5656, A2 => n1756, B1 => n5657, B2 => 
                           n1980, ZN => n2179);
   U3039 : NAND4_X1 port map( A1 => n2180, A2 => n2181, A3 => n2182, A4 => 
                           n2183, ZN => n2170);
   U3040 : AOI221_X1 port map( B1 => n1985, B2 => n6301, C1 => n1986, C2 => 
                           n6333, A => n2184, ZN => n2183);
   U3041 : OAI222_X1 port map( A1 => n5085, A2 => n1988, B1 => n5053, B2 => 
                           n1989, C1 => n5021, C2 => n416, ZN => n2184);
   U3042 : AOI221_X1 port map( B1 => n1990, B2 => n165, C1 => n1991, C2 => n525
                           , A => n2185, ZN => n2182);
   U3043 : OAI22_X1 port map( A1 => n69, A2 => n1993, B1 => n429, B2 => n1994, 
                           ZN => n2185);
   U3044 : AOI221_X1 port map( B1 => n1995, B2 => n6365, C1 => n1996, C2 => 
                           n6397, A => n2186, ZN => n2181);
   U3045 : OAI222_X1 port map( A1 => n5181, A2 => n1998, B1 => n5149, B2 => 
                           n1999, C1 => n5117, C2 => n417, ZN => n2186);
   U3046 : AOI221_X1 port map( B1 => n2000, B2 => n561, C1 => n2001, C2 => n105
                           , A => n2187, ZN => n2180);
   U3047 : OAI22_X1 port map( A1 => n9, A2 => n412, B1 => n465, B2 => n2003, ZN
                           => n2187);
   U3048 : NAND4_X1 port map( A1 => n2188, A2 => n2189, A3 => n2190, A4 => 
                           n2191, ZN => n2169);
   U3049 : AOI221_X1 port map( B1 => n2008, B2 => n6109, C1 => n2009, C2 => 
                           n6141, A => n2192, ZN => n2191);
   U3050 : OAI222_X1 port map( A1 => n4893, A2 => n2011, B1 => n4861, B2 => 
                           n2012, C1 => n4829, C2 => n418, ZN => n2192);
   U3051 : AOI221_X1 port map( B1 => n2013, B2 => n6173, C1 => n2014, C2 => 
                           n6205, A => n2193, ZN => n2190);
   U3052 : OAI22_X1 port map( A1 => n5650, A2 => n2016, B1 => n5651, B2 => 
                           n2017, ZN => n2193);
   U3053 : AOI221_X1 port map( B1 => n1751, B2 => n6237, C1 => n2019, C2 => 
                           n6269, A => n2194, ZN => n2189);
   U3054 : OAI222_X1 port map( A1 => n4989, A2 => n2021, B1 => n4957, B2 => 
                           n2022, C1 => n4925, C2 => n419, ZN => n2194);
   U3055 : AOI221_X1 port map( B1 => n2023, B2 => n562, C1 => n2024, C2 => n106
                           , A => n2195, ZN => n2188);
   U3056 : OAI22_X1 port map( A1 => n10, A2 => n2026, B1 => n466, B2 => n2027, 
                           ZN => n2195);
   U3057 : NAND4_X1 port map( A1 => n2196, A2 => n2197, A3 => n2198, A4 => 
                           n2199, ZN => n2168);
   U3058 : AOI221_X1 port map( B1 => n2032, B2 => n5853, C1 => n2033, C2 => 
                           n5885, A => n2200, ZN => n2199);
   U3059 : OAI222_X1 port map( A1 => n4637, A2 => n2035, B1 => n4605, B2 => 
                           n2036, C1 => n4573, C2 => n1577, ZN => n2200);
   U3060 : AOI221_X1 port map( B1 => n2037, B2 => n5917, C1 => n2038, C2 => 
                           n5949, A => n2201, ZN => n2198);
   U3061 : OAI22_X1 port map( A1 => n4701, A2 => n2040, B1 => n4669, B2 => 
                           n2041, ZN => n2201);
   U3062 : AOI221_X1 port map( B1 => n1752, B2 => n5981, C1 => n2043, C2 => 
                           n6013, A => n2202, ZN => n2197);
   U3063 : OAI222_X1 port map( A1 => n4797, A2 => n411, B1 => n4765, B2 => 
                           n2045, C1 => n4733, C2 => n2046, ZN => n2202);
   U3064 : AOI221_X1 port map( B1 => n1749, B2 => n6045, C1 => n2048, C2 => 
                           n6077, A => n2203, ZN => n2196);
   U3065 : OAI22_X1 port map( A1 => n5648, A2 => n2050, B1 => n5649, B2 => 
                           n2051, ZN => n2203);
   U3066 : OAI21_X1 port map( B1 => n1951, B2 => n1517, A => ENABLE, ZN => 
                           n7664);
   U3067 : OAI222_X1 port map( A1 => n2204, A2 => n1948, B1 => n2205, B2 => 
                           n1950, C1 => n1951, C2 => n1454, ZN => n7663);
   U3068 : NOR4_X1 port map( A1 => n2206, A2 => n2207, A3 => n2208, A4 => n2209
                           , ZN => n2205);
   U3069 : NAND4_X1 port map( A1 => n2210, A2 => n2211, A3 => n2212, A4 => 
                           n2213, ZN => n2209);
   U3070 : AOI221_X1 port map( B1 => n1960, B2 => n6428, C1 => n1961, C2 => 
                           n6460, A => n2214, ZN => n2213);
   U3071 : OAI222_X1 port map( A1 => n5276, A2 => n1963, B1 => n5244, B2 => 
                           n1964, C1 => n5212, C2 => n1965, ZN => n2214);
   U3072 : AOI221_X1 port map( B1 => n1966, B2 => n6492, C1 => n1967, C2 => 
                           n6524, A => n2215, ZN => n2212);
   U3073 : OAI22_X1 port map( A1 => n5644, A2 => n1969, B1 => n5645, B2 => 
                           n1970, ZN => n2215);
   U3074 : AOI221_X1 port map( B1 => n1971, B2 => n6556, C1 => n1972, C2 => 
                           n6588, A => n2216, ZN => n2211);
   U3075 : OAI222_X1 port map( A1 => n5372, A2 => n1974, B1 => n5340, B2 => 
                           n1578, C1 => n5308, C2 => n1975, ZN => n2216);
   U3076 : AOI221_X1 port map( B1 => n1976, B2 => n6620, C1 => n1977, C2 => 
                           n6652, A => n2217, ZN => n2210);
   U3077 : OAI22_X1 port map( A1 => n5646, A2 => n1756, B1 => n5647, B2 => 
                           n1980, ZN => n2217);
   U3078 : NAND4_X1 port map( A1 => n2218, A2 => n2219, A3 => n2220, A4 => 
                           n2221, ZN => n2208);
   U3079 : AOI221_X1 port map( B1 => n1985, B2 => n6300, C1 => n1986, C2 => 
                           n6332, A => n2222, ZN => n2221);
   U3080 : OAI222_X1 port map( A1 => n5084, A2 => n1988, B1 => n5052, B2 => 
                           n1989, C1 => n5020, C2 => n416, ZN => n2222);
   U3081 : AOI221_X1 port map( B1 => n1990, B2 => n166, C1 => n1991, C2 => n526
                           , A => n2223, ZN => n2220);
   U3082 : OAI22_X1 port map( A1 => n70, A2 => n1993, B1 => n430, B2 => n1994, 
                           ZN => n2223);
   U3083 : AOI221_X1 port map( B1 => n1995, B2 => n6364, C1 => n1996, C2 => 
                           n6396, A => n2224, ZN => n2219);
   U3084 : OAI222_X1 port map( A1 => n5180, A2 => n1998, B1 => n5148, B2 => 
                           n1999, C1 => n5116, C2 => n417, ZN => n2224);
   U3085 : AOI221_X1 port map( B1 => n2000, B2 => n563, C1 => n2001, C2 => n107
                           , A => n2225, ZN => n2218);
   U3086 : OAI22_X1 port map( A1 => n11, A2 => n412, B1 => n467, B2 => n2003, 
                           ZN => n2225);
   U3087 : NAND4_X1 port map( A1 => n2226, A2 => n2227, A3 => n2228, A4 => 
                           n2229, ZN => n2207);
   U3088 : AOI221_X1 port map( B1 => n2008, B2 => n6108, C1 => n2009, C2 => 
                           n6140, A => n2230, ZN => n2229);
   U3089 : OAI222_X1 port map( A1 => n4892, A2 => n2011, B1 => n4860, B2 => 
                           n2012, C1 => n4828, C2 => n418, ZN => n2230);
   U3090 : AOI221_X1 port map( B1 => n2013, B2 => n6172, C1 => n2014, C2 => 
                           n6204, A => n2231, ZN => n2228);
   U3091 : OAI22_X1 port map( A1 => n5640, A2 => n2016, B1 => n5641, B2 => 
                           n2017, ZN => n2231);
   U3092 : AOI221_X1 port map( B1 => n1751, B2 => n6236, C1 => n2019, C2 => 
                           n6268, A => n2232, ZN => n2227);
   U3093 : OAI222_X1 port map( A1 => n4988, A2 => n2021, B1 => n4956, B2 => 
                           n2022, C1 => n4924, C2 => n419, ZN => n2232);
   U3094 : AOI221_X1 port map( B1 => n2023, B2 => n564, C1 => n2024, C2 => n108
                           , A => n2233, ZN => n2226);
   U3095 : OAI22_X1 port map( A1 => n12, A2 => n2026, B1 => n468, B2 => n2027, 
                           ZN => n2233);
   U3096 : NAND4_X1 port map( A1 => n2234, A2 => n2235, A3 => n2236, A4 => 
                           n2237, ZN => n2206);
   U3097 : AOI221_X1 port map( B1 => n2032, B2 => n5852, C1 => n2033, C2 => 
                           n5884, A => n2238, ZN => n2237);
   U3098 : OAI222_X1 port map( A1 => n4636, A2 => n2035, B1 => n4604, B2 => 
                           n2036, C1 => n4572, C2 => n1577, ZN => n2238);
   U3099 : AOI221_X1 port map( B1 => n2037, B2 => n5916, C1 => n2038, C2 => 
                           n5948, A => n2239, ZN => n2236);
   U3100 : OAI22_X1 port map( A1 => n4700, A2 => n2040, B1 => n4668, B2 => 
                           n2041, ZN => n2239);
   U3101 : AOI221_X1 port map( B1 => n1752, B2 => n5980, C1 => n2043, C2 => 
                           n6012, A => n2240, ZN => n2235);
   U3102 : OAI222_X1 port map( A1 => n4796, A2 => n411, B1 => n4764, B2 => 
                           n2045, C1 => n4732, C2 => n2046, ZN => n2240);
   U3103 : AOI221_X1 port map( B1 => n1749, B2 => n6044, C1 => n2048, C2 => 
                           n6076, A => n2241, ZN => n2234);
   U3104 : OAI22_X1 port map( A1 => n5638, A2 => n2050, B1 => n5639, B2 => 
                           n2051, ZN => n2241);
   U3105 : OAI21_X1 port map( B1 => n1951, B2 => n1518, A => ENABLE, ZN => 
                           n7662);
   U3106 : OAI222_X1 port map( A1 => n2242, A2 => n1948, B1 => n2243, B2 => 
                           n1950, C1 => n1951, C2 => n1455, ZN => n7661);
   U3107 : NOR4_X1 port map( A1 => n2244, A2 => n2245, A3 => n2246, A4 => n2247
                           , ZN => n2243);
   U3108 : NAND4_X1 port map( A1 => n2248, A2 => n2249, A3 => n2250, A4 => 
                           n2251, ZN => n2247);
   U3109 : AOI221_X1 port map( B1 => n1960, B2 => n6427, C1 => n1961, C2 => 
                           n6459, A => n2252, ZN => n2251);
   U3110 : OAI222_X1 port map( A1 => n5275, A2 => n1963, B1 => n5243, B2 => 
                           n1964, C1 => n5211, C2 => n1965, ZN => n2252);
   U3111 : AOI221_X1 port map( B1 => n1966, B2 => n6491, C1 => n1967, C2 => 
                           n6523, A => n2253, ZN => n2250);
   U3112 : OAI22_X1 port map( A1 => n5634, A2 => n1969, B1 => n5635, B2 => 
                           n1970, ZN => n2253);
   U3113 : AOI221_X1 port map( B1 => n1971, B2 => n6555, C1 => n1972, C2 => 
                           n6587, A => n2254, ZN => n2249);
   U3114 : OAI222_X1 port map( A1 => n5371, A2 => n1974, B1 => n5339, B2 => 
                           n1578, C1 => n5307, C2 => n1975, ZN => n2254);
   U3115 : AOI221_X1 port map( B1 => n1976, B2 => n6619, C1 => n1977, C2 => 
                           n6651, A => n2255, ZN => n2248);
   U3116 : OAI22_X1 port map( A1 => n5636, A2 => n1756, B1 => n5637, B2 => 
                           n1980, ZN => n2255);
   U3117 : NAND4_X1 port map( A1 => n2256, A2 => n2257, A3 => n2258, A4 => 
                           n2259, ZN => n2246);
   U3118 : AOI221_X1 port map( B1 => n1985, B2 => n6299, C1 => n1986, C2 => 
                           n6331, A => n2260, ZN => n2259);
   U3119 : OAI222_X1 port map( A1 => n5083, A2 => n1988, B1 => n5051, B2 => 
                           n1989, C1 => n5019, C2 => n416, ZN => n2260);
   U3120 : AOI221_X1 port map( B1 => n1990, B2 => n167, C1 => n1991, C2 => n527
                           , A => n2261, ZN => n2258);
   U3121 : OAI22_X1 port map( A1 => n71, A2 => n1993, B1 => n431, B2 => n1994, 
                           ZN => n2261);
   U3122 : AOI221_X1 port map( B1 => n1995, B2 => n6363, C1 => n1996, C2 => 
                           n6395, A => n2262, ZN => n2257);
   U3123 : OAI222_X1 port map( A1 => n5179, A2 => n1998, B1 => n5147, B2 => 
                           n1999, C1 => n5115, C2 => n417, ZN => n2262);
   U3124 : AOI221_X1 port map( B1 => n2000, B2 => n565, C1 => n2001, C2 => n109
                           , A => n2263, ZN => n2256);
   U3125 : OAI22_X1 port map( A1 => n13, A2 => n412, B1 => n469, B2 => n2003, 
                           ZN => n2263);
   U3126 : NAND4_X1 port map( A1 => n2264, A2 => n2265, A3 => n2266, A4 => 
                           n2267, ZN => n2245);
   U3127 : AOI221_X1 port map( B1 => n2008, B2 => n6107, C1 => n2009, C2 => 
                           n6139, A => n2268, ZN => n2267);
   U3128 : OAI222_X1 port map( A1 => n4891, A2 => n2011, B1 => n4859, B2 => 
                           n2012, C1 => n4827, C2 => n418, ZN => n2268);
   U3129 : AOI221_X1 port map( B1 => n2013, B2 => n6171, C1 => n2014, C2 => 
                           n6203, A => n2269, ZN => n2266);
   U3130 : OAI22_X1 port map( A1 => n5630, A2 => n2016, B1 => n5631, B2 => 
                           n2017, ZN => n2269);
   U3131 : AOI221_X1 port map( B1 => n1751, B2 => n6235, C1 => n2019, C2 => 
                           n6267, A => n2270, ZN => n2265);
   U3132 : OAI222_X1 port map( A1 => n4987, A2 => n2021, B1 => n4955, B2 => 
                           n2022, C1 => n4923, C2 => n419, ZN => n2270);
   U3133 : AOI221_X1 port map( B1 => n2023, B2 => n566, C1 => n2024, C2 => n110
                           , A => n2271, ZN => n2264);
   U3134 : OAI22_X1 port map( A1 => n14, A2 => n2026, B1 => n470, B2 => n2027, 
                           ZN => n2271);
   U3135 : NAND4_X1 port map( A1 => n2272, A2 => n2273, A3 => n2274, A4 => 
                           n2275, ZN => n2244);
   U3136 : AOI221_X1 port map( B1 => n2032, B2 => n5851, C1 => n2033, C2 => 
                           n5883, A => n2276, ZN => n2275);
   U3137 : OAI222_X1 port map( A1 => n4635, A2 => n2035, B1 => n4603, B2 => 
                           n2036, C1 => n4571, C2 => n1577, ZN => n2276);
   U3138 : AOI221_X1 port map( B1 => n2037, B2 => n5915, C1 => n2038, C2 => 
                           n5947, A => n2277, ZN => n2274);
   U3139 : OAI22_X1 port map( A1 => n4699, A2 => n2040, B1 => n4667, B2 => 
                           n2041, ZN => n2277);
   U3140 : AOI221_X1 port map( B1 => n1752, B2 => n5979, C1 => n2043, C2 => 
                           n6011, A => n2278, ZN => n2273);
   U3141 : OAI222_X1 port map( A1 => n4795, A2 => n411, B1 => n4763, B2 => 
                           n2045, C1 => n4731, C2 => n2046, ZN => n2278);
   U3142 : AOI221_X1 port map( B1 => n1749, B2 => n6043, C1 => n2048, C2 => 
                           n6075, A => n2279, ZN => n2272);
   U3143 : OAI22_X1 port map( A1 => n5628, A2 => n2050, B1 => n5629, B2 => 
                           n2051, ZN => n2279);
   U3144 : OAI21_X1 port map( B1 => n1951, B2 => n1519, A => ENABLE, ZN => 
                           n7660);
   U3145 : OAI222_X1 port map( A1 => n2280, A2 => n1948, B1 => n2281, B2 => 
                           n1950, C1 => n1951, C2 => n1456, ZN => n7659);
   U3146 : NOR4_X1 port map( A1 => n2282, A2 => n2283, A3 => n2284, A4 => n2285
                           , ZN => n2281);
   U3147 : NAND4_X1 port map( A1 => n2286, A2 => n2287, A3 => n2288, A4 => 
                           n2289, ZN => n2285);
   U3148 : AOI221_X1 port map( B1 => n1960, B2 => n6426, C1 => n1961, C2 => 
                           n6458, A => n2290, ZN => n2289);
   U3149 : OAI222_X1 port map( A1 => n5274, A2 => n1963, B1 => n5242, B2 => 
                           n1964, C1 => n5210, C2 => n1965, ZN => n2290);
   U3150 : AOI221_X1 port map( B1 => n1966, B2 => n6490, C1 => n1967, C2 => 
                           n6522, A => n2291, ZN => n2288);
   U3151 : OAI22_X1 port map( A1 => n5624, A2 => n1969, B1 => n5625, B2 => 
                           n1970, ZN => n2291);
   U3152 : AOI221_X1 port map( B1 => n1971, B2 => n6554, C1 => n1972, C2 => 
                           n6586, A => n2292, ZN => n2287);
   U3153 : OAI222_X1 port map( A1 => n5370, A2 => n1974, B1 => n5338, B2 => 
                           n1578, C1 => n5306, C2 => n1975, ZN => n2292);
   U3154 : AOI221_X1 port map( B1 => n1976, B2 => n6618, C1 => n1977, C2 => 
                           n6650, A => n2293, ZN => n2286);
   U3155 : OAI22_X1 port map( A1 => n5626, A2 => n1756, B1 => n5627, B2 => 
                           n1980, ZN => n2293);
   U3156 : NAND4_X1 port map( A1 => n2294, A2 => n2295, A3 => n2296, A4 => 
                           n2297, ZN => n2284);
   U3157 : AOI221_X1 port map( B1 => n1985, B2 => n6298, C1 => n1986, C2 => 
                           n6330, A => n2298, ZN => n2297);
   U3158 : OAI222_X1 port map( A1 => n5082, A2 => n1988, B1 => n5050, B2 => 
                           n1989, C1 => n5018, C2 => n416, ZN => n2298);
   U3159 : AOI221_X1 port map( B1 => n1990, B2 => n168, C1 => n1991, C2 => n528
                           , A => n2299, ZN => n2296);
   U3160 : OAI22_X1 port map( A1 => n72, A2 => n1993, B1 => n432, B2 => n1994, 
                           ZN => n2299);
   U3161 : AOI221_X1 port map( B1 => n1995, B2 => n6362, C1 => n1996, C2 => 
                           n6394, A => n2300, ZN => n2295);
   U3162 : OAI222_X1 port map( A1 => n5178, A2 => n1998, B1 => n5146, B2 => 
                           n1999, C1 => n5114, C2 => n417, ZN => n2300);
   U3163 : AOI221_X1 port map( B1 => n2000, B2 => n567, C1 => n2001, C2 => n111
                           , A => n2301, ZN => n2294);
   U3164 : OAI22_X1 port map( A1 => n15, A2 => n412, B1 => n471, B2 => n2003, 
                           ZN => n2301);
   U3165 : NAND4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2304, A4 => 
                           n2305, ZN => n2283);
   U3166 : AOI221_X1 port map( B1 => n2008, B2 => n6106, C1 => n2009, C2 => 
                           n6138, A => n2306, ZN => n2305);
   U3167 : OAI222_X1 port map( A1 => n4890, A2 => n2011, B1 => n4858, B2 => 
                           n2012, C1 => n4826, C2 => n418, ZN => n2306);
   U3168 : AOI221_X1 port map( B1 => n2013, B2 => n6170, C1 => n2014, C2 => 
                           n6202, A => n2307, ZN => n2304);
   U3169 : OAI22_X1 port map( A1 => n5620, A2 => n2016, B1 => n5621, B2 => 
                           n2017, ZN => n2307);
   U3170 : AOI221_X1 port map( B1 => n2018, B2 => n6234, C1 => n2019, C2 => 
                           n6266, A => n2308, ZN => n2303);
   U3171 : OAI222_X1 port map( A1 => n4986, A2 => n2021, B1 => n4954, B2 => 
                           n2022, C1 => n4922, C2 => n419, ZN => n2308);
   U3172 : AOI221_X1 port map( B1 => n2023, B2 => n568, C1 => n2024, C2 => n112
                           , A => n2309, ZN => n2302);
   U3173 : OAI22_X1 port map( A1 => n16, A2 => n2026, B1 => n472, B2 => n2027, 
                           ZN => n2309);
   U3174 : NAND4_X1 port map( A1 => n2310, A2 => n2311, A3 => n2312, A4 => 
                           n2313, ZN => n2282);
   U3175 : AOI221_X1 port map( B1 => n2032, B2 => n5850, C1 => n2033, C2 => 
                           n5882, A => n2314, ZN => n2313);
   U3176 : OAI222_X1 port map( A1 => n4634, A2 => n2035, B1 => n4602, B2 => 
                           n2036, C1 => n4570, C2 => n1577, ZN => n2314);
   U3177 : AOI221_X1 port map( B1 => n2037, B2 => n5914, C1 => n2038, C2 => 
                           n5946, A => n2315, ZN => n2312);
   U3178 : OAI22_X1 port map( A1 => n4698, A2 => n2040, B1 => n4666, B2 => 
                           n2041, ZN => n2315);
   U3179 : AOI221_X1 port map( B1 => n2042, B2 => n5978, C1 => n2043, C2 => 
                           n6010, A => n2316, ZN => n2311);
   U3180 : OAI222_X1 port map( A1 => n4794, A2 => n411, B1 => n4762, B2 => 
                           n2045, C1 => n4730, C2 => n2046, ZN => n2316);
   U3181 : AOI221_X1 port map( B1 => n2047, B2 => n6042, C1 => n2048, C2 => 
                           n6074, A => n2317, ZN => n2310);
   U3182 : OAI22_X1 port map( A1 => n5618, A2 => n2050, B1 => n5619, B2 => 
                           n2051, ZN => n2317);
   U3183 : OAI21_X1 port map( B1 => n1951, B2 => n1520, A => ENABLE, ZN => 
                           n7658);
   U3184 : OAI222_X1 port map( A1 => n2318, A2 => n1948, B1 => n2319, B2 => 
                           n1950, C1 => n1951, C2 => n1457, ZN => n7657);
   U3185 : NOR4_X1 port map( A1 => n2320, A2 => n2321, A3 => n2322, A4 => n2323
                           , ZN => n2319);
   U3186 : NAND4_X1 port map( A1 => n2324, A2 => n2325, A3 => n2326, A4 => 
                           n2327, ZN => n2323);
   U3187 : AOI221_X1 port map( B1 => n1960, B2 => n6425, C1 => n1961, C2 => 
                           n6457, A => n2328, ZN => n2327);
   U3188 : OAI222_X1 port map( A1 => n5273, A2 => n1963, B1 => n5241, B2 => 
                           n1964, C1 => n5209, C2 => n1965, ZN => n2328);
   U3189 : AOI221_X1 port map( B1 => n1966, B2 => n6489, C1 => n1967, C2 => 
                           n6521, A => n2329, ZN => n2326);
   U3190 : OAI22_X1 port map( A1 => n5614, A2 => n1969, B1 => n5615, B2 => 
                           n1970, ZN => n2329);
   U3191 : AOI221_X1 port map( B1 => n1971, B2 => n6553, C1 => n1972, C2 => 
                           n6585, A => n2330, ZN => n2325);
   U3192 : OAI222_X1 port map( A1 => n5369, A2 => n1974, B1 => n5337, B2 => 
                           n1578, C1 => n5305, C2 => n1975, ZN => n2330);
   U3193 : AOI221_X1 port map( B1 => n1976, B2 => n6617, C1 => n1977, C2 => 
                           n6649, A => n2331, ZN => n2324);
   U3194 : OAI22_X1 port map( A1 => n5616, A2 => n1756, B1 => n5617, B2 => 
                           n1980, ZN => n2331);
   U3195 : NAND4_X1 port map( A1 => n2332, A2 => n2333, A3 => n2334, A4 => 
                           n2335, ZN => n2322);
   U3196 : AOI221_X1 port map( B1 => n1985, B2 => n6297, C1 => n1986, C2 => 
                           n6329, A => n2336, ZN => n2335);
   U3197 : OAI222_X1 port map( A1 => n5081, A2 => n1988, B1 => n5049, B2 => 
                           n1989, C1 => n5017, C2 => n416, ZN => n2336);
   U3198 : AOI221_X1 port map( B1 => n1990, B2 => n169, C1 => n1991, C2 => n529
                           , A => n2337, ZN => n2334);
   U3199 : OAI22_X1 port map( A1 => n73, A2 => n1993, B1 => n433, B2 => n1994, 
                           ZN => n2337);
   U3200 : AOI221_X1 port map( B1 => n1995, B2 => n6361, C1 => n1996, C2 => 
                           n6393, A => n2338, ZN => n2333);
   U3201 : OAI222_X1 port map( A1 => n5177, A2 => n1998, B1 => n5145, B2 => 
                           n1999, C1 => n5113, C2 => n417, ZN => n2338);
   U3202 : AOI221_X1 port map( B1 => n2000, B2 => n569, C1 => n2001, C2 => n113
                           , A => n2339, ZN => n2332);
   U3203 : OAI22_X1 port map( A1 => n17, A2 => n412, B1 => n473, B2 => n2003, 
                           ZN => n2339);
   U3204 : NAND4_X1 port map( A1 => n2340, A2 => n2341, A3 => n2342, A4 => 
                           n2343, ZN => n2321);
   U3205 : AOI221_X1 port map( B1 => n2008, B2 => n6105, C1 => n2009, C2 => 
                           n6137, A => n2344, ZN => n2343);
   U3206 : OAI222_X1 port map( A1 => n4889, A2 => n2011, B1 => n4857, B2 => 
                           n2012, C1 => n4825, C2 => n418, ZN => n2344);
   U3207 : AOI221_X1 port map( B1 => n2013, B2 => n6169, C1 => n2014, C2 => 
                           n6201, A => n2345, ZN => n2342);
   U3208 : OAI22_X1 port map( A1 => n5610, A2 => n2016, B1 => n5611, B2 => 
                           n2017, ZN => n2345);
   U3209 : AOI221_X1 port map( B1 => n2018, B2 => n6233, C1 => n2019, C2 => 
                           n6265, A => n2346, ZN => n2341);
   U3210 : OAI222_X1 port map( A1 => n4985, A2 => n2021, B1 => n4953, B2 => 
                           n2022, C1 => n4921, C2 => n419, ZN => n2346);
   U3211 : AOI221_X1 port map( B1 => n2023, B2 => n570, C1 => n2024, C2 => n114
                           , A => n2347, ZN => n2340);
   U3212 : OAI22_X1 port map( A1 => n18, A2 => n2026, B1 => n474, B2 => n2027, 
                           ZN => n2347);
   U3213 : NAND4_X1 port map( A1 => n2348, A2 => n2349, A3 => n2350, A4 => 
                           n2351, ZN => n2320);
   U3214 : AOI221_X1 port map( B1 => n2032, B2 => n5849, C1 => n2033, C2 => 
                           n5881, A => n2352, ZN => n2351);
   U3215 : OAI222_X1 port map( A1 => n4633, A2 => n2035, B1 => n4601, B2 => 
                           n2036, C1 => n4569, C2 => n1577, ZN => n2352);
   U3216 : AOI221_X1 port map( B1 => n2037, B2 => n5913, C1 => n2038, C2 => 
                           n5945, A => n2353, ZN => n2350);
   U3217 : OAI22_X1 port map( A1 => n4697, A2 => n2040, B1 => n4665, B2 => 
                           n2041, ZN => n2353);
   U3218 : AOI221_X1 port map( B1 => n2042, B2 => n5977, C1 => n2043, C2 => 
                           n6009, A => n2354, ZN => n2349);
   U3219 : OAI222_X1 port map( A1 => n4793, A2 => n411, B1 => n4761, B2 => 
                           n2045, C1 => n4729, C2 => n2046, ZN => n2354);
   U3220 : AOI221_X1 port map( B1 => n2047, B2 => n6041, C1 => n2048, C2 => 
                           n6073, A => n2355, ZN => n2348);
   U3221 : OAI22_X1 port map( A1 => n5608, A2 => n2050, B1 => n5609, B2 => 
                           n2051, ZN => n2355);
   U3222 : OAI21_X1 port map( B1 => n1951, B2 => n1521, A => ENABLE, ZN => 
                           n7656);
   U3223 : OAI222_X1 port map( A1 => n2356, A2 => n1948, B1 => n2357, B2 => 
                           n1950, C1 => n1951, C2 => n1458, ZN => n7655);
   U3224 : NOR4_X1 port map( A1 => n2358, A2 => n2359, A3 => n2360, A4 => n2361
                           , ZN => n2357);
   U3225 : NAND4_X1 port map( A1 => n2362, A2 => n2363, A3 => n2364, A4 => 
                           n2365, ZN => n2361);
   U3226 : AOI221_X1 port map( B1 => n1960, B2 => n6424, C1 => n1961, C2 => 
                           n6456, A => n2366, ZN => n2365);
   U3227 : OAI222_X1 port map( A1 => n5272, A2 => n1963, B1 => n5240, B2 => 
                           n1964, C1 => n5208, C2 => n1965, ZN => n2366);
   U3228 : AOI221_X1 port map( B1 => n1966, B2 => n6488, C1 => n1967, C2 => 
                           n6520, A => n2367, ZN => n2364);
   U3229 : OAI22_X1 port map( A1 => n5604, A2 => n1969, B1 => n5605, B2 => 
                           n1970, ZN => n2367);
   U3230 : AOI221_X1 port map( B1 => n1971, B2 => n6552, C1 => n1972, C2 => 
                           n6584, A => n2368, ZN => n2363);
   U3231 : OAI222_X1 port map( A1 => n5368, A2 => n1974, B1 => n5336, B2 => 
                           n1578, C1 => n5304, C2 => n1975, ZN => n2368);
   U3232 : AOI221_X1 port map( B1 => n1976, B2 => n6616, C1 => n1977, C2 => 
                           n6648, A => n2369, ZN => n2362);
   U3233 : OAI22_X1 port map( A1 => n5606, A2 => n1756, B1 => n5607, B2 => 
                           n1980, ZN => n2369);
   U3234 : NAND4_X1 port map( A1 => n2370, A2 => n2371, A3 => n2372, A4 => 
                           n2373, ZN => n2360);
   U3235 : AOI221_X1 port map( B1 => n1985, B2 => n6296, C1 => n1986, C2 => 
                           n6328, A => n2374, ZN => n2373);
   U3236 : OAI222_X1 port map( A1 => n5080, A2 => n1988, B1 => n5048, B2 => 
                           n1989, C1 => n5016, C2 => n416, ZN => n2374);
   U3237 : AOI221_X1 port map( B1 => n1990, B2 => n170, C1 => n1991, C2 => n530
                           , A => n2375, ZN => n2372);
   U3238 : OAI22_X1 port map( A1 => n74, A2 => n1993, B1 => n434, B2 => n1994, 
                           ZN => n2375);
   U3239 : AOI221_X1 port map( B1 => n1995, B2 => n6360, C1 => n1996, C2 => 
                           n6392, A => n2376, ZN => n2371);
   U3240 : OAI222_X1 port map( A1 => n5176, A2 => n1998, B1 => n5144, B2 => 
                           n1999, C1 => n5112, C2 => n417, ZN => n2376);
   U3241 : AOI221_X1 port map( B1 => n2000, B2 => n571, C1 => n2001, C2 => n115
                           , A => n2377, ZN => n2370);
   U3242 : OAI22_X1 port map( A1 => n19, A2 => n412, B1 => n475, B2 => n2003, 
                           ZN => n2377);
   U3243 : NAND4_X1 port map( A1 => n2378, A2 => n2379, A3 => n2380, A4 => 
                           n2381, ZN => n2359);
   U3244 : AOI221_X1 port map( B1 => n2008, B2 => n6104, C1 => n2009, C2 => 
                           n6136, A => n2382, ZN => n2381);
   U3245 : OAI222_X1 port map( A1 => n4888, A2 => n2011, B1 => n4856, B2 => 
                           n2012, C1 => n4824, C2 => n418, ZN => n2382);
   U3246 : AOI221_X1 port map( B1 => n2013, B2 => n6168, C1 => n2014, C2 => 
                           n6200, A => n2383, ZN => n2380);
   U3247 : OAI22_X1 port map( A1 => n5600, A2 => n2016, B1 => n5601, B2 => 
                           n2017, ZN => n2383);
   U3248 : AOI221_X1 port map( B1 => n2018, B2 => n6232, C1 => n2019, C2 => 
                           n6264, A => n2384, ZN => n2379);
   U3249 : OAI222_X1 port map( A1 => n4984, A2 => n2021, B1 => n4952, B2 => 
                           n2022, C1 => n4920, C2 => n419, ZN => n2384);
   U3250 : AOI221_X1 port map( B1 => n2023, B2 => n572, C1 => n2024, C2 => n116
                           , A => n2385, ZN => n2378);
   U3251 : OAI22_X1 port map( A1 => n20, A2 => n2026, B1 => n476, B2 => n2027, 
                           ZN => n2385);
   U3252 : NAND4_X1 port map( A1 => n2386, A2 => n2387, A3 => n2388, A4 => 
                           n2389, ZN => n2358);
   U3253 : AOI221_X1 port map( B1 => n2032, B2 => n5848, C1 => n2033, C2 => 
                           n5880, A => n2390, ZN => n2389);
   U3254 : OAI222_X1 port map( A1 => n4632, A2 => n2035, B1 => n4600, B2 => 
                           n2036, C1 => n4568, C2 => n1577, ZN => n2390);
   U3255 : AOI221_X1 port map( B1 => n2037, B2 => n5912, C1 => n2038, C2 => 
                           n5944, A => n2391, ZN => n2388);
   U3256 : OAI22_X1 port map( A1 => n4696, A2 => n2040, B1 => n4664, B2 => 
                           n2041, ZN => n2391);
   U3257 : AOI221_X1 port map( B1 => n2042, B2 => n5976, C1 => n2043, C2 => 
                           n6008, A => n2392, ZN => n2387);
   U3258 : OAI222_X1 port map( A1 => n4792, A2 => n411, B1 => n4760, B2 => 
                           n2045, C1 => n4728, C2 => n2046, ZN => n2392);
   U3259 : AOI221_X1 port map( B1 => n2047, B2 => n6040, C1 => n2048, C2 => 
                           n6072, A => n2393, ZN => n2386);
   U3260 : OAI22_X1 port map( A1 => n5598, A2 => n2050, B1 => n5599, B2 => 
                           n2051, ZN => n2393);
   U3261 : OAI21_X1 port map( B1 => n1951, B2 => n1522, A => ENABLE, ZN => 
                           n7654);
   U3262 : OAI222_X1 port map( A1 => n2394, A2 => n1948, B1 => n2395, B2 => 
                           n1950, C1 => n1951, C2 => n1459, ZN => n7653);
   U3263 : NOR4_X1 port map( A1 => n2396, A2 => n2397, A3 => n2398, A4 => n2399
                           , ZN => n2395);
   U3264 : NAND4_X1 port map( A1 => n2400, A2 => n2401, A3 => n2402, A4 => 
                           n2403, ZN => n2399);
   U3265 : AOI221_X1 port map( B1 => n1960, B2 => n6423, C1 => n1961, C2 => 
                           n6455, A => n2404, ZN => n2403);
   U3266 : OAI222_X1 port map( A1 => n5271, A2 => n1963, B1 => n5239, B2 => 
                           n1964, C1 => n5207, C2 => n1965, ZN => n2404);
   U3267 : AOI221_X1 port map( B1 => n1966, B2 => n6487, C1 => n1967, C2 => 
                           n6519, A => n2405, ZN => n2402);
   U3268 : OAI22_X1 port map( A1 => n5594, A2 => n1969, B1 => n5595, B2 => 
                           n1970, ZN => n2405);
   U3269 : AOI221_X1 port map( B1 => n1971, B2 => n6551, C1 => n1972, C2 => 
                           n6583, A => n2406, ZN => n2401);
   U3270 : OAI222_X1 port map( A1 => n5367, A2 => n1974, B1 => n5335, B2 => 
                           n1578, C1 => n5303, C2 => n1975, ZN => n2406);
   U3271 : AOI221_X1 port map( B1 => n1976, B2 => n6615, C1 => n1977, C2 => 
                           n6647, A => n2407, ZN => n2400);
   U3272 : OAI22_X1 port map( A1 => n5596, A2 => n1756, B1 => n5597, B2 => 
                           n1980, ZN => n2407);
   U3273 : NAND4_X1 port map( A1 => n2408, A2 => n2409, A3 => n2410, A4 => 
                           n2411, ZN => n2398);
   U3274 : AOI221_X1 port map( B1 => n1985, B2 => n6295, C1 => n1986, C2 => 
                           n6327, A => n2412, ZN => n2411);
   U3275 : OAI222_X1 port map( A1 => n5079, A2 => n1988, B1 => n5047, B2 => 
                           n1989, C1 => n5015, C2 => n416, ZN => n2412);
   U3276 : AOI221_X1 port map( B1 => n1990, B2 => n171, C1 => n1991, C2 => n531
                           , A => n2413, ZN => n2410);
   U3277 : OAI22_X1 port map( A1 => n75, A2 => n1993, B1 => n435, B2 => n1994, 
                           ZN => n2413);
   U3278 : AOI221_X1 port map( B1 => n1995, B2 => n6359, C1 => n1996, C2 => 
                           n6391, A => n2414, ZN => n2409);
   U3279 : OAI222_X1 port map( A1 => n5175, A2 => n1998, B1 => n5143, B2 => 
                           n1999, C1 => n5111, C2 => n417, ZN => n2414);
   U3280 : AOI221_X1 port map( B1 => n2000, B2 => n573, C1 => n2001, C2 => n117
                           , A => n2415, ZN => n2408);
   U3281 : OAI22_X1 port map( A1 => n21, A2 => n412, B1 => n477, B2 => n2003, 
                           ZN => n2415);
   U3282 : NAND4_X1 port map( A1 => n2416, A2 => n2417, A3 => n2418, A4 => 
                           n2419, ZN => n2397);
   U3283 : AOI221_X1 port map( B1 => n2008, B2 => n6103, C1 => n2009, C2 => 
                           n6135, A => n2420, ZN => n2419);
   U3284 : OAI222_X1 port map( A1 => n4887, A2 => n2011, B1 => n4855, B2 => 
                           n2012, C1 => n4823, C2 => n418, ZN => n2420);
   U3285 : AOI221_X1 port map( B1 => n2013, B2 => n6167, C1 => n2014, C2 => 
                           n6199, A => n2421, ZN => n2418);
   U3286 : OAI22_X1 port map( A1 => n5590, A2 => n2016, B1 => n5591, B2 => 
                           n2017, ZN => n2421);
   U3287 : AOI221_X1 port map( B1 => n2018, B2 => n6231, C1 => n2019, C2 => 
                           n6263, A => n2422, ZN => n2417);
   U3288 : OAI222_X1 port map( A1 => n4983, A2 => n2021, B1 => n4951, B2 => 
                           n2022, C1 => n4919, C2 => n419, ZN => n2422);
   U3289 : AOI221_X1 port map( B1 => n2023, B2 => n574, C1 => n2024, C2 => n118
                           , A => n2423, ZN => n2416);
   U3290 : OAI22_X1 port map( A1 => n22, A2 => n2026, B1 => n478, B2 => n2027, 
                           ZN => n2423);
   U3291 : NAND4_X1 port map( A1 => n2424, A2 => n2425, A3 => n2426, A4 => 
                           n2427, ZN => n2396);
   U3292 : AOI221_X1 port map( B1 => n2032, B2 => n5847, C1 => n2033, C2 => 
                           n5879, A => n2428, ZN => n2427);
   U3293 : OAI222_X1 port map( A1 => n4631, A2 => n2035, B1 => n4599, B2 => 
                           n2036, C1 => n4567, C2 => n1577, ZN => n2428);
   U3294 : AOI221_X1 port map( B1 => n2037, B2 => n5911, C1 => n2038, C2 => 
                           n5943, A => n2429, ZN => n2426);
   U3295 : OAI22_X1 port map( A1 => n4695, A2 => n2040, B1 => n4663, B2 => 
                           n2041, ZN => n2429);
   U3296 : AOI221_X1 port map( B1 => n2042, B2 => n5975, C1 => n2043, C2 => 
                           n6007, A => n2430, ZN => n2425);
   U3297 : OAI222_X1 port map( A1 => n4791, A2 => n411, B1 => n4759, B2 => 
                           n2045, C1 => n4727, C2 => n2046, ZN => n2430);
   U3298 : AOI221_X1 port map( B1 => n2047, B2 => n6039, C1 => n2048, C2 => 
                           n6071, A => n2431, ZN => n2424);
   U3299 : OAI22_X1 port map( A1 => n5588, A2 => n2050, B1 => n5589, B2 => 
                           n2051, ZN => n2431);
   U3300 : OAI21_X1 port map( B1 => n1951, B2 => n1523, A => ENABLE, ZN => 
                           n7652);
   U3301 : OAI222_X1 port map( A1 => n2432, A2 => n1948, B1 => n2433, B2 => 
                           n1950, C1 => n1951, C2 => n1460, ZN => n7651);
   U3302 : NOR4_X1 port map( A1 => n2434, A2 => n2435, A3 => n2436, A4 => n2437
                           , ZN => n2433);
   U3303 : NAND4_X1 port map( A1 => n2438, A2 => n2439, A3 => n2440, A4 => 
                           n2441, ZN => n2437);
   U3304 : AOI221_X1 port map( B1 => n1960, B2 => n6422, C1 => n1961, C2 => 
                           n6454, A => n2442, ZN => n2441);
   U3305 : OAI222_X1 port map( A1 => n5270, A2 => n1963, B1 => n5238, B2 => 
                           n1964, C1 => n5206, C2 => n1965, ZN => n2442);
   U3306 : AOI221_X1 port map( B1 => n1966, B2 => n6486, C1 => n1967, C2 => 
                           n6518, A => n2443, ZN => n2440);
   U3307 : OAI22_X1 port map( A1 => n5584, A2 => n1969, B1 => n5585, B2 => 
                           n1970, ZN => n2443);
   U3308 : AOI221_X1 port map( B1 => n1971, B2 => n6550, C1 => n1972, C2 => 
                           n6582, A => n2444, ZN => n2439);
   U3309 : OAI222_X1 port map( A1 => n5366, A2 => n1974, B1 => n5334, B2 => 
                           n1578, C1 => n5302, C2 => n1975, ZN => n2444);
   U3310 : AOI221_X1 port map( B1 => n1976, B2 => n6614, C1 => n1977, C2 => 
                           n6646, A => n2445, ZN => n2438);
   U3311 : OAI22_X1 port map( A1 => n5586, A2 => n1756, B1 => n5587, B2 => 
                           n1980, ZN => n2445);
   U3312 : NAND4_X1 port map( A1 => n2446, A2 => n2447, A3 => n2448, A4 => 
                           n2449, ZN => n2436);
   U3313 : AOI221_X1 port map( B1 => n1985, B2 => n6294, C1 => n1986, C2 => 
                           n6326, A => n2450, ZN => n2449);
   U3314 : OAI222_X1 port map( A1 => n5078, A2 => n1988, B1 => n5046, B2 => 
                           n1989, C1 => n5014, C2 => n416, ZN => n2450);
   U3315 : AOI221_X1 port map( B1 => n1990, B2 => n172, C1 => n1991, C2 => n532
                           , A => n2451, ZN => n2448);
   U3316 : OAI22_X1 port map( A1 => n76, A2 => n1993, B1 => n436, B2 => n1994, 
                           ZN => n2451);
   U3317 : AOI221_X1 port map( B1 => n1995, B2 => n6358, C1 => n1996, C2 => 
                           n6390, A => n2452, ZN => n2447);
   U3318 : OAI222_X1 port map( A1 => n5174, A2 => n1998, B1 => n5142, B2 => 
                           n1999, C1 => n5110, C2 => n417, ZN => n2452);
   U3319 : AOI221_X1 port map( B1 => n2000, B2 => n575, C1 => n2001, C2 => n119
                           , A => n2453, ZN => n2446);
   U3320 : OAI22_X1 port map( A1 => n23, A2 => n412, B1 => n479, B2 => n2003, 
                           ZN => n2453);
   U3321 : NAND4_X1 port map( A1 => n2454, A2 => n2455, A3 => n2456, A4 => 
                           n2457, ZN => n2435);
   U3322 : AOI221_X1 port map( B1 => n2008, B2 => n6102, C1 => n2009, C2 => 
                           n6134, A => n2458, ZN => n2457);
   U3323 : OAI222_X1 port map( A1 => n4886, A2 => n2011, B1 => n4854, B2 => 
                           n2012, C1 => n4822, C2 => n418, ZN => n2458);
   U3324 : AOI221_X1 port map( B1 => n2013, B2 => n6166, C1 => n2014, C2 => 
                           n6198, A => n2459, ZN => n2456);
   U3325 : OAI22_X1 port map( A1 => n5580, A2 => n2016, B1 => n5581, B2 => 
                           n2017, ZN => n2459);
   U3326 : AOI221_X1 port map( B1 => n2018, B2 => n6230, C1 => n2019, C2 => 
                           n6262, A => n2460, ZN => n2455);
   U3327 : OAI222_X1 port map( A1 => n4982, A2 => n2021, B1 => n4950, B2 => 
                           n2022, C1 => n4918, C2 => n419, ZN => n2460);
   U3328 : AOI221_X1 port map( B1 => n2023, B2 => n576, C1 => n2024, C2 => n120
                           , A => n2461, ZN => n2454);
   U3329 : OAI22_X1 port map( A1 => n24, A2 => n2026, B1 => n480, B2 => n2027, 
                           ZN => n2461);
   U3330 : NAND4_X1 port map( A1 => n2462, A2 => n2463, A3 => n2464, A4 => 
                           n2465, ZN => n2434);
   U3331 : AOI221_X1 port map( B1 => n2032, B2 => n5846, C1 => n2033, C2 => 
                           n5878, A => n2466, ZN => n2465);
   U3332 : OAI222_X1 port map( A1 => n4630, A2 => n2035, B1 => n4598, B2 => 
                           n2036, C1 => n4566, C2 => n1577, ZN => n2466);
   U3333 : AOI221_X1 port map( B1 => n2037, B2 => n5910, C1 => n2038, C2 => 
                           n5942, A => n2467, ZN => n2464);
   U3334 : OAI22_X1 port map( A1 => n4694, A2 => n2040, B1 => n4662, B2 => 
                           n2041, ZN => n2467);
   U3335 : AOI221_X1 port map( B1 => n2042, B2 => n5974, C1 => n2043, C2 => 
                           n6006, A => n2468, ZN => n2463);
   U3336 : OAI222_X1 port map( A1 => n4790, A2 => n411, B1 => n4758, B2 => 
                           n2045, C1 => n4726, C2 => n2046, ZN => n2468);
   U3337 : AOI221_X1 port map( B1 => n2047, B2 => n6038, C1 => n2048, C2 => 
                           n6070, A => n2469, ZN => n2462);
   U3338 : OAI22_X1 port map( A1 => n5578, A2 => n2050, B1 => n5579, B2 => 
                           n2051, ZN => n2469);
   U3339 : OAI21_X1 port map( B1 => n1951, B2 => n1524, A => ENABLE, ZN => 
                           n7650);
   U3340 : OAI222_X1 port map( A1 => n2470, A2 => n1948, B1 => n2471, B2 => 
                           n1950, C1 => n1951, C2 => n1461, ZN => n7649);
   U3341 : NOR4_X1 port map( A1 => n2472, A2 => n2473, A3 => n2474, A4 => n2475
                           , ZN => n2471);
   U3342 : NAND4_X1 port map( A1 => n2476, A2 => n2477, A3 => n2478, A4 => 
                           n2479, ZN => n2475);
   U3343 : AOI221_X1 port map( B1 => n1960, B2 => n6421, C1 => n1961, C2 => 
                           n6453, A => n2480, ZN => n2479);
   U3344 : OAI222_X1 port map( A1 => n5269, A2 => n1963, B1 => n5237, B2 => 
                           n1964, C1 => n5205, C2 => n1965, ZN => n2480);
   U3345 : AOI221_X1 port map( B1 => n1966, B2 => n6485, C1 => n1967, C2 => 
                           n6517, A => n2481, ZN => n2478);
   U3346 : OAI22_X1 port map( A1 => n5574, A2 => n1969, B1 => n5575, B2 => 
                           n1970, ZN => n2481);
   U3347 : AOI221_X1 port map( B1 => n1971, B2 => n6549, C1 => n1972, C2 => 
                           n6581, A => n2482, ZN => n2477);
   U3348 : OAI222_X1 port map( A1 => n5365, A2 => n1974, B1 => n5333, B2 => 
                           n1578, C1 => n5301, C2 => n1975, ZN => n2482);
   U3349 : AOI221_X1 port map( B1 => n1976, B2 => n6613, C1 => n1977, C2 => 
                           n6645, A => n2483, ZN => n2476);
   U3350 : OAI22_X1 port map( A1 => n5576, A2 => n1756, B1 => n5577, B2 => 
                           n1980, ZN => n2483);
   U3351 : NAND4_X1 port map( A1 => n2484, A2 => n2485, A3 => n2486, A4 => 
                           n2487, ZN => n2474);
   U3352 : AOI221_X1 port map( B1 => n1985, B2 => n6293, C1 => n1986, C2 => 
                           n6325, A => n2488, ZN => n2487);
   U3353 : OAI222_X1 port map( A1 => n5077, A2 => n1988, B1 => n5045, B2 => 
                           n1989, C1 => n5013, C2 => n416, ZN => n2488);
   U3354 : AOI221_X1 port map( B1 => n1990, B2 => n173, C1 => n1991, C2 => n533
                           , A => n2489, ZN => n2486);
   U3355 : OAI22_X1 port map( A1 => n77, A2 => n1993, B1 => n437, B2 => n1994, 
                           ZN => n2489);
   U3356 : AOI221_X1 port map( B1 => n1995, B2 => n6357, C1 => n1996, C2 => 
                           n6389, A => n2490, ZN => n2485);
   U3357 : OAI222_X1 port map( A1 => n5173, A2 => n1998, B1 => n5141, B2 => 
                           n1999, C1 => n5109, C2 => n417, ZN => n2490);
   U3358 : AOI221_X1 port map( B1 => n2000, B2 => n577, C1 => n2001, C2 => n121
                           , A => n2491, ZN => n2484);
   U3359 : OAI22_X1 port map( A1 => n25, A2 => n412, B1 => n481, B2 => n2003, 
                           ZN => n2491);
   U3360 : NAND4_X1 port map( A1 => n2492, A2 => n2493, A3 => n2494, A4 => 
                           n2495, ZN => n2473);
   U3361 : AOI221_X1 port map( B1 => n2008, B2 => n6101, C1 => n2009, C2 => 
                           n6133, A => n2496, ZN => n2495);
   U3362 : OAI222_X1 port map( A1 => n4885, A2 => n2011, B1 => n4853, B2 => 
                           n2012, C1 => n4821, C2 => n418, ZN => n2496);
   U3363 : AOI221_X1 port map( B1 => n2013, B2 => n6165, C1 => n2014, C2 => 
                           n6197, A => n2497, ZN => n2494);
   U3364 : OAI22_X1 port map( A1 => n5570, A2 => n2016, B1 => n5571, B2 => 
                           n2017, ZN => n2497);
   U3365 : AOI221_X1 port map( B1 => n2018, B2 => n6229, C1 => n2019, C2 => 
                           n6261, A => n2498, ZN => n2493);
   U3366 : OAI222_X1 port map( A1 => n4981, A2 => n2021, B1 => n4949, B2 => 
                           n2022, C1 => n4917, C2 => n419, ZN => n2498);
   U3367 : AOI221_X1 port map( B1 => n2023, B2 => n578, C1 => n2024, C2 => n122
                           , A => n2499, ZN => n2492);
   U3368 : OAI22_X1 port map( A1 => n26, A2 => n2026, B1 => n482, B2 => n2027, 
                           ZN => n2499);
   U3369 : NAND4_X1 port map( A1 => n2500, A2 => n2501, A3 => n2502, A4 => 
                           n2503, ZN => n2472);
   U3370 : AOI221_X1 port map( B1 => n2032, B2 => n5845, C1 => n2033, C2 => 
                           n5877, A => n2504, ZN => n2503);
   U3371 : OAI222_X1 port map( A1 => n4629, A2 => n2035, B1 => n4597, B2 => 
                           n2036, C1 => n4565, C2 => n1577, ZN => n2504);
   U3372 : AOI221_X1 port map( B1 => n2037, B2 => n5909, C1 => n2038, C2 => 
                           n5941, A => n2505, ZN => n2502);
   U3373 : OAI22_X1 port map( A1 => n4693, A2 => n2040, B1 => n4661, B2 => 
                           n2041, ZN => n2505);
   U3374 : AOI221_X1 port map( B1 => n2042, B2 => n5973, C1 => n2043, C2 => 
                           n6005, A => n2506, ZN => n2501);
   U3375 : OAI222_X1 port map( A1 => n4789, A2 => n411, B1 => n4757, B2 => 
                           n2045, C1 => n4725, C2 => n2046, ZN => n2506);
   U3376 : AOI221_X1 port map( B1 => n2047, B2 => n6037, C1 => n2048, C2 => 
                           n6069, A => n2507, ZN => n2500);
   U3377 : OAI22_X1 port map( A1 => n5568, A2 => n2050, B1 => n5569, B2 => 
                           n2051, ZN => n2507);
   U3378 : OAI21_X1 port map( B1 => n1951, B2 => n1525, A => ENABLE, ZN => 
                           n7648);
   U3379 : OAI222_X1 port map( A1 => n2508, A2 => n1948, B1 => n2509, B2 => 
                           n1950, C1 => n1951, C2 => n1462, ZN => n7647);
   U3380 : NOR4_X1 port map( A1 => n2510, A2 => n2511, A3 => n2512, A4 => n2513
                           , ZN => n2509);
   U3381 : NAND4_X1 port map( A1 => n2514, A2 => n2515, A3 => n2516, A4 => 
                           n2517, ZN => n2513);
   U3382 : AOI221_X1 port map( B1 => n1960, B2 => n6420, C1 => n1961, C2 => 
                           n6452, A => n2518, ZN => n2517);
   U3383 : OAI222_X1 port map( A1 => n5268, A2 => n1963, B1 => n5236, B2 => 
                           n1964, C1 => n5204, C2 => n1965, ZN => n2518);
   U3384 : AOI221_X1 port map( B1 => n1966, B2 => n6484, C1 => n1967, C2 => 
                           n6516, A => n2519, ZN => n2516);
   U3385 : OAI22_X1 port map( A1 => n5564, A2 => n1969, B1 => n5565, B2 => 
                           n1970, ZN => n2519);
   U3386 : AOI221_X1 port map( B1 => n1971, B2 => n6548, C1 => n1972, C2 => 
                           n6580, A => n2520, ZN => n2515);
   U3387 : OAI222_X1 port map( A1 => n5364, A2 => n1974, B1 => n5332, B2 => 
                           n1578, C1 => n5300, C2 => n1975, ZN => n2520);
   U3388 : AOI221_X1 port map( B1 => n1976, B2 => n6612, C1 => n1977, C2 => 
                           n6644, A => n2521, ZN => n2514);
   U3389 : OAI22_X1 port map( A1 => n5566, A2 => n1756, B1 => n5567, B2 => 
                           n1980, ZN => n2521);
   U3390 : NAND4_X1 port map( A1 => n2522, A2 => n2523, A3 => n2524, A4 => 
                           n2525, ZN => n2512);
   U3391 : AOI221_X1 port map( B1 => n1985, B2 => n6292, C1 => n1986, C2 => 
                           n6324, A => n2526, ZN => n2525);
   U3392 : OAI222_X1 port map( A1 => n5076, A2 => n1988, B1 => n5044, B2 => 
                           n1989, C1 => n5012, C2 => n416, ZN => n2526);
   U3393 : AOI221_X1 port map( B1 => n1990, B2 => n174, C1 => n1991, C2 => n534
                           , A => n2527, ZN => n2524);
   U3394 : OAI22_X1 port map( A1 => n78, A2 => n1993, B1 => n438, B2 => n1994, 
                           ZN => n2527);
   U3395 : AOI221_X1 port map( B1 => n1995, B2 => n6356, C1 => n1996, C2 => 
                           n6388, A => n2528, ZN => n2523);
   U3396 : OAI222_X1 port map( A1 => n5172, A2 => n1998, B1 => n5140, B2 => 
                           n1999, C1 => n5108, C2 => n417, ZN => n2528);
   U3397 : AOI221_X1 port map( B1 => n2000, B2 => n579, C1 => n2001, C2 => n123
                           , A => n2529, ZN => n2522);
   U3398 : OAI22_X1 port map( A1 => n27, A2 => n412, B1 => n483, B2 => n2003, 
                           ZN => n2529);
   U3399 : NAND4_X1 port map( A1 => n2530, A2 => n2531, A3 => n2532, A4 => 
                           n2533, ZN => n2511);
   U3400 : AOI221_X1 port map( B1 => n2008, B2 => n6100, C1 => n2009, C2 => 
                           n6132, A => n2534, ZN => n2533);
   U3401 : OAI222_X1 port map( A1 => n4884, A2 => n2011, B1 => n4852, B2 => 
                           n2012, C1 => n4820, C2 => n418, ZN => n2534);
   U3402 : AOI221_X1 port map( B1 => n2013, B2 => n6164, C1 => n2014, C2 => 
                           n6196, A => n2535, ZN => n2532);
   U3403 : OAI22_X1 port map( A1 => n5560, A2 => n2016, B1 => n5561, B2 => 
                           n2017, ZN => n2535);
   U3404 : AOI221_X1 port map( B1 => n2018, B2 => n6228, C1 => n2019, C2 => 
                           n6260, A => n2536, ZN => n2531);
   U3405 : OAI222_X1 port map( A1 => n4980, A2 => n2021, B1 => n4948, B2 => 
                           n2022, C1 => n4916, C2 => n419, ZN => n2536);
   U3406 : AOI221_X1 port map( B1 => n2023, B2 => n580, C1 => n2024, C2 => n124
                           , A => n2537, ZN => n2530);
   U3407 : OAI22_X1 port map( A1 => n28, A2 => n2026, B1 => n484, B2 => n2027, 
                           ZN => n2537);
   U3408 : NAND4_X1 port map( A1 => n2538, A2 => n2539, A3 => n2540, A4 => 
                           n2541, ZN => n2510);
   U3409 : AOI221_X1 port map( B1 => n2032, B2 => n5844, C1 => n2033, C2 => 
                           n5876, A => n2542, ZN => n2541);
   U3410 : OAI222_X1 port map( A1 => n4628, A2 => n2035, B1 => n4596, B2 => 
                           n2036, C1 => n4564, C2 => n1577, ZN => n2542);
   U3411 : AOI221_X1 port map( B1 => n2037, B2 => n5908, C1 => n2038, C2 => 
                           n5940, A => n2543, ZN => n2540);
   U3412 : OAI22_X1 port map( A1 => n4692, A2 => n2040, B1 => n4660, B2 => 
                           n2041, ZN => n2543);
   U3413 : AOI221_X1 port map( B1 => n2042, B2 => n5972, C1 => n2043, C2 => 
                           n6004, A => n2544, ZN => n2539);
   U3414 : OAI222_X1 port map( A1 => n4788, A2 => n411, B1 => n4756, B2 => 
                           n2045, C1 => n4724, C2 => n2046, ZN => n2544);
   U3415 : AOI221_X1 port map( B1 => n2047, B2 => n6036, C1 => n2048, C2 => 
                           n6068, A => n2545, ZN => n2538);
   U3416 : OAI22_X1 port map( A1 => n5558, A2 => n2050, B1 => n5559, B2 => 
                           n2051, ZN => n2545);
   U3417 : OAI21_X1 port map( B1 => n1951, B2 => n1526, A => ENABLE, ZN => 
                           n7646);
   U3418 : OAI222_X1 port map( A1 => n2546, A2 => n1948, B1 => n2547, B2 => 
                           n1950, C1 => n1951, C2 => n1463, ZN => n7645);
   U3419 : NOR4_X1 port map( A1 => n2548, A2 => n2549, A3 => n2550, A4 => n2551
                           , ZN => n2547);
   U3420 : NAND4_X1 port map( A1 => n2552, A2 => n2553, A3 => n2554, A4 => 
                           n2555, ZN => n2551);
   U3421 : AOI221_X1 port map( B1 => n1960, B2 => n6419, C1 => n1961, C2 => 
                           n6451, A => n2556, ZN => n2555);
   U3422 : OAI222_X1 port map( A1 => n5267, A2 => n1963, B1 => n5235, B2 => 
                           n1964, C1 => n5203, C2 => n1965, ZN => n2556);
   U3423 : AOI221_X1 port map( B1 => n1966, B2 => n6483, C1 => n1967, C2 => 
                           n6515, A => n2557, ZN => n2554);
   U3424 : OAI22_X1 port map( A1 => n5554, A2 => n1969, B1 => n5555, B2 => 
                           n1970, ZN => n2557);
   U3425 : AOI221_X1 port map( B1 => n1971, B2 => n6547, C1 => n1972, C2 => 
                           n6579, A => n2558, ZN => n2553);
   U3426 : OAI222_X1 port map( A1 => n5363, A2 => n1974, B1 => n5331, B2 => 
                           n1578, C1 => n5299, C2 => n1975, ZN => n2558);
   U3427 : AOI221_X1 port map( B1 => n1976, B2 => n6611, C1 => n1977, C2 => 
                           n6643, A => n2559, ZN => n2552);
   U3428 : OAI22_X1 port map( A1 => n5556, A2 => n1756, B1 => n5557, B2 => 
                           n1980, ZN => n2559);
   U3429 : NAND4_X1 port map( A1 => n2560, A2 => n2561, A3 => n2562, A4 => 
                           n2563, ZN => n2550);
   U3430 : AOI221_X1 port map( B1 => n1985, B2 => n6291, C1 => n1986, C2 => 
                           n6323, A => n2564, ZN => n2563);
   U3431 : OAI222_X1 port map( A1 => n5075, A2 => n1988, B1 => n5043, B2 => 
                           n1989, C1 => n5011, C2 => n416, ZN => n2564);
   U3432 : AOI221_X1 port map( B1 => n1990, B2 => n175, C1 => n1991, C2 => n535
                           , A => n2565, ZN => n2562);
   U3433 : OAI22_X1 port map( A1 => n79, A2 => n1993, B1 => n439, B2 => n1994, 
                           ZN => n2565);
   U3434 : AOI221_X1 port map( B1 => n1995, B2 => n6355, C1 => n1996, C2 => 
                           n6387, A => n2566, ZN => n2561);
   U3435 : OAI222_X1 port map( A1 => n5171, A2 => n1998, B1 => n5139, B2 => 
                           n1999, C1 => n5107, C2 => n417, ZN => n2566);
   U3436 : AOI221_X1 port map( B1 => n2000, B2 => n581, C1 => n2001, C2 => n125
                           , A => n2567, ZN => n2560);
   U3437 : OAI22_X1 port map( A1 => n29, A2 => n412, B1 => n485, B2 => n2003, 
                           ZN => n2567);
   U3438 : NAND4_X1 port map( A1 => n2568, A2 => n2569, A3 => n2570, A4 => 
                           n2571, ZN => n2549);
   U3439 : AOI221_X1 port map( B1 => n2008, B2 => n6099, C1 => n2009, C2 => 
                           n6131, A => n2572, ZN => n2571);
   U3440 : OAI222_X1 port map( A1 => n4883, A2 => n2011, B1 => n4851, B2 => 
                           n2012, C1 => n4819, C2 => n418, ZN => n2572);
   U3441 : AOI221_X1 port map( B1 => n2013, B2 => n6163, C1 => n2014, C2 => 
                           n6195, A => n2573, ZN => n2570);
   U3442 : OAI22_X1 port map( A1 => n5550, A2 => n2016, B1 => n5551, B2 => 
                           n2017, ZN => n2573);
   U3443 : AOI221_X1 port map( B1 => n2018, B2 => n6227, C1 => n2019, C2 => 
                           n6259, A => n2574, ZN => n2569);
   U3444 : OAI222_X1 port map( A1 => n4979, A2 => n2021, B1 => n4947, B2 => 
                           n2022, C1 => n4915, C2 => n419, ZN => n2574);
   U3445 : AOI221_X1 port map( B1 => n2023, B2 => n582, C1 => n2024, C2 => n126
                           , A => n2575, ZN => n2568);
   U3446 : OAI22_X1 port map( A1 => n30, A2 => n2026, B1 => n486, B2 => n2027, 
                           ZN => n2575);
   U3447 : NAND4_X1 port map( A1 => n2576, A2 => n2577, A3 => n2578, A4 => 
                           n2579, ZN => n2548);
   U3448 : AOI221_X1 port map( B1 => n2032, B2 => n5843, C1 => n2033, C2 => 
                           n5875, A => n2580, ZN => n2579);
   U3449 : OAI222_X1 port map( A1 => n4627, A2 => n2035, B1 => n4595, B2 => 
                           n2036, C1 => n4563, C2 => n1577, ZN => n2580);
   U3450 : AOI221_X1 port map( B1 => n2037, B2 => n5907, C1 => n2038, C2 => 
                           n5939, A => n2581, ZN => n2578);
   U3451 : OAI22_X1 port map( A1 => n4691, A2 => n2040, B1 => n4659, B2 => 
                           n2041, ZN => n2581);
   U3452 : AOI221_X1 port map( B1 => n2042, B2 => n5971, C1 => n2043, C2 => 
                           n6003, A => n2582, ZN => n2577);
   U3453 : OAI222_X1 port map( A1 => n4787, A2 => n411, B1 => n4755, B2 => 
                           n2045, C1 => n4723, C2 => n2046, ZN => n2582);
   U3454 : AOI221_X1 port map( B1 => n2047, B2 => n6035, C1 => n2048, C2 => 
                           n6067, A => n2583, ZN => n2576);
   U3455 : OAI22_X1 port map( A1 => n5548, A2 => n2050, B1 => n5549, B2 => 
                           n2051, ZN => n2583);
   U3456 : OAI21_X1 port map( B1 => n1951, B2 => n1527, A => ENABLE, ZN => 
                           n7644);
   U3457 : OAI222_X1 port map( A1 => n2584, A2 => n1948, B1 => n2585, B2 => 
                           n1950, C1 => n1951, C2 => n1464, ZN => n7643);
   U3458 : NOR4_X1 port map( A1 => n2586, A2 => n2587, A3 => n2588, A4 => n2589
                           , ZN => n2585);
   U3459 : NAND4_X1 port map( A1 => n2590, A2 => n2591, A3 => n2592, A4 => 
                           n2593, ZN => n2589);
   U3460 : AOI221_X1 port map( B1 => n1960, B2 => n6418, C1 => n1961, C2 => 
                           n6450, A => n2594, ZN => n2593);
   U3461 : OAI222_X1 port map( A1 => n5266, A2 => n1963, B1 => n5234, B2 => 
                           n1964, C1 => n5202, C2 => n1965, ZN => n2594);
   U3462 : AOI221_X1 port map( B1 => n1966, B2 => n6482, C1 => n1967, C2 => 
                           n6514, A => n2595, ZN => n2592);
   U3463 : OAI22_X1 port map( A1 => n5544, A2 => n1969, B1 => n5545, B2 => 
                           n1970, ZN => n2595);
   U3464 : AOI221_X1 port map( B1 => n1971, B2 => n6546, C1 => n1972, C2 => 
                           n6578, A => n2596, ZN => n2591);
   U3465 : OAI222_X1 port map( A1 => n5362, A2 => n1974, B1 => n5330, B2 => 
                           n1578, C1 => n5298, C2 => n1975, ZN => n2596);
   U3466 : AOI221_X1 port map( B1 => n1976, B2 => n6610, C1 => n1977, C2 => 
                           n6642, A => n2597, ZN => n2590);
   U3467 : OAI22_X1 port map( A1 => n5546, A2 => n1756, B1 => n5547, B2 => 
                           n1980, ZN => n2597);
   U3468 : NAND4_X1 port map( A1 => n2598, A2 => n2599, A3 => n2600, A4 => 
                           n2601, ZN => n2588);
   U3469 : AOI221_X1 port map( B1 => n1985, B2 => n6290, C1 => n1986, C2 => 
                           n6322, A => n2602, ZN => n2601);
   U3470 : OAI222_X1 port map( A1 => n5074, A2 => n1988, B1 => n5042, B2 => 
                           n1989, C1 => n5010, C2 => n416, ZN => n2602);
   U3471 : AOI221_X1 port map( B1 => n1990, B2 => n176, C1 => n1991, C2 => n536
                           , A => n2603, ZN => n2600);
   U3472 : OAI22_X1 port map( A1 => n80, A2 => n1993, B1 => n440, B2 => n1994, 
                           ZN => n2603);
   U3473 : AOI221_X1 port map( B1 => n1995, B2 => n6354, C1 => n1996, C2 => 
                           n6386, A => n2604, ZN => n2599);
   U3474 : OAI222_X1 port map( A1 => n5170, A2 => n1998, B1 => n5138, B2 => 
                           n1999, C1 => n5106, C2 => n417, ZN => n2604);
   U3475 : AOI221_X1 port map( B1 => n2000, B2 => n583, C1 => n2001, C2 => n127
                           , A => n2605, ZN => n2598);
   U3476 : OAI22_X1 port map( A1 => n31, A2 => n412, B1 => n487, B2 => n2003, 
                           ZN => n2605);
   U3477 : NAND4_X1 port map( A1 => n2606, A2 => n2607, A3 => n2608, A4 => 
                           n2609, ZN => n2587);
   U3478 : AOI221_X1 port map( B1 => n2008, B2 => n6098, C1 => n2009, C2 => 
                           n6130, A => n2610, ZN => n2609);
   U3479 : OAI222_X1 port map( A1 => n4882, A2 => n2011, B1 => n4850, B2 => 
                           n2012, C1 => n4818, C2 => n418, ZN => n2610);
   U3480 : AOI221_X1 port map( B1 => n2013, B2 => n6162, C1 => n2014, C2 => 
                           n6194, A => n2611, ZN => n2608);
   U3481 : OAI22_X1 port map( A1 => n5540, A2 => n2016, B1 => n5541, B2 => 
                           n2017, ZN => n2611);
   U3482 : AOI221_X1 port map( B1 => n2018, B2 => n6226, C1 => n2019, C2 => 
                           n6258, A => n2612, ZN => n2607);
   U3483 : OAI222_X1 port map( A1 => n4978, A2 => n2021, B1 => n4946, B2 => 
                           n2022, C1 => n4914, C2 => n419, ZN => n2612);
   U3484 : AOI221_X1 port map( B1 => n2023, B2 => n584, C1 => n2024, C2 => n128
                           , A => n2613, ZN => n2606);
   U3485 : OAI22_X1 port map( A1 => n32, A2 => n2026, B1 => n488, B2 => n2027, 
                           ZN => n2613);
   U3486 : NAND4_X1 port map( A1 => n2614, A2 => n2615, A3 => n2616, A4 => 
                           n2617, ZN => n2586);
   U3487 : AOI221_X1 port map( B1 => n2032, B2 => n5842, C1 => n2033, C2 => 
                           n5874, A => n2618, ZN => n2617);
   U3488 : OAI222_X1 port map( A1 => n4626, A2 => n2035, B1 => n4594, B2 => 
                           n2036, C1 => n4562, C2 => n1577, ZN => n2618);
   U3489 : AOI221_X1 port map( B1 => n2037, B2 => n5906, C1 => n2038, C2 => 
                           n5938, A => n2619, ZN => n2616);
   U3490 : OAI22_X1 port map( A1 => n4690, A2 => n2040, B1 => n4658, B2 => 
                           n2041, ZN => n2619);
   U3491 : AOI221_X1 port map( B1 => n2042, B2 => n5970, C1 => n2043, C2 => 
                           n6002, A => n2620, ZN => n2615);
   U3492 : OAI222_X1 port map( A1 => n4786, A2 => n411, B1 => n4754, B2 => 
                           n2045, C1 => n4722, C2 => n2046, ZN => n2620);
   U3493 : AOI221_X1 port map( B1 => n2047, B2 => n6034, C1 => n2048, C2 => 
                           n6066, A => n2621, ZN => n2614);
   U3494 : OAI22_X1 port map( A1 => n5538, A2 => n2050, B1 => n5539, B2 => 
                           n2051, ZN => n2621);
   U3495 : OAI21_X1 port map( B1 => n1951, B2 => n1528, A => ENABLE, ZN => 
                           n7642);
   U3496 : OAI222_X1 port map( A1 => n2622, A2 => n1948, B1 => n2623, B2 => 
                           n1950, C1 => n1951, C2 => n1465, ZN => n7641);
   U3497 : NOR4_X1 port map( A1 => n2624, A2 => n2625, A3 => n2626, A4 => n2627
                           , ZN => n2623);
   U3498 : NAND4_X1 port map( A1 => n2628, A2 => n2629, A3 => n2630, A4 => 
                           n2631, ZN => n2627);
   U3499 : AOI221_X1 port map( B1 => n1960, B2 => n6417, C1 => n1961, C2 => 
                           n6449, A => n2632, ZN => n2631);
   U3500 : OAI222_X1 port map( A1 => n5265, A2 => n1963, B1 => n5233, B2 => 
                           n1964, C1 => n5201, C2 => n1965, ZN => n2632);
   U3501 : AOI221_X1 port map( B1 => n1966, B2 => n6481, C1 => n1967, C2 => 
                           n6513, A => n2633, ZN => n2630);
   U3502 : OAI22_X1 port map( A1 => n5534, A2 => n1969, B1 => n5535, B2 => 
                           n1970, ZN => n2633);
   U3503 : AOI221_X1 port map( B1 => n1971, B2 => n6545, C1 => n1972, C2 => 
                           n6577, A => n2634, ZN => n2629);
   U3504 : OAI222_X1 port map( A1 => n5361, A2 => n1974, B1 => n5329, B2 => 
                           n1578, C1 => n5297, C2 => n1975, ZN => n2634);
   U3505 : AOI221_X1 port map( B1 => n1976, B2 => n6609, C1 => n1977, C2 => 
                           n6641, A => n2635, ZN => n2628);
   U3506 : OAI22_X1 port map( A1 => n5536, A2 => n1756, B1 => n5537, B2 => 
                           n1980, ZN => n2635);
   U3507 : NAND4_X1 port map( A1 => n2636, A2 => n2637, A3 => n2638, A4 => 
                           n2639, ZN => n2626);
   U3508 : AOI221_X1 port map( B1 => n1985, B2 => n6289, C1 => n1986, C2 => 
                           n6321, A => n2640, ZN => n2639);
   U3509 : OAI222_X1 port map( A1 => n5073, A2 => n1988, B1 => n5041, B2 => 
                           n1989, C1 => n5009, C2 => n416, ZN => n2640);
   U3510 : AOI221_X1 port map( B1 => n1990, B2 => n177, C1 => n1991, C2 => n537
                           , A => n2641, ZN => n2638);
   U3511 : OAI22_X1 port map( A1 => n81, A2 => n1993, B1 => n441, B2 => n1994, 
                           ZN => n2641);
   U3512 : AOI221_X1 port map( B1 => n1995, B2 => n6353, C1 => n1996, C2 => 
                           n6385, A => n2642, ZN => n2637);
   U3513 : OAI222_X1 port map( A1 => n5169, A2 => n1998, B1 => n5137, B2 => 
                           n1999, C1 => n5105, C2 => n417, ZN => n2642);
   U3514 : AOI221_X1 port map( B1 => n2000, B2 => n585, C1 => n2001, C2 => n129
                           , A => n2643, ZN => n2636);
   U3515 : OAI22_X1 port map( A1 => n33, A2 => n412, B1 => n489, B2 => n2003, 
                           ZN => n2643);
   U3516 : NAND4_X1 port map( A1 => n2644, A2 => n2645, A3 => n2646, A4 => 
                           n2647, ZN => n2625);
   U3517 : AOI221_X1 port map( B1 => n2008, B2 => n6097, C1 => n2009, C2 => 
                           n6129, A => n2648, ZN => n2647);
   U3518 : OAI222_X1 port map( A1 => n4881, A2 => n2011, B1 => n4849, B2 => 
                           n2012, C1 => n4817, C2 => n418, ZN => n2648);
   U3519 : AOI221_X1 port map( B1 => n2013, B2 => n6161, C1 => n2014, C2 => 
                           n6193, A => n2649, ZN => n2646);
   U3520 : OAI22_X1 port map( A1 => n5530, A2 => n2016, B1 => n5531, B2 => 
                           n2017, ZN => n2649);
   U3521 : AOI221_X1 port map( B1 => n2018, B2 => n6225, C1 => n2019, C2 => 
                           n6257, A => n2650, ZN => n2645);
   U3522 : OAI222_X1 port map( A1 => n4977, A2 => n2021, B1 => n4945, B2 => 
                           n2022, C1 => n4913, C2 => n419, ZN => n2650);
   U3523 : AOI221_X1 port map( B1 => n2023, B2 => n586, C1 => n2024, C2 => n130
                           , A => n2651, ZN => n2644);
   U3524 : OAI22_X1 port map( A1 => n34, A2 => n2026, B1 => n490, B2 => n2027, 
                           ZN => n2651);
   U3525 : NAND4_X1 port map( A1 => n2652, A2 => n2653, A3 => n2654, A4 => 
                           n2655, ZN => n2624);
   U3526 : AOI221_X1 port map( B1 => n2032, B2 => n5841, C1 => n2033, C2 => 
                           n5873, A => n2656, ZN => n2655);
   U3527 : OAI222_X1 port map( A1 => n4625, A2 => n2035, B1 => n4593, B2 => 
                           n2036, C1 => n4561, C2 => n1577, ZN => n2656);
   U3528 : AOI221_X1 port map( B1 => n2037, B2 => n5905, C1 => n2038, C2 => 
                           n5937, A => n2657, ZN => n2654);
   U3529 : OAI22_X1 port map( A1 => n4689, A2 => n2040, B1 => n4657, B2 => 
                           n2041, ZN => n2657);
   U3530 : AOI221_X1 port map( B1 => n2042, B2 => n5969, C1 => n2043, C2 => 
                           n6001, A => n2658, ZN => n2653);
   U3531 : OAI222_X1 port map( A1 => n4785, A2 => n411, B1 => n4753, B2 => 
                           n2045, C1 => n4721, C2 => n2046, ZN => n2658);
   U3532 : AOI221_X1 port map( B1 => n2047, B2 => n6033, C1 => n2048, C2 => 
                           n6065, A => n2659, ZN => n2652);
   U3533 : OAI22_X1 port map( A1 => n5528, A2 => n2050, B1 => n5529, B2 => 
                           n2051, ZN => n2659);
   U3534 : OAI21_X1 port map( B1 => n1951, B2 => n1529, A => ENABLE, ZN => 
                           n7640);
   U3535 : OAI222_X1 port map( A1 => n2660, A2 => n1948, B1 => n2661, B2 => 
                           n1950, C1 => n1951, C2 => n1466, ZN => n7639);
   U3536 : NOR4_X1 port map( A1 => n2662, A2 => n2663, A3 => n2664, A4 => n2665
                           , ZN => n2661);
   U3537 : NAND4_X1 port map( A1 => n2666, A2 => n2667, A3 => n2668, A4 => 
                           n2669, ZN => n2665);
   U3538 : AOI221_X1 port map( B1 => n1960, B2 => n6416, C1 => n1961, C2 => 
                           n6448, A => n2670, ZN => n2669);
   U3539 : OAI222_X1 port map( A1 => n5264, A2 => n1963, B1 => n5232, B2 => 
                           n1964, C1 => n5200, C2 => n1965, ZN => n2670);
   U3540 : AOI221_X1 port map( B1 => n1966, B2 => n6480, C1 => n1967, C2 => 
                           n6512, A => n2671, ZN => n2668);
   U3541 : OAI22_X1 port map( A1 => n5524, A2 => n1969, B1 => n5525, B2 => 
                           n1970, ZN => n2671);
   U3542 : AOI221_X1 port map( B1 => n1971, B2 => n6544, C1 => n1972, C2 => 
                           n6576, A => n2672, ZN => n2667);
   U3543 : OAI222_X1 port map( A1 => n5360, A2 => n1974, B1 => n5328, B2 => 
                           n1578, C1 => n5296, C2 => n1975, ZN => n2672);
   U3544 : AOI221_X1 port map( B1 => n1976, B2 => n6608, C1 => n1977, C2 => 
                           n6640, A => n2673, ZN => n2666);
   U3545 : OAI22_X1 port map( A1 => n5526, A2 => n1756, B1 => n5527, B2 => 
                           n1980, ZN => n2673);
   U3546 : NAND4_X1 port map( A1 => n2674, A2 => n2675, A3 => n2676, A4 => 
                           n2677, ZN => n2664);
   U3547 : AOI221_X1 port map( B1 => n1985, B2 => n6288, C1 => n1986, C2 => 
                           n6320, A => n2678, ZN => n2677);
   U3548 : OAI222_X1 port map( A1 => n5072, A2 => n1988, B1 => n5040, B2 => 
                           n1989, C1 => n5008, C2 => n416, ZN => n2678);
   U3549 : AOI221_X1 port map( B1 => n1990, B2 => n178, C1 => n1991, C2 => n538
                           , A => n2679, ZN => n2676);
   U3550 : OAI22_X1 port map( A1 => n82, A2 => n1993, B1 => n442, B2 => n1994, 
                           ZN => n2679);
   U3551 : AOI221_X1 port map( B1 => n1995, B2 => n6352, C1 => n1996, C2 => 
                           n6384, A => n2680, ZN => n2675);
   U3552 : OAI222_X1 port map( A1 => n5168, A2 => n1998, B1 => n5136, B2 => 
                           n1999, C1 => n5104, C2 => n417, ZN => n2680);
   U3553 : AOI221_X1 port map( B1 => n2000, B2 => n587, C1 => n2001, C2 => n131
                           , A => n2681, ZN => n2674);
   U3554 : OAI22_X1 port map( A1 => n35, A2 => n412, B1 => n491, B2 => n2003, 
                           ZN => n2681);
   U3555 : NAND4_X1 port map( A1 => n2682, A2 => n2683, A3 => n2684, A4 => 
                           n2685, ZN => n2663);
   U3556 : AOI221_X1 port map( B1 => n2008, B2 => n6096, C1 => n2009, C2 => 
                           n6128, A => n2686, ZN => n2685);
   U3557 : OAI222_X1 port map( A1 => n4880, A2 => n2011, B1 => n4848, B2 => 
                           n2012, C1 => n4816, C2 => n418, ZN => n2686);
   U3558 : AOI221_X1 port map( B1 => n2013, B2 => n6160, C1 => n2014, C2 => 
                           n6192, A => n2687, ZN => n2684);
   U3559 : OAI22_X1 port map( A1 => n5520, A2 => n2016, B1 => n5521, B2 => 
                           n2017, ZN => n2687);
   U3560 : AOI221_X1 port map( B1 => n2018, B2 => n6224, C1 => n2019, C2 => 
                           n6256, A => n2688, ZN => n2683);
   U3561 : OAI222_X1 port map( A1 => n4976, A2 => n2021, B1 => n4944, B2 => 
                           n2022, C1 => n4912, C2 => n419, ZN => n2688);
   U3562 : AOI221_X1 port map( B1 => n2023, B2 => n588, C1 => n2024, C2 => n132
                           , A => n2689, ZN => n2682);
   U3563 : OAI22_X1 port map( A1 => n36, A2 => n2026, B1 => n492, B2 => n2027, 
                           ZN => n2689);
   U3564 : NAND4_X1 port map( A1 => n2690, A2 => n2691, A3 => n2692, A4 => 
                           n2693, ZN => n2662);
   U3565 : AOI221_X1 port map( B1 => n2032, B2 => n5840, C1 => n2033, C2 => 
                           n5872, A => n2694, ZN => n2693);
   U3566 : OAI222_X1 port map( A1 => n4624, A2 => n2035, B1 => n4592, B2 => 
                           n2036, C1 => n4560, C2 => n1577, ZN => n2694);
   U3567 : AOI221_X1 port map( B1 => n2037, B2 => n5904, C1 => n2038, C2 => 
                           n5936, A => n2695, ZN => n2692);
   U3568 : OAI22_X1 port map( A1 => n4688, A2 => n2040, B1 => n4656, B2 => 
                           n2041, ZN => n2695);
   U3569 : AOI221_X1 port map( B1 => n2042, B2 => n5968, C1 => n2043, C2 => 
                           n6000, A => n2696, ZN => n2691);
   U3570 : OAI222_X1 port map( A1 => n4784, A2 => n411, B1 => n4752, B2 => 
                           n2045, C1 => n4720, C2 => n2046, ZN => n2696);
   U3571 : AOI221_X1 port map( B1 => n2047, B2 => n6032, C1 => n2048, C2 => 
                           n6064, A => n2697, ZN => n2690);
   U3572 : OAI22_X1 port map( A1 => n5518, A2 => n2050, B1 => n5519, B2 => 
                           n2051, ZN => n2697);
   U3573 : OAI21_X1 port map( B1 => n1951, B2 => n1530, A => ENABLE, ZN => 
                           n7638);
   U3574 : OAI222_X1 port map( A1 => n2698, A2 => n1948, B1 => n2699, B2 => 
                           n1950, C1 => n1951, C2 => n1467, ZN => n7637);
   U3575 : NOR4_X1 port map( A1 => n2700, A2 => n2701, A3 => n2702, A4 => n2703
                           , ZN => n2699);
   U3576 : NAND4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => 
                           n2707, ZN => n2703);
   U3577 : AOI221_X1 port map( B1 => n1960, B2 => n6415, C1 => n1961, C2 => 
                           n6447, A => n2708, ZN => n2707);
   U3578 : OAI222_X1 port map( A1 => n5263, A2 => n1963, B1 => n5231, B2 => 
                           n1964, C1 => n5199, C2 => n1965, ZN => n2708);
   U3579 : AOI221_X1 port map( B1 => n1966, B2 => n6479, C1 => n1967, C2 => 
                           n6511, A => n2709, ZN => n2706);
   U3580 : OAI22_X1 port map( A1 => n5514, A2 => n1969, B1 => n5515, B2 => 
                           n1970, ZN => n2709);
   U3581 : AOI221_X1 port map( B1 => n1971, B2 => n6543, C1 => n1972, C2 => 
                           n6575, A => n2710, ZN => n2705);
   U3582 : OAI222_X1 port map( A1 => n5359, A2 => n1974, B1 => n5327, B2 => 
                           n1578, C1 => n5295, C2 => n1975, ZN => n2710);
   U3583 : AOI221_X1 port map( B1 => n1976, B2 => n6607, C1 => n1977, C2 => 
                           n6639, A => n2711, ZN => n2704);
   U3584 : OAI22_X1 port map( A1 => n5516, A2 => n1756, B1 => n5517, B2 => 
                           n1980, ZN => n2711);
   U3585 : NAND4_X1 port map( A1 => n2712, A2 => n2713, A3 => n2714, A4 => 
                           n2715, ZN => n2702);
   U3586 : AOI221_X1 port map( B1 => n1985, B2 => n6287, C1 => n1986, C2 => 
                           n6319, A => n2716, ZN => n2715);
   U3587 : OAI222_X1 port map( A1 => n5071, A2 => n1988, B1 => n5039, B2 => 
                           n1989, C1 => n5007, C2 => n416, ZN => n2716);
   U3588 : AOI221_X1 port map( B1 => n1990, B2 => n179, C1 => n1991, C2 => n539
                           , A => n2717, ZN => n2714);
   U3589 : OAI22_X1 port map( A1 => n83, A2 => n1993, B1 => n443, B2 => n1994, 
                           ZN => n2717);
   U3590 : AOI221_X1 port map( B1 => n1995, B2 => n6351, C1 => n1996, C2 => 
                           n6383, A => n2718, ZN => n2713);
   U3591 : OAI222_X1 port map( A1 => n5167, A2 => n1998, B1 => n5135, B2 => 
                           n1999, C1 => n5103, C2 => n417, ZN => n2718);
   U3592 : AOI221_X1 port map( B1 => n2000, B2 => n589, C1 => n2001, C2 => n133
                           , A => n2719, ZN => n2712);
   U3593 : OAI22_X1 port map( A1 => n37, A2 => n412, B1 => n493, B2 => n2003, 
                           ZN => n2719);
   U3594 : NAND4_X1 port map( A1 => n2720, A2 => n2721, A3 => n2722, A4 => 
                           n2723, ZN => n2701);
   U3595 : AOI221_X1 port map( B1 => n2008, B2 => n6095, C1 => n2009, C2 => 
                           n6127, A => n2724, ZN => n2723);
   U3596 : OAI222_X1 port map( A1 => n4879, A2 => n2011, B1 => n4847, B2 => 
                           n2012, C1 => n4815, C2 => n418, ZN => n2724);
   U3597 : AOI221_X1 port map( B1 => n2013, B2 => n6159, C1 => n2014, C2 => 
                           n6191, A => n2725, ZN => n2722);
   U3598 : OAI22_X1 port map( A1 => n5510, A2 => n2016, B1 => n5511, B2 => 
                           n2017, ZN => n2725);
   U3599 : AOI221_X1 port map( B1 => n2018, B2 => n6223, C1 => n2019, C2 => 
                           n6255, A => n2726, ZN => n2721);
   U3600 : OAI222_X1 port map( A1 => n4975, A2 => n2021, B1 => n4943, B2 => 
                           n2022, C1 => n4911, C2 => n419, ZN => n2726);
   U3601 : AOI221_X1 port map( B1 => n2023, B2 => n590, C1 => n2024, C2 => n134
                           , A => n2727, ZN => n2720);
   U3602 : OAI22_X1 port map( A1 => n38, A2 => n2026, B1 => n494, B2 => n2027, 
                           ZN => n2727);
   U3603 : NAND4_X1 port map( A1 => n2728, A2 => n2729, A3 => n2730, A4 => 
                           n2731, ZN => n2700);
   U3604 : AOI221_X1 port map( B1 => n2032, B2 => n5839, C1 => n2033, C2 => 
                           n5871, A => n2732, ZN => n2731);
   U3605 : OAI222_X1 port map( A1 => n4623, A2 => n2035, B1 => n4591, B2 => 
                           n2036, C1 => n4559, C2 => n1577, ZN => n2732);
   U3606 : AOI221_X1 port map( B1 => n2037, B2 => n5903, C1 => n2038, C2 => 
                           n5935, A => n2733, ZN => n2730);
   U3607 : OAI22_X1 port map( A1 => n4687, A2 => n2040, B1 => n4655, B2 => 
                           n2041, ZN => n2733);
   U3608 : AOI221_X1 port map( B1 => n2042, B2 => n5967, C1 => n2043, C2 => 
                           n5999, A => n2734, ZN => n2729);
   U3609 : OAI222_X1 port map( A1 => n4783, A2 => n411, B1 => n4751, B2 => 
                           n2045, C1 => n4719, C2 => n2046, ZN => n2734);
   U3610 : AOI221_X1 port map( B1 => n2047, B2 => n6031, C1 => n2048, C2 => 
                           n6063, A => n2735, ZN => n2728);
   U3611 : OAI22_X1 port map( A1 => n5508, A2 => n2050, B1 => n5509, B2 => 
                           n2051, ZN => n2735);
   U3612 : OAI21_X1 port map( B1 => n1951, B2 => n1531, A => ENABLE, ZN => 
                           n7636);
   U3613 : OAI222_X1 port map( A1 => n2736, A2 => n1948, B1 => n2737, B2 => 
                           n1950, C1 => n1951, C2 => n1468, ZN => n7635);
   U3614 : NOR4_X1 port map( A1 => n2738, A2 => n2739, A3 => n2740, A4 => n2741
                           , ZN => n2737);
   U3615 : NAND4_X1 port map( A1 => n2742, A2 => n2743, A3 => n2744, A4 => 
                           n2745, ZN => n2741);
   U3616 : AOI221_X1 port map( B1 => n1960, B2 => n6414, C1 => n1961, C2 => 
                           n6446, A => n2746, ZN => n2745);
   U3617 : OAI222_X1 port map( A1 => n5262, A2 => n1963, B1 => n5230, B2 => 
                           n1964, C1 => n5198, C2 => n1965, ZN => n2746);
   U3618 : AOI221_X1 port map( B1 => n1966, B2 => n6478, C1 => n1967, C2 => 
                           n6510, A => n2747, ZN => n2744);
   U3619 : OAI22_X1 port map( A1 => n5504, A2 => n1969, B1 => n5505, B2 => 
                           n1970, ZN => n2747);
   U3620 : AOI221_X1 port map( B1 => n1971, B2 => n6542, C1 => n1972, C2 => 
                           n6574, A => n2748, ZN => n2743);
   U3621 : OAI222_X1 port map( A1 => n5358, A2 => n1974, B1 => n5326, B2 => 
                           n1578, C1 => n5294, C2 => n1975, ZN => n2748);
   U3622 : AOI221_X1 port map( B1 => n1976, B2 => n6606, C1 => n1977, C2 => 
                           n6638, A => n2749, ZN => n2742);
   U3623 : OAI22_X1 port map( A1 => n5506, A2 => n1756, B1 => n5507, B2 => 
                           n1980, ZN => n2749);
   U3624 : NAND4_X1 port map( A1 => n2750, A2 => n2751, A3 => n2752, A4 => 
                           n2753, ZN => n2740);
   U3625 : AOI221_X1 port map( B1 => n1985, B2 => n6286, C1 => n1986, C2 => 
                           n6318, A => n2754, ZN => n2753);
   U3626 : OAI222_X1 port map( A1 => n5070, A2 => n1988, B1 => n5038, B2 => 
                           n1989, C1 => n5006, C2 => n416, ZN => n2754);
   U3627 : AOI221_X1 port map( B1 => n1990, B2 => n180, C1 => n1991, C2 => n540
                           , A => n2755, ZN => n2752);
   U3628 : OAI22_X1 port map( A1 => n84, A2 => n1993, B1 => n444, B2 => n1994, 
                           ZN => n2755);
   U3629 : AOI221_X1 port map( B1 => n1995, B2 => n6350, C1 => n1996, C2 => 
                           n6382, A => n2756, ZN => n2751);
   U3630 : OAI222_X1 port map( A1 => n5166, A2 => n1998, B1 => n5134, B2 => 
                           n1999, C1 => n5102, C2 => n417, ZN => n2756);
   U3631 : AOI221_X1 port map( B1 => n2000, B2 => n591, C1 => n2001, C2 => n135
                           , A => n2757, ZN => n2750);
   U3632 : OAI22_X1 port map( A1 => n39, A2 => n412, B1 => n495, B2 => n2003, 
                           ZN => n2757);
   U3633 : NAND4_X1 port map( A1 => n2758, A2 => n2759, A3 => n2760, A4 => 
                           n2761, ZN => n2739);
   U3634 : AOI221_X1 port map( B1 => n2008, B2 => n6094, C1 => n2009, C2 => 
                           n6126, A => n2762, ZN => n2761);
   U3635 : OAI222_X1 port map( A1 => n4878, A2 => n2011, B1 => n4846, B2 => 
                           n2012, C1 => n4814, C2 => n418, ZN => n2762);
   U3636 : AOI221_X1 port map( B1 => n2013, B2 => n6158, C1 => n2014, C2 => 
                           n6190, A => n2763, ZN => n2760);
   U3637 : OAI22_X1 port map( A1 => n5500, A2 => n2016, B1 => n5501, B2 => 
                           n2017, ZN => n2763);
   U3638 : AOI221_X1 port map( B1 => n2018, B2 => n6222, C1 => n2019, C2 => 
                           n6254, A => n2764, ZN => n2759);
   U3639 : OAI222_X1 port map( A1 => n4974, A2 => n2021, B1 => n4942, B2 => 
                           n2022, C1 => n4910, C2 => n419, ZN => n2764);
   U3640 : AOI221_X1 port map( B1 => n2023, B2 => n592, C1 => n2024, C2 => n136
                           , A => n2765, ZN => n2758);
   U3641 : OAI22_X1 port map( A1 => n40, A2 => n2026, B1 => n496, B2 => n2027, 
                           ZN => n2765);
   U3642 : NAND4_X1 port map( A1 => n2766, A2 => n2767, A3 => n2768, A4 => 
                           n2769, ZN => n2738);
   U3643 : AOI221_X1 port map( B1 => n2032, B2 => n5838, C1 => n2033, C2 => 
                           n5870, A => n2770, ZN => n2769);
   U3644 : OAI222_X1 port map( A1 => n4622, A2 => n2035, B1 => n4590, B2 => 
                           n2036, C1 => n4558, C2 => n1577, ZN => n2770);
   U3645 : AOI221_X1 port map( B1 => n2037, B2 => n5902, C1 => n2038, C2 => 
                           n5934, A => n2771, ZN => n2768);
   U3646 : OAI22_X1 port map( A1 => n4686, A2 => n2040, B1 => n4654, B2 => 
                           n2041, ZN => n2771);
   U3647 : AOI221_X1 port map( B1 => n2042, B2 => n5966, C1 => n2043, C2 => 
                           n5998, A => n2772, ZN => n2767);
   U3648 : OAI222_X1 port map( A1 => n4782, A2 => n411, B1 => n4750, B2 => 
                           n2045, C1 => n4718, C2 => n2046, ZN => n2772);
   U3649 : AOI221_X1 port map( B1 => n2047, B2 => n6030, C1 => n2048, C2 => 
                           n6062, A => n2773, ZN => n2766);
   U3650 : OAI22_X1 port map( A1 => n5498, A2 => n2050, B1 => n5499, B2 => 
                           n2051, ZN => n2773);
   U3651 : OAI21_X1 port map( B1 => n1951, B2 => n1532, A => ENABLE, ZN => 
                           n7634);
   U3652 : OAI222_X1 port map( A1 => n2774, A2 => n1948, B1 => n2775, B2 => 
                           n1950, C1 => n1951, C2 => n1469, ZN => n7633);
   U3653 : NOR4_X1 port map( A1 => n2776, A2 => n2777, A3 => n2778, A4 => n2779
                           , ZN => n2775);
   U3654 : NAND4_X1 port map( A1 => n2780, A2 => n2781, A3 => n2782, A4 => 
                           n2783, ZN => n2779);
   U3655 : AOI221_X1 port map( B1 => n1960, B2 => n6413, C1 => n1961, C2 => 
                           n6445, A => n2784, ZN => n2783);
   U3656 : OAI222_X1 port map( A1 => n5261, A2 => n1963, B1 => n5229, B2 => 
                           n1964, C1 => n5197, C2 => n1965, ZN => n2784);
   U3657 : AOI221_X1 port map( B1 => n1966, B2 => n6477, C1 => n1967, C2 => 
                           n6509, A => n2785, ZN => n2782);
   U3658 : OAI22_X1 port map( A1 => n5494, A2 => n1969, B1 => n5495, B2 => 
                           n1970, ZN => n2785);
   U3659 : AOI221_X1 port map( B1 => n1971, B2 => n6541, C1 => n1972, C2 => 
                           n6573, A => n2786, ZN => n2781);
   U3660 : OAI222_X1 port map( A1 => n5357, A2 => n1974, B1 => n5325, B2 => 
                           n1578, C1 => n5293, C2 => n1975, ZN => n2786);
   U3661 : AOI221_X1 port map( B1 => n1976, B2 => n6605, C1 => n1977, C2 => 
                           n6637, A => n2787, ZN => n2780);
   U3662 : OAI22_X1 port map( A1 => n5496, A2 => n1756, B1 => n5497, B2 => 
                           n1980, ZN => n2787);
   U3663 : NAND4_X1 port map( A1 => n2788, A2 => n2789, A3 => n2790, A4 => 
                           n2791, ZN => n2778);
   U3664 : AOI221_X1 port map( B1 => n1985, B2 => n6285, C1 => n1986, C2 => 
                           n6317, A => n2792, ZN => n2791);
   U3665 : OAI222_X1 port map( A1 => n5069, A2 => n1988, B1 => n5037, B2 => 
                           n1989, C1 => n5005, C2 => n416, ZN => n2792);
   U3666 : AOI221_X1 port map( B1 => n1990, B2 => n181, C1 => n1991, C2 => n541
                           , A => n2793, ZN => n2790);
   U3667 : OAI22_X1 port map( A1 => n85, A2 => n1993, B1 => n445, B2 => n1994, 
                           ZN => n2793);
   U3668 : AOI221_X1 port map( B1 => n1995, B2 => n6349, C1 => n1996, C2 => 
                           n6381, A => n2794, ZN => n2789);
   U3669 : OAI222_X1 port map( A1 => n5165, A2 => n1998, B1 => n5133, B2 => 
                           n1999, C1 => n5101, C2 => n417, ZN => n2794);
   U3670 : AOI221_X1 port map( B1 => n2000, B2 => n593, C1 => n2001, C2 => n137
                           , A => n2795, ZN => n2788);
   U3671 : OAI22_X1 port map( A1 => n41, A2 => n412, B1 => n497, B2 => n2003, 
                           ZN => n2795);
   U3672 : NAND4_X1 port map( A1 => n2796, A2 => n2797, A3 => n2798, A4 => 
                           n2799, ZN => n2777);
   U3673 : AOI221_X1 port map( B1 => n2008, B2 => n6093, C1 => n2009, C2 => 
                           n6125, A => n2800, ZN => n2799);
   U3674 : OAI222_X1 port map( A1 => n4877, A2 => n2011, B1 => n4845, B2 => 
                           n2012, C1 => n4813, C2 => n418, ZN => n2800);
   U3675 : AOI221_X1 port map( B1 => n2013, B2 => n6157, C1 => n2014, C2 => 
                           n6189, A => n2801, ZN => n2798);
   U3676 : OAI22_X1 port map( A1 => n5490, A2 => n2016, B1 => n5491, B2 => 
                           n2017, ZN => n2801);
   U3677 : AOI221_X1 port map( B1 => n2018, B2 => n6221, C1 => n2019, C2 => 
                           n6253, A => n2802, ZN => n2797);
   U3678 : OAI222_X1 port map( A1 => n4973, A2 => n2021, B1 => n4941, B2 => 
                           n2022, C1 => n4909, C2 => n419, ZN => n2802);
   U3679 : AOI221_X1 port map( B1 => n2023, B2 => n594, C1 => n2024, C2 => n138
                           , A => n2803, ZN => n2796);
   U3680 : OAI22_X1 port map( A1 => n42, A2 => n2026, B1 => n498, B2 => n2027, 
                           ZN => n2803);
   U3681 : NAND4_X1 port map( A1 => n2804, A2 => n2805, A3 => n2806, A4 => 
                           n2807, ZN => n2776);
   U3682 : AOI221_X1 port map( B1 => n2032, B2 => n5837, C1 => n2033, C2 => 
                           n5869, A => n2808, ZN => n2807);
   U3683 : OAI222_X1 port map( A1 => n4621, A2 => n2035, B1 => n4589, B2 => 
                           n2036, C1 => n4557, C2 => n1577, ZN => n2808);
   U3684 : AOI221_X1 port map( B1 => n2037, B2 => n5901, C1 => n2038, C2 => 
                           n5933, A => n2809, ZN => n2806);
   U3685 : OAI22_X1 port map( A1 => n4685, A2 => n2040, B1 => n4653, B2 => 
                           n2041, ZN => n2809);
   U3686 : AOI221_X1 port map( B1 => n2042, B2 => n5965, C1 => n2043, C2 => 
                           n5997, A => n2810, ZN => n2805);
   U3687 : OAI222_X1 port map( A1 => n4781, A2 => n411, B1 => n4749, B2 => 
                           n2045, C1 => n4717, C2 => n2046, ZN => n2810);
   U3688 : AOI221_X1 port map( B1 => n2047, B2 => n6029, C1 => n2048, C2 => 
                           n6061, A => n2811, ZN => n2804);
   U3689 : OAI22_X1 port map( A1 => n5488, A2 => n2050, B1 => n5489, B2 => 
                           n2051, ZN => n2811);
   U3690 : OAI21_X1 port map( B1 => n1951, B2 => n1533, A => ENABLE, ZN => 
                           n7632);
   U3691 : OAI222_X1 port map( A1 => n2812, A2 => n1948, B1 => n2813, B2 => 
                           n1950, C1 => n1951, C2 => n1470, ZN => n7631);
   U3692 : NOR4_X1 port map( A1 => n2814, A2 => n2815, A3 => n2816, A4 => n2817
                           , ZN => n2813);
   U3693 : NAND4_X1 port map( A1 => n2818, A2 => n2819, A3 => n2820, A4 => 
                           n2821, ZN => n2817);
   U3694 : AOI221_X1 port map( B1 => n1960, B2 => n6412, C1 => n1961, C2 => 
                           n6444, A => n2822, ZN => n2821);
   U3695 : OAI222_X1 port map( A1 => n5260, A2 => n1963, B1 => n5228, B2 => 
                           n1964, C1 => n5196, C2 => n1965, ZN => n2822);
   U3696 : AOI221_X1 port map( B1 => n1966, B2 => n6476, C1 => n1967, C2 => 
                           n6508, A => n2823, ZN => n2820);
   U3697 : OAI22_X1 port map( A1 => n5484, A2 => n1969, B1 => n5485, B2 => 
                           n1970, ZN => n2823);
   U3698 : AOI221_X1 port map( B1 => n1971, B2 => n6540, C1 => n1972, C2 => 
                           n6572, A => n2824, ZN => n2819);
   U3699 : OAI222_X1 port map( A1 => n5356, A2 => n1974, B1 => n5324, B2 => 
                           n1578, C1 => n5292, C2 => n1975, ZN => n2824);
   U3700 : AOI221_X1 port map( B1 => n1976, B2 => n6604, C1 => n1977, C2 => 
                           n6636, A => n2825, ZN => n2818);
   U3701 : OAI22_X1 port map( A1 => n5486, A2 => n1756, B1 => n5487, B2 => 
                           n1980, ZN => n2825);
   U3702 : NAND4_X1 port map( A1 => n2826, A2 => n2827, A3 => n2828, A4 => 
                           n2829, ZN => n2816);
   U3703 : AOI221_X1 port map( B1 => n1985, B2 => n6284, C1 => n1986, C2 => 
                           n6316, A => n2830, ZN => n2829);
   U3704 : OAI222_X1 port map( A1 => n5068, A2 => n1988, B1 => n5036, B2 => 
                           n1989, C1 => n5004, C2 => n416, ZN => n2830);
   U3705 : AOI221_X1 port map( B1 => n1990, B2 => n182, C1 => n1991, C2 => n542
                           , A => n2831, ZN => n2828);
   U3706 : OAI22_X1 port map( A1 => n86, A2 => n1993, B1 => n446, B2 => n1994, 
                           ZN => n2831);
   U3707 : AOI221_X1 port map( B1 => n1995, B2 => n6348, C1 => n1996, C2 => 
                           n6380, A => n2832, ZN => n2827);
   U3708 : OAI222_X1 port map( A1 => n5164, A2 => n1998, B1 => n5132, B2 => 
                           n1999, C1 => n5100, C2 => n417, ZN => n2832);
   U3709 : AOI221_X1 port map( B1 => n2000, B2 => n595, C1 => n2001, C2 => n139
                           , A => n2833, ZN => n2826);
   U3710 : OAI22_X1 port map( A1 => n43, A2 => n412, B1 => n499, B2 => n2003, 
                           ZN => n2833);
   U3711 : NAND4_X1 port map( A1 => n2834, A2 => n2835, A3 => n2836, A4 => 
                           n2837, ZN => n2815);
   U3712 : AOI221_X1 port map( B1 => n2008, B2 => n6092, C1 => n2009, C2 => 
                           n6124, A => n2838, ZN => n2837);
   U3713 : OAI222_X1 port map( A1 => n4876, A2 => n2011, B1 => n4844, B2 => 
                           n2012, C1 => n4812, C2 => n418, ZN => n2838);
   U3714 : AOI221_X1 port map( B1 => n2013, B2 => n6156, C1 => n2014, C2 => 
                           n6188, A => n2839, ZN => n2836);
   U3715 : OAI22_X1 port map( A1 => n5480, A2 => n2016, B1 => n5481, B2 => 
                           n2017, ZN => n2839);
   U3716 : AOI221_X1 port map( B1 => n2018, B2 => n6220, C1 => n2019, C2 => 
                           n6252, A => n2840, ZN => n2835);
   U3717 : OAI222_X1 port map( A1 => n4972, A2 => n2021, B1 => n4940, B2 => 
                           n2022, C1 => n4908, C2 => n419, ZN => n2840);
   U3718 : AOI221_X1 port map( B1 => n2023, B2 => n596, C1 => n2024, C2 => n140
                           , A => n2841, ZN => n2834);
   U3719 : OAI22_X1 port map( A1 => n44, A2 => n2026, B1 => n500, B2 => n2027, 
                           ZN => n2841);
   U3720 : NAND4_X1 port map( A1 => n2842, A2 => n2843, A3 => n2844, A4 => 
                           n2845, ZN => n2814);
   U3721 : AOI221_X1 port map( B1 => n2032, B2 => n5836, C1 => n2033, C2 => 
                           n5868, A => n2846, ZN => n2845);
   U3722 : OAI222_X1 port map( A1 => n4620, A2 => n2035, B1 => n4588, B2 => 
                           n2036, C1 => n4556, C2 => n1577, ZN => n2846);
   U3723 : AOI221_X1 port map( B1 => n2037, B2 => n5900, C1 => n2038, C2 => 
                           n5932, A => n2847, ZN => n2844);
   U3724 : OAI22_X1 port map( A1 => n4684, A2 => n2040, B1 => n4652, B2 => 
                           n2041, ZN => n2847);
   U3725 : AOI221_X1 port map( B1 => n2042, B2 => n5964, C1 => n2043, C2 => 
                           n5996, A => n2848, ZN => n2843);
   U3726 : OAI222_X1 port map( A1 => n4780, A2 => n411, B1 => n4748, B2 => 
                           n2045, C1 => n4716, C2 => n2046, ZN => n2848);
   U3727 : AOI221_X1 port map( B1 => n2047, B2 => n6028, C1 => n2048, C2 => 
                           n6060, A => n2849, ZN => n2842);
   U3728 : OAI22_X1 port map( A1 => n5478, A2 => n2050, B1 => n5479, B2 => 
                           n2051, ZN => n2849);
   U3729 : OAI21_X1 port map( B1 => n1951, B2 => n1534, A => ENABLE, ZN => 
                           n7630);
   U3730 : OAI222_X1 port map( A1 => n2850, A2 => n1948, B1 => n2851, B2 => 
                           n1950, C1 => n1951, C2 => n1471, ZN => n7629);
   U3731 : NOR4_X1 port map( A1 => n2852, A2 => n2853, A3 => n2854, A4 => n2855
                           , ZN => n2851);
   U3732 : NAND4_X1 port map( A1 => n2856, A2 => n2857, A3 => n2858, A4 => 
                           n2859, ZN => n2855);
   U3733 : AOI221_X1 port map( B1 => n1960, B2 => n6411, C1 => n1961, C2 => 
                           n6443, A => n2860, ZN => n2859);
   U3734 : OAI222_X1 port map( A1 => n5259, A2 => n1963, B1 => n5227, B2 => 
                           n1964, C1 => n5195, C2 => n1965, ZN => n2860);
   U3735 : AOI221_X1 port map( B1 => n1966, B2 => n6475, C1 => n1967, C2 => 
                           n6507, A => n2861, ZN => n2858);
   U3736 : OAI22_X1 port map( A1 => n5474, A2 => n1969, B1 => n5475, B2 => 
                           n1970, ZN => n2861);
   U3737 : AOI221_X1 port map( B1 => n1971, B2 => n6539, C1 => n1972, C2 => 
                           n6571, A => n2862, ZN => n2857);
   U3738 : OAI222_X1 port map( A1 => n5355, A2 => n1974, B1 => n5323, B2 => 
                           n1578, C1 => n5291, C2 => n1975, ZN => n2862);
   U3739 : AOI221_X1 port map( B1 => n1976, B2 => n6603, C1 => n1977, C2 => 
                           n6635, A => n2863, ZN => n2856);
   U3740 : OAI22_X1 port map( A1 => n5476, A2 => n1756, B1 => n5477, B2 => 
                           n1980, ZN => n2863);
   U3741 : NAND4_X1 port map( A1 => n2864, A2 => n2865, A3 => n2866, A4 => 
                           n2867, ZN => n2854);
   U3742 : AOI221_X1 port map( B1 => n1985, B2 => n6283, C1 => n1986, C2 => 
                           n6315, A => n2868, ZN => n2867);
   U3743 : OAI222_X1 port map( A1 => n5067, A2 => n1988, B1 => n5035, B2 => 
                           n1989, C1 => n5003, C2 => n416, ZN => n2868);
   U3744 : AOI221_X1 port map( B1 => n1990, B2 => n183, C1 => n1991, C2 => n543
                           , A => n2869, ZN => n2866);
   U3745 : OAI22_X1 port map( A1 => n87, A2 => n1993, B1 => n447, B2 => n1994, 
                           ZN => n2869);
   U3746 : AOI221_X1 port map( B1 => n1995, B2 => n6347, C1 => n1996, C2 => 
                           n6379, A => n2870, ZN => n2865);
   U3747 : OAI222_X1 port map( A1 => n5163, A2 => n1998, B1 => n5131, B2 => 
                           n1999, C1 => n5099, C2 => n417, ZN => n2870);
   U3748 : AOI221_X1 port map( B1 => n2000, B2 => n597, C1 => n2001, C2 => n141
                           , A => n2871, ZN => n2864);
   U3749 : OAI22_X1 port map( A1 => n45, A2 => n412, B1 => n501, B2 => n2003, 
                           ZN => n2871);
   U3750 : NAND4_X1 port map( A1 => n2872, A2 => n2873, A3 => n2874, A4 => 
                           n2875, ZN => n2853);
   U3751 : AOI221_X1 port map( B1 => n2008, B2 => n6091, C1 => n2009, C2 => 
                           n6123, A => n2876, ZN => n2875);
   U3752 : OAI222_X1 port map( A1 => n4875, A2 => n2011, B1 => n4843, B2 => 
                           n2012, C1 => n4811, C2 => n418, ZN => n2876);
   U3753 : AOI221_X1 port map( B1 => n2013, B2 => n6155, C1 => n2014, C2 => 
                           n6187, A => n2877, ZN => n2874);
   U3754 : OAI22_X1 port map( A1 => n5470, A2 => n2016, B1 => n5471, B2 => 
                           n2017, ZN => n2877);
   U3755 : AOI221_X1 port map( B1 => n2018, B2 => n6219, C1 => n2019, C2 => 
                           n6251, A => n2878, ZN => n2873);
   U3756 : OAI222_X1 port map( A1 => n4971, A2 => n2021, B1 => n4939, B2 => 
                           n2022, C1 => n4907, C2 => n419, ZN => n2878);
   U3757 : AOI221_X1 port map( B1 => n2023, B2 => n598, C1 => n2024, C2 => n142
                           , A => n2879, ZN => n2872);
   U3758 : OAI22_X1 port map( A1 => n46, A2 => n2026, B1 => n502, B2 => n2027, 
                           ZN => n2879);
   U3759 : NAND4_X1 port map( A1 => n2880, A2 => n2881, A3 => n2882, A4 => 
                           n2883, ZN => n2852);
   U3760 : AOI221_X1 port map( B1 => n2032, B2 => n5835, C1 => n2033, C2 => 
                           n5867, A => n2884, ZN => n2883);
   U3761 : OAI222_X1 port map( A1 => n4619, A2 => n2035, B1 => n4587, B2 => 
                           n2036, C1 => n4555, C2 => n1577, ZN => n2884);
   U3762 : AOI221_X1 port map( B1 => n2037, B2 => n5899, C1 => n2038, C2 => 
                           n5931, A => n2885, ZN => n2882);
   U3763 : OAI22_X1 port map( A1 => n4683, A2 => n2040, B1 => n4651, B2 => 
                           n2041, ZN => n2885);
   U3764 : AOI221_X1 port map( B1 => n2042, B2 => n5963, C1 => n2043, C2 => 
                           n5995, A => n2886, ZN => n2881);
   U3765 : OAI222_X1 port map( A1 => n4779, A2 => n411, B1 => n4747, B2 => 
                           n2045, C1 => n4715, C2 => n2046, ZN => n2886);
   U3766 : AOI221_X1 port map( B1 => n2047, B2 => n6027, C1 => n2048, C2 => 
                           n6059, A => n2887, ZN => n2880);
   U3767 : OAI22_X1 port map( A1 => n5468, A2 => n2050, B1 => n5469, B2 => 
                           n2051, ZN => n2887);
   U3768 : OAI21_X1 port map( B1 => n1951, B2 => n1535, A => ENABLE, ZN => 
                           n7628);
   U3769 : OAI222_X1 port map( A1 => n2888, A2 => n1948, B1 => n2889, B2 => 
                           n1950, C1 => n1951, C2 => n1472, ZN => n7627);
   U3770 : NOR4_X1 port map( A1 => n2890, A2 => n2891, A3 => n2892, A4 => n2893
                           , ZN => n2889);
   U3771 : NAND4_X1 port map( A1 => n2894, A2 => n2895, A3 => n2896, A4 => 
                           n2897, ZN => n2893);
   U3772 : AOI221_X1 port map( B1 => n1960, B2 => n6410, C1 => n1961, C2 => 
                           n6442, A => n2898, ZN => n2897);
   U3773 : OAI222_X1 port map( A1 => n5258, A2 => n1963, B1 => n5226, B2 => 
                           n1964, C1 => n5194, C2 => n1965, ZN => n2898);
   U3774 : AOI221_X1 port map( B1 => n1966, B2 => n6474, C1 => n1967, C2 => 
                           n6506, A => n2899, ZN => n2896);
   U3775 : OAI22_X1 port map( A1 => n5464, A2 => n1969, B1 => n5465, B2 => 
                           n1970, ZN => n2899);
   U3776 : AOI221_X1 port map( B1 => n1971, B2 => n6538, C1 => n1972, C2 => 
                           n6570, A => n2900, ZN => n2895);
   U3777 : OAI222_X1 port map( A1 => n5354, A2 => n1974, B1 => n5322, B2 => 
                           n1578, C1 => n5290, C2 => n1975, ZN => n2900);
   U3778 : AOI221_X1 port map( B1 => n1976, B2 => n6602, C1 => n1977, C2 => 
                           n6634, A => n2901, ZN => n2894);
   U3779 : OAI22_X1 port map( A1 => n5466, A2 => n1756, B1 => n5467, B2 => 
                           n1980, ZN => n2901);
   U3780 : NAND4_X1 port map( A1 => n2902, A2 => n2903, A3 => n2904, A4 => 
                           n2905, ZN => n2892);
   U3781 : AOI221_X1 port map( B1 => n1985, B2 => n6282, C1 => n1986, C2 => 
                           n6314, A => n2906, ZN => n2905);
   U3782 : OAI222_X1 port map( A1 => n5066, A2 => n1988, B1 => n5034, B2 => 
                           n1989, C1 => n5002, C2 => n416, ZN => n2906);
   U3783 : AOI221_X1 port map( B1 => n1990, B2 => n184, C1 => n1991, C2 => n544
                           , A => n2907, ZN => n2904);
   U3784 : OAI22_X1 port map( A1 => n88, A2 => n1993, B1 => n448, B2 => n1994, 
                           ZN => n2907);
   U3785 : AOI221_X1 port map( B1 => n1995, B2 => n6346, C1 => n1996, C2 => 
                           n6378, A => n2908, ZN => n2903);
   U3786 : OAI222_X1 port map( A1 => n5162, A2 => n1998, B1 => n5130, B2 => 
                           n1999, C1 => n5098, C2 => n417, ZN => n2908);
   U3787 : AOI221_X1 port map( B1 => n2000, B2 => n599, C1 => n2001, C2 => n143
                           , A => n2909, ZN => n2902);
   U3788 : OAI22_X1 port map( A1 => n47, A2 => n412, B1 => n503, B2 => n2003, 
                           ZN => n2909);
   U3789 : NAND4_X1 port map( A1 => n2910, A2 => n2911, A3 => n2912, A4 => 
                           n2913, ZN => n2891);
   U3790 : AOI221_X1 port map( B1 => n2008, B2 => n6090, C1 => n2009, C2 => 
                           n6122, A => n2914, ZN => n2913);
   U3791 : OAI222_X1 port map( A1 => n4874, A2 => n2011, B1 => n4842, B2 => 
                           n2012, C1 => n4810, C2 => n418, ZN => n2914);
   U3792 : AOI221_X1 port map( B1 => n2013, B2 => n6154, C1 => n2014, C2 => 
                           n6186, A => n2915, ZN => n2912);
   U3793 : OAI22_X1 port map( A1 => n5460, A2 => n2016, B1 => n5461, B2 => 
                           n2017, ZN => n2915);
   U3794 : AOI221_X1 port map( B1 => n2018, B2 => n6218, C1 => n2019, C2 => 
                           n6250, A => n2916, ZN => n2911);
   U3795 : OAI222_X1 port map( A1 => n4970, A2 => n2021, B1 => n4938, B2 => 
                           n2022, C1 => n4906, C2 => n419, ZN => n2916);
   U3796 : AOI221_X1 port map( B1 => n2023, B2 => n600, C1 => n2024, C2 => n144
                           , A => n2917, ZN => n2910);
   U3797 : OAI22_X1 port map( A1 => n48, A2 => n2026, B1 => n504, B2 => n2027, 
                           ZN => n2917);
   U3798 : NAND4_X1 port map( A1 => n2918, A2 => n2919, A3 => n2920, A4 => 
                           n2921, ZN => n2890);
   U3799 : AOI221_X1 port map( B1 => n2032, B2 => n5834, C1 => n2033, C2 => 
                           n5866, A => n2922, ZN => n2921);
   U3800 : OAI222_X1 port map( A1 => n4618, A2 => n2035, B1 => n4586, B2 => 
                           n2036, C1 => n4554, C2 => n1577, ZN => n2922);
   U3801 : AOI221_X1 port map( B1 => n2037, B2 => n5898, C1 => n2038, C2 => 
                           n5930, A => n2923, ZN => n2920);
   U3802 : OAI22_X1 port map( A1 => n4682, A2 => n2040, B1 => n4650, B2 => 
                           n2041, ZN => n2923);
   U3803 : AOI221_X1 port map( B1 => n2042, B2 => n5962, C1 => n2043, C2 => 
                           n5994, A => n2924, ZN => n2919);
   U3804 : OAI222_X1 port map( A1 => n4778, A2 => n411, B1 => n4746, B2 => 
                           n2045, C1 => n4714, C2 => n2046, ZN => n2924);
   U3805 : AOI221_X1 port map( B1 => n2047, B2 => n6026, C1 => n2048, C2 => 
                           n6058, A => n2925, ZN => n2918);
   U3806 : OAI22_X1 port map( A1 => n5458, A2 => n2050, B1 => n5459, B2 => 
                           n2051, ZN => n2925);
   U3807 : OAI21_X1 port map( B1 => n1951, B2 => n1536, A => ENABLE, ZN => 
                           n7626);
   U3808 : OAI222_X1 port map( A1 => n2926, A2 => n1948, B1 => n2927, B2 => 
                           n1950, C1 => n1951, C2 => n1473, ZN => n7625);
   U3809 : NOR4_X1 port map( A1 => n2928, A2 => n2929, A3 => n2930, A4 => n2931
                           , ZN => n2927);
   U3810 : NAND4_X1 port map( A1 => n2932, A2 => n2933, A3 => n2934, A4 => 
                           n2935, ZN => n2931);
   U3811 : AOI221_X1 port map( B1 => n1960, B2 => n6409, C1 => n1961, C2 => 
                           n6441, A => n2936, ZN => n2935);
   U3812 : OAI222_X1 port map( A1 => n5257, A2 => n1963, B1 => n5225, B2 => 
                           n1964, C1 => n5193, C2 => n1965, ZN => n2936);
   U3813 : AOI221_X1 port map( B1 => n1966, B2 => n6473, C1 => n1967, C2 => 
                           n6505, A => n2937, ZN => n2934);
   U3814 : OAI22_X1 port map( A1 => n5454, A2 => n1969, B1 => n5455, B2 => 
                           n1970, ZN => n2937);
   U3815 : AOI221_X1 port map( B1 => n1971, B2 => n6537, C1 => n1972, C2 => 
                           n6569, A => n2938, ZN => n2933);
   U3816 : OAI222_X1 port map( A1 => n5353, A2 => n1974, B1 => n5321, B2 => 
                           n1578, C1 => n5289, C2 => n1975, ZN => n2938);
   U3817 : AOI221_X1 port map( B1 => n1976, B2 => n6601, C1 => n1977, C2 => 
                           n6633, A => n2939, ZN => n2932);
   U3818 : OAI22_X1 port map( A1 => n5456, A2 => n1756, B1 => n5457, B2 => 
                           n1980, ZN => n2939);
   U3819 : NAND4_X1 port map( A1 => n2940, A2 => n2941, A3 => n2942, A4 => 
                           n2943, ZN => n2930);
   U3820 : AOI221_X1 port map( B1 => n1985, B2 => n6281, C1 => n1986, C2 => 
                           n6313, A => n2944, ZN => n2943);
   U3821 : OAI222_X1 port map( A1 => n5065, A2 => n1988, B1 => n5033, B2 => 
                           n1989, C1 => n5001, C2 => n416, ZN => n2944);
   U3822 : AOI221_X1 port map( B1 => n1990, B2 => n185, C1 => n1991, C2 => n545
                           , A => n2945, ZN => n2942);
   U3823 : OAI22_X1 port map( A1 => n89, A2 => n1993, B1 => n449, B2 => n1994, 
                           ZN => n2945);
   U3824 : AOI221_X1 port map( B1 => n1995, B2 => n6345, C1 => n1996, C2 => 
                           n6377, A => n2946, ZN => n2941);
   U3825 : OAI222_X1 port map( A1 => n5161, A2 => n1998, B1 => n5129, B2 => 
                           n1999, C1 => n5097, C2 => n417, ZN => n2946);
   U3826 : AOI221_X1 port map( B1 => n2000, B2 => n601, C1 => n2001, C2 => n145
                           , A => n2947, ZN => n2940);
   U3827 : OAI22_X1 port map( A1 => n49, A2 => n412, B1 => n505, B2 => n2003, 
                           ZN => n2947);
   U3828 : NAND4_X1 port map( A1 => n2948, A2 => n2949, A3 => n2950, A4 => 
                           n2951, ZN => n2929);
   U3829 : AOI221_X1 port map( B1 => n2008, B2 => n6089, C1 => n2009, C2 => 
                           n6121, A => n2952, ZN => n2951);
   U3830 : OAI222_X1 port map( A1 => n4873, A2 => n2011, B1 => n4841, B2 => 
                           n2012, C1 => n4809, C2 => n418, ZN => n2952);
   U3831 : AOI221_X1 port map( B1 => n2013, B2 => n6153, C1 => n2014, C2 => 
                           n6185, A => n2953, ZN => n2950);
   U3832 : OAI22_X1 port map( A1 => n5450, A2 => n2016, B1 => n5451, B2 => 
                           n2017, ZN => n2953);
   U3833 : AOI221_X1 port map( B1 => n2018, B2 => n6217, C1 => n2019, C2 => 
                           n6249, A => n2954, ZN => n2949);
   U3834 : OAI222_X1 port map( A1 => n4969, A2 => n2021, B1 => n4937, B2 => 
                           n2022, C1 => n4905, C2 => n419, ZN => n2954);
   U3835 : AOI221_X1 port map( B1 => n2023, B2 => n602, C1 => n2024, C2 => n146
                           , A => n2955, ZN => n2948);
   U3836 : OAI22_X1 port map( A1 => n50, A2 => n2026, B1 => n506, B2 => n2027, 
                           ZN => n2955);
   U3837 : NAND4_X1 port map( A1 => n2956, A2 => n2957, A3 => n2958, A4 => 
                           n2959, ZN => n2928);
   U3838 : AOI221_X1 port map( B1 => n2032, B2 => n5833, C1 => n2033, C2 => 
                           n5865, A => n2960, ZN => n2959);
   U3839 : OAI222_X1 port map( A1 => n4617, A2 => n2035, B1 => n4585, B2 => 
                           n2036, C1 => n4553, C2 => n1577, ZN => n2960);
   U3840 : AOI221_X1 port map( B1 => n2037, B2 => n5897, C1 => n2038, C2 => 
                           n5929, A => n2961, ZN => n2958);
   U3841 : OAI22_X1 port map( A1 => n4681, A2 => n2040, B1 => n4649, B2 => 
                           n2041, ZN => n2961);
   U3842 : AOI221_X1 port map( B1 => n2042, B2 => n5961, C1 => n2043, C2 => 
                           n5993, A => n2962, ZN => n2957);
   U3843 : OAI222_X1 port map( A1 => n4777, A2 => n411, B1 => n4745, B2 => 
                           n2045, C1 => n4713, C2 => n2046, ZN => n2962);
   U3844 : AOI221_X1 port map( B1 => n2047, B2 => n6025, C1 => n2048, C2 => 
                           n6057, A => n2963, ZN => n2956);
   U3845 : OAI22_X1 port map( A1 => n5448, A2 => n2050, B1 => n5449, B2 => 
                           n2051, ZN => n2963);
   U3846 : OAI21_X1 port map( B1 => n1951, B2 => n1537, A => ENABLE, ZN => 
                           n7624);
   U3847 : OAI222_X1 port map( A1 => n2964, A2 => n1948, B1 => n2965, B2 => 
                           n1950, C1 => n1951, C2 => n1474, ZN => n7623);
   U3848 : NOR4_X1 port map( A1 => n2966, A2 => n2967, A3 => n2968, A4 => n2969
                           , ZN => n2965);
   U3849 : NAND4_X1 port map( A1 => n2970, A2 => n2971, A3 => n2972, A4 => 
                           n2973, ZN => n2969);
   U3850 : AOI221_X1 port map( B1 => n1960, B2 => n6408, C1 => n1961, C2 => 
                           n6440, A => n2974, ZN => n2973);
   U3851 : OAI222_X1 port map( A1 => n5256, A2 => n1963, B1 => n5224, B2 => 
                           n1964, C1 => n5192, C2 => n1965, ZN => n2974);
   U3852 : AOI221_X1 port map( B1 => n1966, B2 => n6472, C1 => n1967, C2 => 
                           n6504, A => n2975, ZN => n2972);
   U3853 : OAI22_X1 port map( A1 => n5444, A2 => n1969, B1 => n5445, B2 => 
                           n1970, ZN => n2975);
   U3854 : AOI221_X1 port map( B1 => n1971, B2 => n6536, C1 => n1972, C2 => 
                           n6568, A => n2976, ZN => n2971);
   U3855 : OAI222_X1 port map( A1 => n5352, A2 => n1974, B1 => n5320, B2 => 
                           n1578, C1 => n5288, C2 => n1975, ZN => n2976);
   U3856 : AOI221_X1 port map( B1 => n1976, B2 => n6600, C1 => n1977, C2 => 
                           n6632, A => n2977, ZN => n2970);
   U3857 : OAI22_X1 port map( A1 => n5446, A2 => n1756, B1 => n5447, B2 => 
                           n1980, ZN => n2977);
   U3858 : NAND4_X1 port map( A1 => n2978, A2 => n2979, A3 => n2980, A4 => 
                           n2981, ZN => n2968);
   U3859 : AOI221_X1 port map( B1 => n1985, B2 => n6280, C1 => n1986, C2 => 
                           n6312, A => n2982, ZN => n2981);
   U3860 : OAI222_X1 port map( A1 => n5064, A2 => n1988, B1 => n5032, B2 => 
                           n1989, C1 => n5000, C2 => n416, ZN => n2982);
   U3861 : AOI221_X1 port map( B1 => n1990, B2 => n186, C1 => n1991, C2 => n546
                           , A => n2983, ZN => n2980);
   U3862 : OAI22_X1 port map( A1 => n90, A2 => n1993, B1 => n450, B2 => n1994, 
                           ZN => n2983);
   U3863 : AOI221_X1 port map( B1 => n1995, B2 => n6344, C1 => n1996, C2 => 
                           n6376, A => n2984, ZN => n2979);
   U3864 : OAI222_X1 port map( A1 => n5160, A2 => n1998, B1 => n5128, B2 => 
                           n1999, C1 => n5096, C2 => n417, ZN => n2984);
   U3865 : AOI221_X1 port map( B1 => n2000, B2 => n603, C1 => n2001, C2 => n147
                           , A => n2985, ZN => n2978);
   U3866 : OAI22_X1 port map( A1 => n51, A2 => n412, B1 => n507, B2 => n2003, 
                           ZN => n2985);
   U3867 : NAND4_X1 port map( A1 => n2986, A2 => n2987, A3 => n2988, A4 => 
                           n2989, ZN => n2967);
   U3868 : AOI221_X1 port map( B1 => n2008, B2 => n6088, C1 => n2009, C2 => 
                           n6120, A => n2990, ZN => n2989);
   U3869 : OAI222_X1 port map( A1 => n4872, A2 => n2011, B1 => n4840, B2 => 
                           n2012, C1 => n4808, C2 => n418, ZN => n2990);
   U3870 : AOI221_X1 port map( B1 => n2013, B2 => n6152, C1 => n2014, C2 => 
                           n6184, A => n2991, ZN => n2988);
   U3871 : OAI22_X1 port map( A1 => n5440, A2 => n2016, B1 => n5441, B2 => 
                           n2017, ZN => n2991);
   U3872 : AOI221_X1 port map( B1 => n2018, B2 => n6216, C1 => n2019, C2 => 
                           n6248, A => n2992, ZN => n2987);
   U3873 : OAI222_X1 port map( A1 => n4968, A2 => n2021, B1 => n4936, B2 => 
                           n2022, C1 => n4904, C2 => n419, ZN => n2992);
   U3874 : AOI221_X1 port map( B1 => n2023, B2 => n604, C1 => n2024, C2 => n148
                           , A => n2993, ZN => n2986);
   U3875 : OAI22_X1 port map( A1 => n52, A2 => n2026, B1 => n508, B2 => n2027, 
                           ZN => n2993);
   U3876 : NAND4_X1 port map( A1 => n2994, A2 => n2995, A3 => n2996, A4 => 
                           n2997, ZN => n2966);
   U3877 : AOI221_X1 port map( B1 => n2032, B2 => n5832, C1 => n2033, C2 => 
                           n5864, A => n2998, ZN => n2997);
   U3878 : OAI222_X1 port map( A1 => n4616, A2 => n2035, B1 => n4584, B2 => 
                           n2036, C1 => n4552, C2 => n1577, ZN => n2998);
   U3879 : AOI221_X1 port map( B1 => n2037, B2 => n5896, C1 => n2038, C2 => 
                           n5928, A => n2999, ZN => n2996);
   U3880 : OAI22_X1 port map( A1 => n4680, A2 => n2040, B1 => n4648, B2 => 
                           n2041, ZN => n2999);
   U3881 : AOI221_X1 port map( B1 => n2042, B2 => n5960, C1 => n2043, C2 => 
                           n5992, A => n3000, ZN => n2995);
   U3882 : OAI222_X1 port map( A1 => n4776, A2 => n411, B1 => n4744, B2 => 
                           n2045, C1 => n4712, C2 => n2046, ZN => n3000);
   U3883 : AOI221_X1 port map( B1 => n2047, B2 => n6024, C1 => n2048, C2 => 
                           n6056, A => n3001, ZN => n2994);
   U3884 : OAI22_X1 port map( A1 => n5438, A2 => n2050, B1 => n5439, B2 => 
                           n2051, ZN => n3001);
   U3885 : OAI21_X1 port map( B1 => n1951, B2 => n1538, A => ENABLE, ZN => 
                           n7622);
   U3886 : OAI222_X1 port map( A1 => n3002, A2 => n1948, B1 => n3003, B2 => 
                           n1950, C1 => n1951, C2 => n1475, ZN => n7621);
   U3887 : NOR4_X1 port map( A1 => n3004, A2 => n3005, A3 => n3006, A4 => n3007
                           , ZN => n3003);
   U3888 : NAND4_X1 port map( A1 => n3008, A2 => n3009, A3 => n3010, A4 => 
                           n3011, ZN => n3007);
   U3889 : AOI221_X1 port map( B1 => n1960, B2 => n6407, C1 => n1961, C2 => 
                           n6439, A => n3012, ZN => n3011);
   U3890 : OAI222_X1 port map( A1 => n5255, A2 => n1963, B1 => n5223, B2 => 
                           n1964, C1 => n5191, C2 => n1965, ZN => n3012);
   U3891 : AOI221_X1 port map( B1 => n1966, B2 => n6471, C1 => n1967, C2 => 
                           n6503, A => n3013, ZN => n3010);
   U3892 : OAI22_X1 port map( A1 => n5434, A2 => n1969, B1 => n5435, B2 => 
                           n1970, ZN => n3013);
   U3893 : AOI221_X1 port map( B1 => n1971, B2 => n6535, C1 => n1972, C2 => 
                           n6567, A => n3014, ZN => n3009);
   U3894 : OAI222_X1 port map( A1 => n5351, A2 => n1974, B1 => n5319, B2 => 
                           n1578, C1 => n5287, C2 => n1975, ZN => n3014);
   U3895 : AOI221_X1 port map( B1 => n1976, B2 => n6599, C1 => n1977, C2 => 
                           n6631, A => n3015, ZN => n3008);
   U3896 : OAI22_X1 port map( A1 => n5436, A2 => n1756, B1 => n5437, B2 => 
                           n1980, ZN => n3015);
   U3897 : NAND4_X1 port map( A1 => n3016, A2 => n3017, A3 => n3018, A4 => 
                           n3019, ZN => n3006);
   U3898 : AOI221_X1 port map( B1 => n1985, B2 => n6279, C1 => n1986, C2 => 
                           n6311, A => n3020, ZN => n3019);
   U3899 : OAI222_X1 port map( A1 => n5063, A2 => n1988, B1 => n5031, B2 => 
                           n1989, C1 => n4999, C2 => n416, ZN => n3020);
   U3900 : AOI221_X1 port map( B1 => n1990, B2 => n187, C1 => n1991, C2 => n547
                           , A => n3021, ZN => n3018);
   U3901 : OAI22_X1 port map( A1 => n91, A2 => n1993, B1 => n451, B2 => n1994, 
                           ZN => n3021);
   U3902 : AOI221_X1 port map( B1 => n1995, B2 => n6343, C1 => n1996, C2 => 
                           n6375, A => n3022, ZN => n3017);
   U3903 : OAI222_X1 port map( A1 => n5159, A2 => n1998, B1 => n5127, B2 => 
                           n1999, C1 => n5095, C2 => n417, ZN => n3022);
   U3904 : AOI221_X1 port map( B1 => n2000, B2 => n605, C1 => n2001, C2 => n149
                           , A => n3023, ZN => n3016);
   U3905 : OAI22_X1 port map( A1 => n53, A2 => n412, B1 => n509, B2 => n2003, 
                           ZN => n3023);
   U3906 : NAND4_X1 port map( A1 => n3024, A2 => n3025, A3 => n3026, A4 => 
                           n3027, ZN => n3005);
   U3907 : AOI221_X1 port map( B1 => n2008, B2 => n6087, C1 => n2009, C2 => 
                           n6119, A => n3028, ZN => n3027);
   U3908 : OAI222_X1 port map( A1 => n4871, A2 => n2011, B1 => n4839, B2 => 
                           n2012, C1 => n4807, C2 => n418, ZN => n3028);
   U3909 : AOI221_X1 port map( B1 => n2013, B2 => n6151, C1 => n2014, C2 => 
                           n6183, A => n3029, ZN => n3026);
   U3910 : OAI22_X1 port map( A1 => n5430, A2 => n2016, B1 => n5431, B2 => 
                           n2017, ZN => n3029);
   U3911 : AOI221_X1 port map( B1 => n2018, B2 => n6215, C1 => n2019, C2 => 
                           n6247, A => n3030, ZN => n3025);
   U3912 : OAI222_X1 port map( A1 => n4967, A2 => n2021, B1 => n4935, B2 => 
                           n2022, C1 => n4903, C2 => n419, ZN => n3030);
   U3913 : AOI221_X1 port map( B1 => n2023, B2 => n606, C1 => n2024, C2 => n150
                           , A => n3031, ZN => n3024);
   U3914 : OAI22_X1 port map( A1 => n54, A2 => n2026, B1 => n510, B2 => n2027, 
                           ZN => n3031);
   U3915 : NAND4_X1 port map( A1 => n3032, A2 => n3033, A3 => n3034, A4 => 
                           n3035, ZN => n3004);
   U3916 : AOI221_X1 port map( B1 => n2032, B2 => n5831, C1 => n2033, C2 => 
                           n5863, A => n3036, ZN => n3035);
   U3917 : OAI222_X1 port map( A1 => n4615, A2 => n2035, B1 => n4583, B2 => 
                           n2036, C1 => n4551, C2 => n1577, ZN => n3036);
   U3918 : AOI221_X1 port map( B1 => n2037, B2 => n5895, C1 => n2038, C2 => 
                           n5927, A => n3037, ZN => n3034);
   U3919 : OAI22_X1 port map( A1 => n4679, A2 => n2040, B1 => n4647, B2 => 
                           n2041, ZN => n3037);
   U3920 : AOI221_X1 port map( B1 => n2042, B2 => n5959, C1 => n2043, C2 => 
                           n5991, A => n3038, ZN => n3033);
   U3921 : OAI222_X1 port map( A1 => n4775, A2 => n411, B1 => n4743, B2 => 
                           n2045, C1 => n4711, C2 => n2046, ZN => n3038);
   U3922 : AOI221_X1 port map( B1 => n2047, B2 => n6023, C1 => n2048, C2 => 
                           n6055, A => n3039, ZN => n3032);
   U3923 : OAI22_X1 port map( A1 => n5428, A2 => n2050, B1 => n5429, B2 => 
                           n2051, ZN => n3039);
   U3924 : OAI21_X1 port map( B1 => n1951, B2 => n1539, A => ENABLE, ZN => 
                           n7620);
   U3925 : OAI222_X1 port map( A1 => n3040, A2 => n1948, B1 => n3041, B2 => 
                           n1950, C1 => n1951, C2 => n1476, ZN => n7619);
   U3926 : NOR4_X1 port map( A1 => n3042, A2 => n3043, A3 => n3044, A4 => n3045
                           , ZN => n3041);
   U3927 : NAND4_X1 port map( A1 => n3046, A2 => n3047, A3 => n3048, A4 => 
                           n3049, ZN => n3045);
   U3928 : AOI221_X1 port map( B1 => n1960, B2 => n6406, C1 => n1961, C2 => 
                           n6438, A => n3050, ZN => n3049);
   U3929 : OAI222_X1 port map( A1 => n5254, A2 => n1963, B1 => n5222, B2 => 
                           n1964, C1 => n5190, C2 => n1965, ZN => n3050);
   U3930 : AOI221_X1 port map( B1 => n1966, B2 => n6470, C1 => n1967, C2 => 
                           n6502, A => n3051, ZN => n3048);
   U3931 : OAI22_X1 port map( A1 => n5424, A2 => n1969, B1 => n5425, B2 => 
                           n1970, ZN => n3051);
   U3932 : AOI221_X1 port map( B1 => n1971, B2 => n6534, C1 => n1972, C2 => 
                           n6566, A => n3052, ZN => n3047);
   U3933 : OAI222_X1 port map( A1 => n5350, A2 => n1974, B1 => n5318, B2 => 
                           n1578, C1 => n5286, C2 => n1975, ZN => n3052);
   U3934 : AOI221_X1 port map( B1 => n1976, B2 => n6598, C1 => n1977, C2 => 
                           n6630, A => n3053, ZN => n3046);
   U3935 : OAI22_X1 port map( A1 => n5426, A2 => n1756, B1 => n5427, B2 => 
                           n1980, ZN => n3053);
   U3936 : NAND4_X1 port map( A1 => n3054, A2 => n3055, A3 => n3056, A4 => 
                           n3057, ZN => n3044);
   U3937 : AOI221_X1 port map( B1 => n1985, B2 => n6278, C1 => n1986, C2 => 
                           n6310, A => n3058, ZN => n3057);
   U3938 : OAI222_X1 port map( A1 => n5062, A2 => n1988, B1 => n5030, B2 => 
                           n1989, C1 => n4998, C2 => n416, ZN => n3058);
   U3939 : AOI221_X1 port map( B1 => n1990, B2 => n188, C1 => n1991, C2 => n548
                           , A => n3059, ZN => n3056);
   U3940 : OAI22_X1 port map( A1 => n92, A2 => n1993, B1 => n452, B2 => n1994, 
                           ZN => n3059);
   U3941 : AOI221_X1 port map( B1 => n1995, B2 => n6342, C1 => n1996, C2 => 
                           n6374, A => n3060, ZN => n3055);
   U3942 : OAI222_X1 port map( A1 => n5158, A2 => n1998, B1 => n5126, B2 => 
                           n1999, C1 => n5094, C2 => n417, ZN => n3060);
   U3943 : AOI221_X1 port map( B1 => n2000, B2 => n607, C1 => n2001, C2 => n151
                           , A => n3061, ZN => n3054);
   U3944 : OAI22_X1 port map( A1 => n55, A2 => n412, B1 => n511, B2 => n2003, 
                           ZN => n3061);
   U3945 : NAND4_X1 port map( A1 => n3062, A2 => n3063, A3 => n3064, A4 => 
                           n3065, ZN => n3043);
   U3946 : AOI221_X1 port map( B1 => n2008, B2 => n6086, C1 => n2009, C2 => 
                           n6118, A => n3066, ZN => n3065);
   U3947 : OAI222_X1 port map( A1 => n4870, A2 => n2011, B1 => n4838, B2 => 
                           n2012, C1 => n4806, C2 => n418, ZN => n3066);
   U3948 : AOI221_X1 port map( B1 => n2013, B2 => n6150, C1 => n2014, C2 => 
                           n6182, A => n3067, ZN => n3064);
   U3949 : OAI22_X1 port map( A1 => n5420, A2 => n2016, B1 => n5421, B2 => 
                           n2017, ZN => n3067);
   U3950 : AOI221_X1 port map( B1 => n2018, B2 => n6214, C1 => n2019, C2 => 
                           n6246, A => n3068, ZN => n3063);
   U3951 : OAI222_X1 port map( A1 => n4966, A2 => n2021, B1 => n4934, B2 => 
                           n2022, C1 => n4902, C2 => n419, ZN => n3068);
   U3952 : AOI221_X1 port map( B1 => n2023, B2 => n608, C1 => n2024, C2 => n152
                           , A => n3069, ZN => n3062);
   U3953 : OAI22_X1 port map( A1 => n56, A2 => n2026, B1 => n512, B2 => n2027, 
                           ZN => n3069);
   U3954 : NAND4_X1 port map( A1 => n3070, A2 => n3071, A3 => n3072, A4 => 
                           n3073, ZN => n3042);
   U3955 : AOI221_X1 port map( B1 => n2032, B2 => n5830, C1 => n2033, C2 => 
                           n5862, A => n3074, ZN => n3073);
   U3956 : OAI222_X1 port map( A1 => n4614, A2 => n2035, B1 => n4582, B2 => 
                           n2036, C1 => n4550, C2 => n1577, ZN => n3074);
   U3957 : AOI221_X1 port map( B1 => n2037, B2 => n5894, C1 => n2038, C2 => 
                           n5926, A => n3075, ZN => n3072);
   U3958 : OAI22_X1 port map( A1 => n4678, A2 => n2040, B1 => n4646, B2 => 
                           n2041, ZN => n3075);
   U3959 : AOI221_X1 port map( B1 => n2042, B2 => n5958, C1 => n2043, C2 => 
                           n5990, A => n3076, ZN => n3071);
   U3960 : OAI222_X1 port map( A1 => n4774, A2 => n411, B1 => n4742, B2 => 
                           n2045, C1 => n4710, C2 => n2046, ZN => n3076);
   U3961 : AOI221_X1 port map( B1 => n2047, B2 => n6022, C1 => n2048, C2 => 
                           n6054, A => n3077, ZN => n3070);
   U3962 : OAI22_X1 port map( A1 => n5418, A2 => n2050, B1 => n5419, B2 => 
                           n2051, ZN => n3077);
   U3963 : OAI21_X1 port map( B1 => n1951, B2 => n1540, A => ENABLE, ZN => 
                           n7618);
   U3964 : OAI222_X1 port map( A1 => n3078, A2 => n1948, B1 => n3079, B2 => 
                           n1950, C1 => n1951, C2 => n1477, ZN => n7617);
   U3965 : NOR4_X1 port map( A1 => n3080, A2 => n3081, A3 => n3082, A4 => n3083
                           , ZN => n3079);
   U3966 : NAND4_X1 port map( A1 => n3084, A2 => n3085, A3 => n3086, A4 => 
                           n3087, ZN => n3083);
   U3967 : AOI221_X1 port map( B1 => n1960, B2 => n6405, C1 => n1961, C2 => 
                           n6437, A => n3088, ZN => n3087);
   U3968 : OAI222_X1 port map( A1 => n5253, A2 => n1963, B1 => n5221, B2 => 
                           n1964, C1 => n5189, C2 => n1965, ZN => n3088);
   U3969 : AOI221_X1 port map( B1 => n1966, B2 => n6469, C1 => n1967, C2 => 
                           n6501, A => n3089, ZN => n3086);
   U3970 : OAI22_X1 port map( A1 => n5414, A2 => n1969, B1 => n5415, B2 => 
                           n1970, ZN => n3089);
   U3971 : AOI221_X1 port map( B1 => n1971, B2 => n6533, C1 => n1972, C2 => 
                           n6565, A => n3090, ZN => n3085);
   U3972 : OAI222_X1 port map( A1 => n5349, A2 => n1974, B1 => n5317, B2 => 
                           n1578, C1 => n5285, C2 => n1975, ZN => n3090);
   U3973 : AOI221_X1 port map( B1 => n1976, B2 => n6597, C1 => n1977, C2 => 
                           n6629, A => n3091, ZN => n3084);
   U3974 : OAI22_X1 port map( A1 => n5416, A2 => n1756, B1 => n5417, B2 => 
                           n1980, ZN => n3091);
   U3975 : NAND4_X1 port map( A1 => n3092, A2 => n3093, A3 => n3094, A4 => 
                           n3095, ZN => n3082);
   U3976 : AOI221_X1 port map( B1 => n1985, B2 => n6277, C1 => n1986, C2 => 
                           n6309, A => n3096, ZN => n3095);
   U3977 : OAI222_X1 port map( A1 => n5061, A2 => n1988, B1 => n5029, B2 => 
                           n1989, C1 => n4997, C2 => n416, ZN => n3096);
   U3978 : AOI221_X1 port map( B1 => n1990, B2 => n189, C1 => n1991, C2 => n549
                           , A => n3097, ZN => n3094);
   U3979 : OAI22_X1 port map( A1 => n93, A2 => n1993, B1 => n453, B2 => n1994, 
                           ZN => n3097);
   U3980 : AOI221_X1 port map( B1 => n1995, B2 => n6341, C1 => n1996, C2 => 
                           n6373, A => n3098, ZN => n3093);
   U3981 : OAI222_X1 port map( A1 => n5157, A2 => n1998, B1 => n5125, B2 => 
                           n1999, C1 => n5093, C2 => n417, ZN => n3098);
   U3982 : AOI221_X1 port map( B1 => n2000, B2 => n609, C1 => n2001, C2 => n153
                           , A => n3099, ZN => n3092);
   U3983 : OAI22_X1 port map( A1 => n57, A2 => n412, B1 => n513, B2 => n2003, 
                           ZN => n3099);
   U3984 : NAND4_X1 port map( A1 => n3100, A2 => n3101, A3 => n3102, A4 => 
                           n3103, ZN => n3081);
   U3985 : AOI221_X1 port map( B1 => n2008, B2 => n6085, C1 => n2009, C2 => 
                           n6117, A => n3104, ZN => n3103);
   U3986 : OAI222_X1 port map( A1 => n4869, A2 => n2011, B1 => n4837, B2 => 
                           n2012, C1 => n4805, C2 => n418, ZN => n3104);
   U3987 : AOI221_X1 port map( B1 => n2013, B2 => n6149, C1 => n2014, C2 => 
                           n6181, A => n3105, ZN => n3102);
   U3988 : OAI22_X1 port map( A1 => n5410, A2 => n2016, B1 => n5411, B2 => 
                           n2017, ZN => n3105);
   U3989 : AOI221_X1 port map( B1 => n2018, B2 => n6213, C1 => n2019, C2 => 
                           n6245, A => n3106, ZN => n3101);
   U3990 : OAI222_X1 port map( A1 => n4965, A2 => n2021, B1 => n4933, B2 => 
                           n2022, C1 => n4901, C2 => n419, ZN => n3106);
   U3991 : AOI221_X1 port map( B1 => n2023, B2 => n610, C1 => n2024, C2 => n154
                           , A => n3107, ZN => n3100);
   U3992 : OAI22_X1 port map( A1 => n58, A2 => n2026, B1 => n514, B2 => n2027, 
                           ZN => n3107);
   U3993 : NAND4_X1 port map( A1 => n3108, A2 => n3109, A3 => n3110, A4 => 
                           n3111, ZN => n3080);
   U3994 : AOI221_X1 port map( B1 => n2032, B2 => n5829, C1 => n2033, C2 => 
                           n5861, A => n3112, ZN => n3111);
   U3995 : OAI222_X1 port map( A1 => n4613, A2 => n2035, B1 => n4581, B2 => 
                           n2036, C1 => n4549, C2 => n1577, ZN => n3112);
   U3996 : AOI221_X1 port map( B1 => n2037, B2 => n5893, C1 => n2038, C2 => 
                           n5925, A => n3113, ZN => n3110);
   U3997 : OAI22_X1 port map( A1 => n4677, A2 => n2040, B1 => n4645, B2 => 
                           n2041, ZN => n3113);
   U3998 : AOI221_X1 port map( B1 => n2042, B2 => n5957, C1 => n2043, C2 => 
                           n5989, A => n3114, ZN => n3109);
   U3999 : OAI222_X1 port map( A1 => n4773, A2 => n411, B1 => n4741, B2 => 
                           n2045, C1 => n4709, C2 => n2046, ZN => n3114);
   U4000 : AOI221_X1 port map( B1 => n2047, B2 => n6021, C1 => n2048, C2 => 
                           n6053, A => n3115, ZN => n3108);
   U4001 : OAI22_X1 port map( A1 => n5408, A2 => n2050, B1 => n5409, B2 => 
                           n2051, ZN => n3115);
   U4002 : OAI21_X1 port map( B1 => n1951, B2 => n1541, A => ENABLE, ZN => 
                           n7616);
   U4003 : OAI222_X1 port map( A1 => n3116, A2 => n1948, B1 => n3117, B2 => 
                           n1950, C1 => n1951, C2 => n1478, ZN => n7615);
   U4004 : NOR4_X1 port map( A1 => n3118, A2 => n3119, A3 => n3120, A4 => n3121
                           , ZN => n3117);
   U4005 : NAND4_X1 port map( A1 => n3122, A2 => n3123, A3 => n3124, A4 => 
                           n3125, ZN => n3121);
   U4006 : AOI221_X1 port map( B1 => n1960, B2 => n6404, C1 => n1961, C2 => 
                           n6436, A => n3126, ZN => n3125);
   U4007 : OAI222_X1 port map( A1 => n5252, A2 => n1963, B1 => n5220, B2 => 
                           n1964, C1 => n5188, C2 => n1965, ZN => n3126);
   U4008 : AOI221_X1 port map( B1 => n1966, B2 => n6468, C1 => n1967, C2 => 
                           n6500, A => n3127, ZN => n3124);
   U4009 : OAI22_X1 port map( A1 => n5404, A2 => n1969, B1 => n5405, B2 => 
                           n1970, ZN => n3127);
   U4010 : AOI221_X1 port map( B1 => n1971, B2 => n6532, C1 => n1972, C2 => 
                           n6564, A => n3128, ZN => n3123);
   U4011 : OAI222_X1 port map( A1 => n5348, A2 => n1974, B1 => n5316, B2 => 
                           n1578, C1 => n5284, C2 => n1975, ZN => n3128);
   U4012 : AOI221_X1 port map( B1 => n1976, B2 => n6596, C1 => n1977, C2 => 
                           n6628, A => n3129, ZN => n3122);
   U4013 : OAI22_X1 port map( A1 => n5406, A2 => n1756, B1 => n5407, B2 => 
                           n1980, ZN => n3129);
   U4014 : NAND4_X1 port map( A1 => n3130, A2 => n3131, A3 => n3132, A4 => 
                           n3133, ZN => n3120);
   U4015 : AOI221_X1 port map( B1 => n1985, B2 => n6276, C1 => n1986, C2 => 
                           n6308, A => n3134, ZN => n3133);
   U4016 : OAI222_X1 port map( A1 => n5060, A2 => n1988, B1 => n5028, B2 => 
                           n1989, C1 => n4996, C2 => n416, ZN => n3134);
   U4017 : AOI221_X1 port map( B1 => n1990, B2 => n190, C1 => n1991, C2 => n550
                           , A => n3135, ZN => n3132);
   U4018 : OAI22_X1 port map( A1 => n94, A2 => n1993, B1 => n454, B2 => n1994, 
                           ZN => n3135);
   U4019 : AOI221_X1 port map( B1 => n1995, B2 => n6340, C1 => n1996, C2 => 
                           n6372, A => n3136, ZN => n3131);
   U4020 : OAI222_X1 port map( A1 => n5156, A2 => n1998, B1 => n5124, B2 => 
                           n1999, C1 => n5092, C2 => n417, ZN => n3136);
   U4021 : AOI221_X1 port map( B1 => n2000, B2 => n611, C1 => n2001, C2 => n155
                           , A => n3137, ZN => n3130);
   U4022 : OAI22_X1 port map( A1 => n59, A2 => n412, B1 => n515, B2 => n2003, 
                           ZN => n3137);
   U4023 : NAND4_X1 port map( A1 => n3138, A2 => n3139, A3 => n3140, A4 => 
                           n3141, ZN => n3119);
   U4024 : AOI221_X1 port map( B1 => n2008, B2 => n6084, C1 => n2009, C2 => 
                           n6116, A => n3142, ZN => n3141);
   U4025 : OAI222_X1 port map( A1 => n4868, A2 => n2011, B1 => n4836, B2 => 
                           n2012, C1 => n4804, C2 => n418, ZN => n3142);
   U4026 : AOI221_X1 port map( B1 => n2013, B2 => n6148, C1 => n2014, C2 => 
                           n6180, A => n3143, ZN => n3140);
   U4027 : OAI22_X1 port map( A1 => n5400, A2 => n2016, B1 => n5401, B2 => 
                           n2017, ZN => n3143);
   U4028 : AOI221_X1 port map( B1 => n2018, B2 => n6212, C1 => n2019, C2 => 
                           n6244, A => n3144, ZN => n3139);
   U4029 : OAI222_X1 port map( A1 => n4964, A2 => n2021, B1 => n4932, B2 => 
                           n2022, C1 => n4900, C2 => n419, ZN => n3144);
   U4030 : AOI221_X1 port map( B1 => n2023, B2 => n612, C1 => n2024, C2 => n156
                           , A => n3145, ZN => n3138);
   U4031 : OAI22_X1 port map( A1 => n60, A2 => n2026, B1 => n516, B2 => n2027, 
                           ZN => n3145);
   U4032 : NAND4_X1 port map( A1 => n3146, A2 => n3147, A3 => n3148, A4 => 
                           n3149, ZN => n3118);
   U4033 : AOI221_X1 port map( B1 => n2032, B2 => n5828, C1 => n2033, C2 => 
                           n5860, A => n3150, ZN => n3149);
   U4034 : OAI222_X1 port map( A1 => n4612, A2 => n2035, B1 => n4580, B2 => 
                           n2036, C1 => n4548, C2 => n1577, ZN => n3150);
   U4035 : AOI221_X1 port map( B1 => n2037, B2 => n5892, C1 => n2038, C2 => 
                           n5924, A => n3151, ZN => n3148);
   U4036 : OAI22_X1 port map( A1 => n4676, A2 => n2040, B1 => n4644, B2 => 
                           n2041, ZN => n3151);
   U4037 : AOI221_X1 port map( B1 => n2042, B2 => n5956, C1 => n2043, C2 => 
                           n5988, A => n3152, ZN => n3147);
   U4038 : OAI222_X1 port map( A1 => n4772, A2 => n411, B1 => n4740, B2 => 
                           n2045, C1 => n4708, C2 => n2046, ZN => n3152);
   U4039 : AOI221_X1 port map( B1 => n2047, B2 => n6020, C1 => n2048, C2 => 
                           n6052, A => n3153, ZN => n3146);
   U4040 : OAI22_X1 port map( A1 => n5398, A2 => n2050, B1 => n5399, B2 => 
                           n2051, ZN => n3153);
   U4041 : OAI21_X1 port map( B1 => n1951, B2 => n1542, A => ENABLE, ZN => 
                           n7614);
   U4042 : OAI222_X1 port map( A1 => n3154, A2 => n1948, B1 => n3155, B2 => 
                           n1950, C1 => n1951, C2 => n1479, ZN => n7613);
   U4043 : NOR4_X1 port map( A1 => n3156, A2 => n3157, A3 => n3158, A4 => n3159
                           , ZN => n3155);
   U4044 : NAND4_X1 port map( A1 => n3160, A2 => n3161, A3 => n3162, A4 => 
                           n3163, ZN => n3159);
   U4045 : AOI221_X1 port map( B1 => n1960, B2 => n6403, C1 => n1961, C2 => 
                           n6435, A => n3164, ZN => n3163);
   U4046 : OAI222_X1 port map( A1 => n5251, A2 => n1963, B1 => n5219, B2 => 
                           n1964, C1 => n5187, C2 => n1965, ZN => n3164);
   U4047 : AOI221_X1 port map( B1 => n1966, B2 => n6467, C1 => n1967, C2 => 
                           n6499, A => n3165, ZN => n3162);
   U4048 : OAI22_X1 port map( A1 => n5394, A2 => n1969, B1 => n5395, B2 => 
                           n1970, ZN => n3165);
   U4049 : AOI221_X1 port map( B1 => n1971, B2 => n6531, C1 => n1972, C2 => 
                           n6563, A => n3166, ZN => n3161);
   U4050 : OAI222_X1 port map( A1 => n5347, A2 => n1974, B1 => n5315, B2 => 
                           n1578, C1 => n5283, C2 => n1975, ZN => n3166);
   U4051 : AOI221_X1 port map( B1 => n1976, B2 => n6595, C1 => n1977, C2 => 
                           n6627, A => n3167, ZN => n3160);
   U4052 : OAI22_X1 port map( A1 => n5396, A2 => n1756, B1 => n5397, B2 => 
                           n1980, ZN => n3167);
   U4053 : NAND4_X1 port map( A1 => n3168, A2 => n3169, A3 => n3170, A4 => 
                           n3171, ZN => n3158);
   U4054 : AOI221_X1 port map( B1 => n1985, B2 => n6275, C1 => n1986, C2 => 
                           n6307, A => n3172, ZN => n3171);
   U4055 : OAI222_X1 port map( A1 => n5059, A2 => n1988, B1 => n5027, B2 => 
                           n1989, C1 => n4995, C2 => n416, ZN => n3172);
   U4056 : AOI221_X1 port map( B1 => n1990, B2 => n191, C1 => n1991, C2 => n551
                           , A => n3173, ZN => n3170);
   U4057 : OAI22_X1 port map( A1 => n95, A2 => n1993, B1 => n455, B2 => n1994, 
                           ZN => n3173);
   U4058 : AOI221_X1 port map( B1 => n1995, B2 => n6339, C1 => n1996, C2 => 
                           n6371, A => n3174, ZN => n3169);
   U4059 : OAI222_X1 port map( A1 => n5155, A2 => n1998, B1 => n5123, B2 => 
                           n1999, C1 => n5091, C2 => n417, ZN => n3174);
   U4060 : AOI221_X1 port map( B1 => n2000, B2 => n613, C1 => n2001, C2 => n157
                           , A => n3175, ZN => n3168);
   U4061 : OAI22_X1 port map( A1 => n61, A2 => n412, B1 => n517, B2 => n2003, 
                           ZN => n3175);
   U4062 : NAND4_X1 port map( A1 => n3176, A2 => n3177, A3 => n3178, A4 => 
                           n3179, ZN => n3157);
   U4063 : AOI221_X1 port map( B1 => n2008, B2 => n6083, C1 => n2009, C2 => 
                           n6115, A => n3180, ZN => n3179);
   U4064 : OAI222_X1 port map( A1 => n4867, A2 => n2011, B1 => n4835, B2 => 
                           n2012, C1 => n4803, C2 => n418, ZN => n3180);
   U4065 : AOI221_X1 port map( B1 => n2013, B2 => n6147, C1 => n2014, C2 => 
                           n6179, A => n3181, ZN => n3178);
   U4066 : OAI22_X1 port map( A1 => n5390, A2 => n2016, B1 => n5391, B2 => 
                           n2017, ZN => n3181);
   U4067 : AOI221_X1 port map( B1 => n2018, B2 => n6211, C1 => n2019, C2 => 
                           n6243, A => n3182, ZN => n3177);
   U4068 : OAI222_X1 port map( A1 => n4963, A2 => n2021, B1 => n4931, B2 => 
                           n2022, C1 => n4899, C2 => n419, ZN => n3182);
   U4069 : AOI221_X1 port map( B1 => n2023, B2 => n614, C1 => n2024, C2 => n158
                           , A => n3183, ZN => n3176);
   U4070 : OAI22_X1 port map( A1 => n62, A2 => n2026, B1 => n518, B2 => n2027, 
                           ZN => n3183);
   U4071 : NAND4_X1 port map( A1 => n3184, A2 => n3185, A3 => n3186, A4 => 
                           n3187, ZN => n3156);
   U4072 : AOI221_X1 port map( B1 => n2032, B2 => n5827, C1 => n2033, C2 => 
                           n5859, A => n3188, ZN => n3187);
   U4073 : OAI222_X1 port map( A1 => n4611, A2 => n2035, B1 => n4579, B2 => 
                           n2036, C1 => n4547, C2 => n1577, ZN => n3188);
   U4074 : AOI221_X1 port map( B1 => n2037, B2 => n5891, C1 => n2038, C2 => 
                           n5923, A => n3189, ZN => n3186);
   U4075 : OAI22_X1 port map( A1 => n4675, A2 => n2040, B1 => n4643, B2 => 
                           n2041, ZN => n3189);
   U4076 : AOI221_X1 port map( B1 => n2042, B2 => n5955, C1 => n2043, C2 => 
                           n5987, A => n3190, ZN => n3185);
   U4077 : OAI222_X1 port map( A1 => n4771, A2 => n411, B1 => n4739, B2 => 
                           n2045, C1 => n4707, C2 => n2046, ZN => n3190);
   U4078 : AOI221_X1 port map( B1 => n2047, B2 => n6019, C1 => n2048, C2 => 
                           n6051, A => n3191, ZN => n3184);
   U4079 : OAI22_X1 port map( A1 => n5388, A2 => n2050, B1 => n5389, B2 => 
                           n2051, ZN => n3191);
   U4080 : OAI21_X1 port map( B1 => n1951, B2 => n1543, A => ENABLE, ZN => 
                           n7612);
   U4081 : OAI222_X1 port map( A1 => n3192, A2 => n1948, B1 => n3193, B2 => 
                           n1950, C1 => n1951, C2 => n1480, ZN => n7611);
   U4082 : NOR4_X1 port map( A1 => n3194, A2 => n3195, A3 => n3196, A4 => n3197
                           , ZN => n3193);
   U4083 : NAND4_X1 port map( A1 => n3198, A2 => n3199, A3 => n3200, A4 => 
                           n3201, ZN => n3197);
   U4084 : AOI221_X1 port map( B1 => n1960, B2 => n6402, C1 => n1961, C2 => 
                           n6434, A => n3202, ZN => n3201);
   U4085 : OAI222_X1 port map( A1 => n5250, A2 => n1963, B1 => n5218, B2 => 
                           n1964, C1 => n5186, C2 => n1965, ZN => n3202);
   U4086 : AOI221_X1 port map( B1 => n1966, B2 => n6466, C1 => n1967, C2 => 
                           n6498, A => n3210, ZN => n3200);
   U4087 : OAI22_X1 port map( A1 => n5384, A2 => n1969, B1 => n5385, B2 => 
                           n1970, ZN => n3210);
   U4088 : AOI221_X1 port map( B1 => n1971, B2 => n6530, C1 => n1972, C2 => 
                           n6562, A => n3214, ZN => n3199);
   U4089 : OAI222_X1 port map( A1 => n5346, A2 => n1974, B1 => n5314, B2 => 
                           n1578, C1 => n5282, C2 => n1975, ZN => n3214);
   U4090 : AOI221_X1 port map( B1 => n1976, B2 => n6594, C1 => n1977, C2 => 
                           n6626, A => n3217, ZN => n3198);
   U4091 : OAI22_X1 port map( A1 => n5386, A2 => n1756, B1 => n5387, B2 => 
                           n1980, ZN => n3217);
   U4092 : NAND4_X1 port map( A1 => n3218, A2 => n3219, A3 => n3220, A4 => 
                           n3221, ZN => n3196);
   U4093 : AOI221_X1 port map( B1 => n1985, B2 => n6274, C1 => n1986, C2 => 
                           n6306, A => n3222, ZN => n3221);
   U4094 : OAI222_X1 port map( A1 => n5058, A2 => n1988, B1 => n5026, B2 => 
                           n1989, C1 => n4994, C2 => n416, ZN => n3222);
   U4095 : AOI221_X1 port map( B1 => n1990, B2 => n192, C1 => n1991, C2 => n552
                           , A => n3225, ZN => n3220);
   U4096 : OAI22_X1 port map( A1 => n96, A2 => n1993, B1 => n456, B2 => n1994, 
                           ZN => n3225);
   U4097 : AOI221_X1 port map( B1 => n1995, B2 => n6338, C1 => n1996, C2 => 
                           n6370, A => n3226, ZN => n3219);
   U4098 : OAI222_X1 port map( A1 => n5154, A2 => n1998, B1 => n5122, B2 => 
                           n1999, C1 => n5090, C2 => n417, ZN => n3226);
   U4099 : AOI221_X1 port map( B1 => n2000, B2 => n615, C1 => n2001, C2 => n159
                           , A => n3228, ZN => n3218);
   U4100 : OAI22_X1 port map( A1 => n63, A2 => n412, B1 => n519, B2 => n2003, 
                           ZN => n3228);
   U4101 : NAND4_X1 port map( A1 => n3229, A2 => n3230, A3 => n3231, A4 => 
                           n3232, ZN => n3195);
   U4102 : AOI221_X1 port map( B1 => n2008, B2 => n6082, C1 => n2009, C2 => 
                           n6114, A => n3233, ZN => n3232);
   U4103 : OAI222_X1 port map( A1 => n4866, A2 => n2011, B1 => n4834, B2 => 
                           n2012, C1 => n4802, C2 => n418, ZN => n3233);
   U4104 : AOI221_X1 port map( B1 => n2013, B2 => n6146, C1 => n2014, C2 => 
                           n6178, A => n3235, ZN => n3231);
   U4105 : OAI22_X1 port map( A1 => n5380, A2 => n2016, B1 => n5381, B2 => 
                           n2017, ZN => n3235);
   U4106 : AOI221_X1 port map( B1 => n2018, B2 => n6210, C1 => n2019, C2 => 
                           n6242, A => n3237, ZN => n3230);
   U4107 : OAI222_X1 port map( A1 => n4962, A2 => n2021, B1 => n4930, B2 => 
                           n2022, C1 => n4898, C2 => n419, ZN => n3237);
   U4108 : AND2_X1 port map( A1 => n3236, A2 => n3204, ZN => n2018);
   U4109 : AOI221_X1 port map( B1 => n2023, B2 => n616, C1 => n2024, C2 => n160
                           , A => n3239, ZN => n3229);
   U4110 : OAI22_X1 port map( A1 => n64, A2 => n2026, B1 => n520, B2 => n2027, 
                           ZN => n3239);
   U4111 : NAND4_X1 port map( A1 => n3240, A2 => n3241, A3 => n3242, A4 => 
                           n3243, ZN => n3194);
   U4112 : AOI221_X1 port map( B1 => n2032, B2 => n5826, C1 => n2033, C2 => 
                           n5858, A => n3244, ZN => n3243);
   U4113 : OAI222_X1 port map( A1 => n4610, A2 => n2035, B1 => n4578, B2 => 
                           n2036, C1 => n4546, C2 => n1577, ZN => n3244);
   U4114 : AOI221_X1 port map( B1 => n2037, B2 => n5890, C1 => n2038, C2 => 
                           n5922, A => n3245, ZN => n3242);
   U4115 : OAI22_X1 port map( A1 => n4674, A2 => n2040, B1 => n4642, B2 => 
                           n2041, ZN => n3245);
   U4116 : AOI221_X1 port map( B1 => n2042, B2 => n5954, C1 => n2043, C2 => 
                           n5986, A => n3247, ZN => n3241);
   U4117 : OAI222_X1 port map( A1 => n4770, A2 => n411, B1 => n4738, B2 => 
                           n2045, C1 => n4706, C2 => n2046, ZN => n3247);
   U4118 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n3250, 
                           ZN => n3213);
   U4119 : AND2_X1 port map( A1 => n3246, A2 => n3212, ZN => n2042);
   U4120 : AOI221_X1 port map( B1 => n2047, B2 => n6018, C1 => n2048, C2 => 
                           n6050, A => n3251, ZN => n3240);
   U4121 : OAI22_X1 port map( A1 => n5378, A2 => n2050, B1 => n5379, B2 => 
                           n2051, ZN => n3251);
   U4122 : NOR3_X1 port map( A1 => n3250, A2 => ADD_RD1(0), A3 => n3249, ZN => 
                           n3209);
   U4123 : INV_X1 port map( A => ADD_RD1(2), ZN => n3249);
   U4124 : INV_X1 port map( A => ADD_RD1(1), ZN => n3250);
   U4125 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n3205);
   U4126 : AND2_X1 port map( A1 => n3246, A2 => n3204, ZN => n2047);
   U4127 : INV_X1 port map( A => ADD_RD1(0), ZN => n3248);
   U4128 : INV_X1 port map( A => ADD_RD1(5), ZN => n3238);
   U4129 : INV_X1 port map( A => ADD_RD1(3), ZN => n3215);
   U4130 : INV_X1 port map( A => ADD_RD1(4), ZN => n3227);
   U4131 : NOR4_X1 port map( A1 => n3256, A2 => n3257, A3 => n3258, A4 => n3259
                           , ZN => n3255);
   U4132 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD1(6), Z => n3259);
   U4133 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD1(5), Z => n3258);
   U4134 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD1(4), Z => n3257);
   U4135 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD1(3), Z => n3256);
   U4136 : NOR3_X1 port map( A1 => n3260, A2 => n3261, A3 => n3262, ZN => n3254
                           );
   U4137 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD1(0), Z => n3260);
   U4138 : XOR2_X1 port map( A => n1943, B => ADD_RD1(1), Z => n3253);
   U4139 : XOR2_X1 port map( A => n1915, B => ADD_RD1(2), Z => n3252);
   U4140 : OAI21_X1 port map( B1 => n1951, B2 => n1544, A => ENABLE, ZN => 
                           n7610);
   U4141 : INV_X1 port map( A => RD1, ZN => n3262);
   U4142 : OAI222_X1 port map( A1 => n1947, A2 => n3263, B1 => n3264, B2 => 
                           n3265, C1 => n3266, C2 => n1481, ZN => n7609);
   U4143 : NOR4_X1 port map( A1 => n3267, A2 => n3268, A3 => n3269, A4 => n3270
                           , ZN => n3264);
   U4144 : NAND4_X1 port map( A1 => n3271, A2 => n3272, A3 => n3273, A4 => 
                           n3274, ZN => n3270);
   U4145 : AOI221_X1 port map( B1 => n1748, B2 => n6433, C1 => n3276, C2 => 
                           n6465, A => n3277, ZN => n3274);
   U4146 : OAI222_X1 port map( A1 => n5281, A2 => n3278, B1 => n5249, B2 => 
                           n3279, C1 => n5217, C2 => n421, ZN => n3277);
   U4147 : AOI221_X1 port map( B1 => n3280, B2 => n713, C1 => n3281, C2 => n289
                           , A => n3282, ZN => n3273);
   U4148 : OAI22_X1 port map( A1 => n193, A2 => n413, B1 => n617, B2 => n3283, 
                           ZN => n3282);
   U4149 : AOI221_X1 port map( B1 => n1754, B2 => n6561, C1 => n3285, C2 => 
                           n6593, A => n3286, ZN => n3272);
   U4150 : OAI222_X1 port map( A1 => n5377, A2 => n3287, B1 => n5345, B2 => 
                           n1579, C1 => n5313, C2 => n3288, ZN => n3286);
   U4151 : AOI221_X1 port map( B1 => n3289, B2 => n714, C1 => n3290, C2 => n290
                           , A => n3291, ZN => n3271);
   U4152 : OAI22_X1 port map( A1 => n194, A2 => n414, B1 => n618, B2 => n3292, 
                           ZN => n3291);
   U4153 : NAND4_X1 port map( A1 => n3293, A2 => n3294, A3 => n3295, A4 => 
                           n3296, ZN => n3269);
   U4154 : AOI221_X1 port map( B1 => n3297, B2 => n6305, C1 => n3298, C2 => 
                           n6337, A => n3299, ZN => n3296);
   U4155 : OAI222_X1 port map( A1 => n5089, A2 => n3300, B1 => n5057, B2 => 
                           n3301, C1 => n5025, C2 => n3302, ZN => n3299);
   U4156 : AOI221_X1 port map( B1 => n3303, B2 => n521, C1 => n3304, C2 => n161
                           , A => n3305, ZN => n3295);
   U4157 : OAI22_X1 port map( A1 => n425, A2 => n3306, B1 => n65, B2 => n3307, 
                           ZN => n3305);
   U4158 : AOI221_X1 port map( B1 => n3308, B2 => n6369, C1 => n3309, C2 => 
                           n6401, A => n3310, ZN => n3294);
   U4159 : OAI222_X1 port map( A1 => n5185, A2 => n3311, B1 => n5153, B2 => 
                           n3312, C1 => n5121, C2 => n422, ZN => n3310);
   U4160 : AOI221_X1 port map( B1 => n3313, B2 => n553, C1 => n3314, C2 => n97,
                           A => n3315, ZN => n3293);
   U4161 : OAI22_X1 port map( A1 => n1, A2 => n415, B1 => n457, B2 => n3316, ZN
                           => n3315);
   U4162 : NAND4_X1 port map( A1 => n3317, A2 => n3318, A3 => n3319, A4 => 
                           n3320, ZN => n3268);
   U4163 : AOI221_X1 port map( B1 => n3321, B2 => n6113, C1 => n3322, C2 => 
                           n6145, A => n3323, ZN => n3320);
   U4164 : OAI222_X1 port map( A1 => n4897, A2 => n3324, B1 => n4865, B2 => 
                           n3325, C1 => n4833, C2 => n423, ZN => n3323);
   U4165 : AOI221_X1 port map( B1 => n3326, B2 => n715, C1 => n3327, C2 => n291
                           , A => n3328, ZN => n3319);
   U4166 : OAI22_X1 port map( A1 => n195, A2 => n3329, B1 => n619, B2 => n3330,
                           ZN => n3328);
   U4167 : AOI221_X1 port map( B1 => n3331, B2 => n6241, C1 => n3332, C2 => 
                           n6273, A => n3333, ZN => n3318);
   U4168 : OAI222_X1 port map( A1 => n4993, A2 => n3334, B1 => n4961, B2 => 
                           n3335, C1 => n4929, C2 => n3336, ZN => n3333);
   U4169 : AOI221_X1 port map( B1 => n3337, B2 => n554, C1 => n3338, C2 => n98,
                           A => n3339, ZN => n3317);
   U4170 : OAI22_X1 port map( A1 => n2, A2 => n3340, B1 => n458, B2 => n3341, 
                           ZN => n3339);
   U4171 : NAND4_X1 port map( A1 => n3342, A2 => n3343, A3 => n3344, A4 => 
                           n3345, ZN => n3267);
   U4172 : AOI221_X1 port map( B1 => n3346, B2 => n5857, C1 => n3347, C2 => 
                           n5889, A => n3348, ZN => n3345);
   U4173 : OAI222_X1 port map( A1 => n4641, A2 => n3349, B1 => n4609, B2 => 
                           n3350, C1 => n4577, C2 => n3351, ZN => n3348);
   U4174 : AOI221_X1 port map( B1 => n3352, B2 => n5921, C1 => n3353, C2 => 
                           n5953, A => n3354, ZN => n3344);
   U4175 : OAI22_X1 port map( A1 => n4705, A2 => n3355, B1 => n4673, B2 => 
                           n3356, ZN => n3354);
   U4176 : AOI221_X1 port map( B1 => n1753, B2 => n5985, C1 => n3358, C2 => 
                           n6017, A => n3359, ZN => n3343);
   U4177 : OAI222_X1 port map( A1 => n4801, A2 => n3360, B1 => n4769, B2 => 
                           n3361, C1 => n4737, C2 => n424, ZN => n3359);
   U4178 : AOI221_X1 port map( B1 => n3362, B2 => n6081, C1 => n3363, C2 => 
                           n6049, A => n3364, ZN => n3342);
   U4179 : OAI22_X1 port map( A1 => n5689, A2 => n3365, B1 => n5688, B2 => 
                           n3366, ZN => n3364);
   U4180 : INV_X1 port map( A => DATAIN(31), ZN => n1947);
   U4181 : OAI21_X1 port map( B1 => n3266, B2 => n1545, A => ENABLE, ZN => 
                           n7608);
   U4182 : OAI222_X1 port map( A1 => n2052, A2 => n3263, B1 => n3367, B2 => 
                           n3265, C1 => n3266, C2 => n1482, ZN => n7607);
   U4183 : NOR4_X1 port map( A1 => n3368, A2 => n3369, A3 => n3370, A4 => n3371
                           , ZN => n3367);
   U4184 : NAND4_X1 port map( A1 => n3372, A2 => n3373, A3 => n3374, A4 => 
                           n3375, ZN => n3371);
   U4185 : AOI221_X1 port map( B1 => n1748, B2 => n6432, C1 => n3276, C2 => 
                           n6464, A => n3376, ZN => n3375);
   U4186 : OAI222_X1 port map( A1 => n5280, A2 => n3278, B1 => n5248, B2 => 
                           n3279, C1 => n5216, C2 => n421, ZN => n3376);
   U4187 : AOI221_X1 port map( B1 => n3280, B2 => n716, C1 => n3281, C2 => n292
                           , A => n3377, ZN => n3374);
   U4188 : OAI22_X1 port map( A1 => n196, A2 => n413, B1 => n620, B2 => n3283, 
                           ZN => n3377);
   U4189 : AOI221_X1 port map( B1 => n1754, B2 => n6560, C1 => n3285, C2 => 
                           n6592, A => n3378, ZN => n3373);
   U4190 : OAI222_X1 port map( A1 => n5376, A2 => n3287, B1 => n5344, B2 => 
                           n1579, C1 => n5312, C2 => n3288, ZN => n3378);
   U4191 : AOI221_X1 port map( B1 => n3289, B2 => n717, C1 => n3290, C2 => n293
                           , A => n3379, ZN => n3372);
   U4192 : OAI22_X1 port map( A1 => n197, A2 => n414, B1 => n621, B2 => n3292, 
                           ZN => n3379);
   U4193 : NAND4_X1 port map( A1 => n3380, A2 => n3381, A3 => n3382, A4 => 
                           n3383, ZN => n3370);
   U4194 : AOI221_X1 port map( B1 => n3297, B2 => n6304, C1 => n3298, C2 => 
                           n6336, A => n3384, ZN => n3383);
   U4195 : OAI222_X1 port map( A1 => n5088, A2 => n3300, B1 => n5056, B2 => 
                           n3301, C1 => n5024, C2 => n3302, ZN => n3384);
   U4196 : AOI221_X1 port map( B1 => n3303, B2 => n522, C1 => n3304, C2 => n162
                           , A => n3385, ZN => n3382);
   U4197 : OAI22_X1 port map( A1 => n426, A2 => n3306, B1 => n66, B2 => n3307, 
                           ZN => n3385);
   U4198 : AOI221_X1 port map( B1 => n3308, B2 => n6368, C1 => n3309, C2 => 
                           n6400, A => n3386, ZN => n3381);
   U4199 : OAI222_X1 port map( A1 => n5184, A2 => n3311, B1 => n5152, B2 => 
                           n3312, C1 => n5120, C2 => n422, ZN => n3386);
   U4200 : AOI221_X1 port map( B1 => n3313, B2 => n555, C1 => n3314, C2 => n99,
                           A => n3387, ZN => n3380);
   U4201 : OAI22_X1 port map( A1 => n3, A2 => n415, B1 => n459, B2 => n3316, ZN
                           => n3387);
   U4202 : NAND4_X1 port map( A1 => n3388, A2 => n3389, A3 => n3390, A4 => 
                           n3391, ZN => n3369);
   U4203 : AOI221_X1 port map( B1 => n3321, B2 => n6112, C1 => n3322, C2 => 
                           n6144, A => n3392, ZN => n3391);
   U4204 : OAI222_X1 port map( A1 => n4896, A2 => n3324, B1 => n4864, B2 => 
                           n3325, C1 => n4832, C2 => n423, ZN => n3392);
   U4205 : AOI221_X1 port map( B1 => n3326, B2 => n718, C1 => n3327, C2 => n294
                           , A => n3393, ZN => n3390);
   U4206 : OAI22_X1 port map( A1 => n198, A2 => n3329, B1 => n622, B2 => n3330,
                           ZN => n3393);
   U4207 : AOI221_X1 port map( B1 => n3331, B2 => n6240, C1 => n3332, C2 => 
                           n6272, A => n3394, ZN => n3389);
   U4208 : OAI222_X1 port map( A1 => n4992, A2 => n3334, B1 => n4960, B2 => 
                           n3335, C1 => n4928, C2 => n3336, ZN => n3394);
   U4209 : AOI221_X1 port map( B1 => n3337, B2 => n556, C1 => n3338, C2 => n100
                           , A => n3395, ZN => n3388);
   U4210 : OAI22_X1 port map( A1 => n4, A2 => n3340, B1 => n460, B2 => n3341, 
                           ZN => n3395);
   U4211 : NAND4_X1 port map( A1 => n3396, A2 => n3397, A3 => n3398, A4 => 
                           n3399, ZN => n3368);
   U4212 : AOI221_X1 port map( B1 => n3346, B2 => n5856, C1 => n3347, C2 => 
                           n5888, A => n3400, ZN => n3399);
   U4213 : OAI222_X1 port map( A1 => n4640, A2 => n3349, B1 => n4608, B2 => 
                           n3350, C1 => n4576, C2 => n3351, ZN => n3400);
   U4214 : AOI221_X1 port map( B1 => n3352, B2 => n5920, C1 => n3353, C2 => 
                           n5952, A => n3401, ZN => n3398);
   U4215 : OAI22_X1 port map( A1 => n4704, A2 => n3355, B1 => n4672, B2 => 
                           n3356, ZN => n3401);
   U4216 : AOI221_X1 port map( B1 => n1753, B2 => n5984, C1 => n3358, C2 => 
                           n6016, A => n3402, ZN => n3397);
   U4217 : OAI222_X1 port map( A1 => n4800, A2 => n3360, B1 => n4768, B2 => 
                           n3361, C1 => n4736, C2 => n424, ZN => n3402);
   U4218 : AOI221_X1 port map( B1 => n3362, B2 => n6080, C1 => n3363, C2 => 
                           n6048, A => n3403, ZN => n3396);
   U4219 : OAI22_X1 port map( A1 => n5679, A2 => n3365, B1 => n5678, B2 => 
                           n3366, ZN => n3403);
   U4220 : INV_X1 port map( A => DATAIN(30), ZN => n2052);
   U4221 : OAI21_X1 port map( B1 => n3266, B2 => n1546, A => ENABLE, ZN => 
                           n7606);
   U4222 : OAI222_X1 port map( A1 => n2090, A2 => n3263, B1 => n3404, B2 => 
                           n3265, C1 => n3266, C2 => n1483, ZN => n7605);
   U4223 : NOR4_X1 port map( A1 => n3405, A2 => n3406, A3 => n3407, A4 => n3408
                           , ZN => n3404);
   U4224 : NAND4_X1 port map( A1 => n3409, A2 => n3410, A3 => n3411, A4 => 
                           n3412, ZN => n3408);
   U4225 : AOI221_X1 port map( B1 => n1748, B2 => n6431, C1 => n3276, C2 => 
                           n6463, A => n3413, ZN => n3412);
   U4226 : OAI222_X1 port map( A1 => n5279, A2 => n3278, B1 => n5247, B2 => 
                           n3279, C1 => n5215, C2 => n421, ZN => n3413);
   U4227 : AOI221_X1 port map( B1 => n3280, B2 => n719, C1 => n3281, C2 => n295
                           , A => n3414, ZN => n3411);
   U4228 : OAI22_X1 port map( A1 => n199, A2 => n413, B1 => n623, B2 => n3283, 
                           ZN => n3414);
   U4229 : AOI221_X1 port map( B1 => n1754, B2 => n6559, C1 => n3285, C2 => 
                           n6591, A => n3415, ZN => n3410);
   U4230 : OAI222_X1 port map( A1 => n5375, A2 => n3287, B1 => n5343, B2 => 
                           n1579, C1 => n5311, C2 => n3288, ZN => n3415);
   U4231 : AOI221_X1 port map( B1 => n3289, B2 => n720, C1 => n3290, C2 => n296
                           , A => n3416, ZN => n3409);
   U4232 : OAI22_X1 port map( A1 => n200, A2 => n414, B1 => n624, B2 => n3292, 
                           ZN => n3416);
   U4233 : NAND4_X1 port map( A1 => n3417, A2 => n3418, A3 => n3419, A4 => 
                           n3420, ZN => n3407);
   U4234 : AOI221_X1 port map( B1 => n3297, B2 => n6303, C1 => n3298, C2 => 
                           n6335, A => n3421, ZN => n3420);
   U4235 : OAI222_X1 port map( A1 => n5087, A2 => n3300, B1 => n5055, B2 => 
                           n3301, C1 => n5023, C2 => n3302, ZN => n3421);
   U4236 : AOI221_X1 port map( B1 => n3303, B2 => n523, C1 => n3304, C2 => n163
                           , A => n3422, ZN => n3419);
   U4237 : OAI22_X1 port map( A1 => n427, A2 => n3306, B1 => n67, B2 => n3307, 
                           ZN => n3422);
   U4238 : AOI221_X1 port map( B1 => n3308, B2 => n6367, C1 => n3309, C2 => 
                           n6399, A => n3423, ZN => n3418);
   U4239 : OAI222_X1 port map( A1 => n5183, A2 => n3311, B1 => n5151, B2 => 
                           n3312, C1 => n5119, C2 => n422, ZN => n3423);
   U4240 : AOI221_X1 port map( B1 => n3313, B2 => n557, C1 => n3314, C2 => n101
                           , A => n3424, ZN => n3417);
   U4241 : OAI22_X1 port map( A1 => n5, A2 => n415, B1 => n461, B2 => n3316, ZN
                           => n3424);
   U4242 : NAND4_X1 port map( A1 => n3425, A2 => n3426, A3 => n3427, A4 => 
                           n3428, ZN => n3406);
   U4243 : AOI221_X1 port map( B1 => n3321, B2 => n6111, C1 => n3322, C2 => 
                           n6143, A => n3429, ZN => n3428);
   U4244 : OAI222_X1 port map( A1 => n4895, A2 => n3324, B1 => n4863, B2 => 
                           n3325, C1 => n4831, C2 => n423, ZN => n3429);
   U4245 : AOI221_X1 port map( B1 => n3326, B2 => n721, C1 => n3327, C2 => n297
                           , A => n3430, ZN => n3427);
   U4246 : OAI22_X1 port map( A1 => n201, A2 => n3329, B1 => n625, B2 => n3330,
                           ZN => n3430);
   U4247 : AOI221_X1 port map( B1 => n3331, B2 => n6239, C1 => n3332, C2 => 
                           n6271, A => n3431, ZN => n3426);
   U4248 : OAI222_X1 port map( A1 => n4991, A2 => n3334, B1 => n4959, B2 => 
                           n3335, C1 => n4927, C2 => n3336, ZN => n3431);
   U4249 : AOI221_X1 port map( B1 => n3337, B2 => n558, C1 => n3338, C2 => n102
                           , A => n3432, ZN => n3425);
   U4250 : OAI22_X1 port map( A1 => n6, A2 => n3340, B1 => n462, B2 => n3341, 
                           ZN => n3432);
   U4251 : NAND4_X1 port map( A1 => n3433, A2 => n3434, A3 => n3435, A4 => 
                           n3436, ZN => n3405);
   U4252 : AOI221_X1 port map( B1 => n3346, B2 => n5855, C1 => n3347, C2 => 
                           n5887, A => n3437, ZN => n3436);
   U4253 : OAI222_X1 port map( A1 => n4639, A2 => n3349, B1 => n4607, B2 => 
                           n3350, C1 => n4575, C2 => n3351, ZN => n3437);
   U4254 : AOI221_X1 port map( B1 => n3352, B2 => n5919, C1 => n3353, C2 => 
                           n5951, A => n3438, ZN => n3435);
   U4255 : OAI22_X1 port map( A1 => n4703, A2 => n3355, B1 => n4671, B2 => 
                           n3356, ZN => n3438);
   U4256 : AOI221_X1 port map( B1 => n1753, B2 => n5983, C1 => n3358, C2 => 
                           n6015, A => n3439, ZN => n3434);
   U4257 : OAI222_X1 port map( A1 => n4799, A2 => n3360, B1 => n4767, B2 => 
                           n3361, C1 => n4735, C2 => n424, ZN => n3439);
   U4258 : AOI221_X1 port map( B1 => n3362, B2 => n6079, C1 => n3363, C2 => 
                           n6047, A => n3440, ZN => n3433);
   U4259 : OAI22_X1 port map( A1 => n5669, A2 => n3365, B1 => n5668, B2 => 
                           n3366, ZN => n3440);
   U4260 : INV_X1 port map( A => DATAIN(29), ZN => n2090);
   U4261 : OAI21_X1 port map( B1 => n3266, B2 => n1547, A => ENABLE, ZN => 
                           n7604);
   U4262 : OAI222_X1 port map( A1 => n2128, A2 => n3263, B1 => n3441, B2 => 
                           n3265, C1 => n3266, C2 => n1484, ZN => n7603);
   U4263 : NOR4_X1 port map( A1 => n3442, A2 => n3443, A3 => n3444, A4 => n3445
                           , ZN => n3441);
   U4264 : NAND4_X1 port map( A1 => n3446, A2 => n3447, A3 => n3448, A4 => 
                           n3449, ZN => n3445);
   U4265 : AOI221_X1 port map( B1 => n1748, B2 => n6430, C1 => n3276, C2 => 
                           n6462, A => n3450, ZN => n3449);
   U4266 : OAI222_X1 port map( A1 => n5278, A2 => n3278, B1 => n5246, B2 => 
                           n3279, C1 => n5214, C2 => n421, ZN => n3450);
   U4267 : AOI221_X1 port map( B1 => n3280, B2 => n722, C1 => n3281, C2 => n298
                           , A => n3451, ZN => n3448);
   U4268 : OAI22_X1 port map( A1 => n202, A2 => n413, B1 => n626, B2 => n3283, 
                           ZN => n3451);
   U4269 : AOI221_X1 port map( B1 => n1754, B2 => n6558, C1 => n3285, C2 => 
                           n6590, A => n3452, ZN => n3447);
   U4270 : OAI222_X1 port map( A1 => n5374, A2 => n3287, B1 => n5342, B2 => 
                           n1579, C1 => n5310, C2 => n3288, ZN => n3452);
   U4271 : AOI221_X1 port map( B1 => n3289, B2 => n723, C1 => n3290, C2 => n299
                           , A => n3453, ZN => n3446);
   U4272 : OAI22_X1 port map( A1 => n203, A2 => n414, B1 => n627, B2 => n3292, 
                           ZN => n3453);
   U4273 : NAND4_X1 port map( A1 => n3454, A2 => n3455, A3 => n3456, A4 => 
                           n3457, ZN => n3444);
   U4274 : AOI221_X1 port map( B1 => n3297, B2 => n6302, C1 => n3298, C2 => 
                           n6334, A => n3458, ZN => n3457);
   U4275 : OAI222_X1 port map( A1 => n5086, A2 => n3300, B1 => n5054, B2 => 
                           n3301, C1 => n5022, C2 => n3302, ZN => n3458);
   U4276 : AOI221_X1 port map( B1 => n3303, B2 => n524, C1 => n3304, C2 => n164
                           , A => n3459, ZN => n3456);
   U4277 : OAI22_X1 port map( A1 => n428, A2 => n3306, B1 => n68, B2 => n3307, 
                           ZN => n3459);
   U4278 : AOI221_X1 port map( B1 => n3308, B2 => n6366, C1 => n3309, C2 => 
                           n6398, A => n3460, ZN => n3455);
   U4279 : OAI222_X1 port map( A1 => n5182, A2 => n3311, B1 => n5150, B2 => 
                           n3312, C1 => n5118, C2 => n422, ZN => n3460);
   U4280 : AOI221_X1 port map( B1 => n3313, B2 => n559, C1 => n3314, C2 => n103
                           , A => n3461, ZN => n3454);
   U4281 : OAI22_X1 port map( A1 => n7, A2 => n415, B1 => n463, B2 => n3316, ZN
                           => n3461);
   U4282 : NAND4_X1 port map( A1 => n3462, A2 => n3463, A3 => n3464, A4 => 
                           n3465, ZN => n3443);
   U4283 : AOI221_X1 port map( B1 => n3321, B2 => n6110, C1 => n3322, C2 => 
                           n6142, A => n3466, ZN => n3465);
   U4284 : OAI222_X1 port map( A1 => n4894, A2 => n3324, B1 => n4862, B2 => 
                           n3325, C1 => n4830, C2 => n423, ZN => n3466);
   U4285 : AOI221_X1 port map( B1 => n3326, B2 => n724, C1 => n3327, C2 => n300
                           , A => n3467, ZN => n3464);
   U4286 : OAI22_X1 port map( A1 => n204, A2 => n3329, B1 => n628, B2 => n3330,
                           ZN => n3467);
   U4287 : AOI221_X1 port map( B1 => n3331, B2 => n6238, C1 => n3332, C2 => 
                           n6270, A => n3468, ZN => n3463);
   U4288 : OAI222_X1 port map( A1 => n4990, A2 => n3334, B1 => n4958, B2 => 
                           n3335, C1 => n4926, C2 => n3336, ZN => n3468);
   U4289 : AOI221_X1 port map( B1 => n3337, B2 => n560, C1 => n3338, C2 => n104
                           , A => n3469, ZN => n3462);
   U4290 : OAI22_X1 port map( A1 => n8, A2 => n3340, B1 => n464, B2 => n3341, 
                           ZN => n3469);
   U4291 : NAND4_X1 port map( A1 => n3470, A2 => n3471, A3 => n3472, A4 => 
                           n3473, ZN => n3442);
   U4292 : AOI221_X1 port map( B1 => n3346, B2 => n5854, C1 => n3347, C2 => 
                           n5886, A => n3474, ZN => n3473);
   U4293 : OAI222_X1 port map( A1 => n4638, A2 => n3349, B1 => n4606, B2 => 
                           n3350, C1 => n4574, C2 => n3351, ZN => n3474);
   U4294 : AOI221_X1 port map( B1 => n3352, B2 => n5918, C1 => n3353, C2 => 
                           n5950, A => n3475, ZN => n3472);
   U4295 : OAI22_X1 port map( A1 => n4702, A2 => n3355, B1 => n4670, B2 => 
                           n3356, ZN => n3475);
   U4296 : AOI221_X1 port map( B1 => n1753, B2 => n5982, C1 => n3358, C2 => 
                           n6014, A => n3476, ZN => n3471);
   U4297 : OAI222_X1 port map( A1 => n4798, A2 => n3360, B1 => n4766, B2 => 
                           n3361, C1 => n4734, C2 => n424, ZN => n3476);
   U4298 : AOI221_X1 port map( B1 => n3362, B2 => n6078, C1 => n3363, C2 => 
                           n6046, A => n3477, ZN => n3470);
   U4299 : OAI22_X1 port map( A1 => n5659, A2 => n3365, B1 => n5658, B2 => 
                           n3366, ZN => n3477);
   U4300 : INV_X1 port map( A => DATAIN(28), ZN => n2128);
   U4301 : OAI21_X1 port map( B1 => n3266, B2 => n1548, A => ENABLE, ZN => 
                           n7602);
   U4302 : OAI222_X1 port map( A1 => n2166, A2 => n3263, B1 => n3478, B2 => 
                           n3265, C1 => n3266, C2 => n1485, ZN => n7601);
   U4303 : NOR4_X1 port map( A1 => n3479, A2 => n3480, A3 => n3481, A4 => n3482
                           , ZN => n3478);
   U4304 : NAND4_X1 port map( A1 => n3483, A2 => n3484, A3 => n3485, A4 => 
                           n3486, ZN => n3482);
   U4305 : AOI221_X1 port map( B1 => n1748, B2 => n6429, C1 => n3276, C2 => 
                           n6461, A => n3487, ZN => n3486);
   U4306 : OAI222_X1 port map( A1 => n5277, A2 => n3278, B1 => n5245, B2 => 
                           n3279, C1 => n5213, C2 => n421, ZN => n3487);
   U4307 : AOI221_X1 port map( B1 => n3280, B2 => n725, C1 => n3281, C2 => n301
                           , A => n3488, ZN => n3485);
   U4308 : OAI22_X1 port map( A1 => n205, A2 => n413, B1 => n629, B2 => n3283, 
                           ZN => n3488);
   U4309 : AOI221_X1 port map( B1 => n1754, B2 => n6557, C1 => n3285, C2 => 
                           n6589, A => n3489, ZN => n3484);
   U4310 : OAI222_X1 port map( A1 => n5373, A2 => n3287, B1 => n5341, B2 => 
                           n1579, C1 => n5309, C2 => n3288, ZN => n3489);
   U4311 : AOI221_X1 port map( B1 => n3289, B2 => n726, C1 => n3290, C2 => n302
                           , A => n3490, ZN => n3483);
   U4312 : OAI22_X1 port map( A1 => n206, A2 => n414, B1 => n630, B2 => n3292, 
                           ZN => n3490);
   U4313 : NAND4_X1 port map( A1 => n3491, A2 => n3492, A3 => n3493, A4 => 
                           n3494, ZN => n3481);
   U4314 : AOI221_X1 port map( B1 => n3297, B2 => n6301, C1 => n3298, C2 => 
                           n6333, A => n3495, ZN => n3494);
   U4315 : OAI222_X1 port map( A1 => n5085, A2 => n3300, B1 => n5053, B2 => 
                           n3301, C1 => n5021, C2 => n3302, ZN => n3495);
   U4316 : AOI221_X1 port map( B1 => n3303, B2 => n525, C1 => n3304, C2 => n165
                           , A => n3496, ZN => n3493);
   U4317 : OAI22_X1 port map( A1 => n429, A2 => n3306, B1 => n69, B2 => n3307, 
                           ZN => n3496);
   U4318 : AOI221_X1 port map( B1 => n3308, B2 => n6365, C1 => n3309, C2 => 
                           n6397, A => n3497, ZN => n3492);
   U4319 : OAI222_X1 port map( A1 => n5181, A2 => n3311, B1 => n5149, B2 => 
                           n3312, C1 => n5117, C2 => n422, ZN => n3497);
   U4320 : AOI221_X1 port map( B1 => n3313, B2 => n561, C1 => n3314, C2 => n105
                           , A => n3498, ZN => n3491);
   U4321 : OAI22_X1 port map( A1 => n9, A2 => n415, B1 => n465, B2 => n3316, ZN
                           => n3498);
   U4322 : NAND4_X1 port map( A1 => n3499, A2 => n3500, A3 => n3501, A4 => 
                           n3502, ZN => n3480);
   U4323 : AOI221_X1 port map( B1 => n3321, B2 => n6109, C1 => n3322, C2 => 
                           n6141, A => n3503, ZN => n3502);
   U4324 : OAI222_X1 port map( A1 => n4893, A2 => n3324, B1 => n4861, B2 => 
                           n3325, C1 => n4829, C2 => n423, ZN => n3503);
   U4325 : AOI221_X1 port map( B1 => n3326, B2 => n727, C1 => n3327, C2 => n303
                           , A => n3504, ZN => n3501);
   U4326 : OAI22_X1 port map( A1 => n207, A2 => n3329, B1 => n631, B2 => n3330,
                           ZN => n3504);
   U4327 : AOI221_X1 port map( B1 => n3331, B2 => n6237, C1 => n3332, C2 => 
                           n6269, A => n3505, ZN => n3500);
   U4328 : OAI222_X1 port map( A1 => n4989, A2 => n3334, B1 => n4957, B2 => 
                           n3335, C1 => n4925, C2 => n3336, ZN => n3505);
   U4329 : AOI221_X1 port map( B1 => n3337, B2 => n562, C1 => n3338, C2 => n106
                           , A => n3506, ZN => n3499);
   U4330 : OAI22_X1 port map( A1 => n10, A2 => n3340, B1 => n466, B2 => n3341, 
                           ZN => n3506);
   U4331 : NAND4_X1 port map( A1 => n3507, A2 => n3508, A3 => n3509, A4 => 
                           n3510, ZN => n3479);
   U4332 : AOI221_X1 port map( B1 => n3346, B2 => n5853, C1 => n3347, C2 => 
                           n5885, A => n3511, ZN => n3510);
   U4333 : OAI222_X1 port map( A1 => n4637, A2 => n3349, B1 => n4605, B2 => 
                           n3350, C1 => n4573, C2 => n3351, ZN => n3511);
   U4334 : AOI221_X1 port map( B1 => n3352, B2 => n5917, C1 => n3353, C2 => 
                           n5949, A => n3512, ZN => n3509);
   U4335 : OAI22_X1 port map( A1 => n4701, A2 => n3355, B1 => n4669, B2 => 
                           n3356, ZN => n3512);
   U4336 : AOI221_X1 port map( B1 => n1753, B2 => n5981, C1 => n3358, C2 => 
                           n6013, A => n3513, ZN => n3508);
   U4337 : OAI222_X1 port map( A1 => n4797, A2 => n3360, B1 => n4765, B2 => 
                           n3361, C1 => n4733, C2 => n424, ZN => n3513);
   U4338 : AOI221_X1 port map( B1 => n3362, B2 => n6077, C1 => n3363, C2 => 
                           n6045, A => n3514, ZN => n3507);
   U4339 : OAI22_X1 port map( A1 => n5649, A2 => n3365, B1 => n5648, B2 => 
                           n3366, ZN => n3514);
   U4340 : INV_X1 port map( A => DATAIN(27), ZN => n2166);
   U4341 : OAI21_X1 port map( B1 => n3266, B2 => n1549, A => ENABLE, ZN => 
                           n7600);
   U4342 : OAI222_X1 port map( A1 => n2204, A2 => n3263, B1 => n3515, B2 => 
                           n3265, C1 => n3266, C2 => n1486, ZN => n7599);
   U4343 : NOR4_X1 port map( A1 => n3516, A2 => n3517, A3 => n3518, A4 => n3519
                           , ZN => n3515);
   U4344 : NAND4_X1 port map( A1 => n3520, A2 => n3521, A3 => n3522, A4 => 
                           n3523, ZN => n3519);
   U4345 : AOI221_X1 port map( B1 => n1748, B2 => n6428, C1 => n3276, C2 => 
                           n6460, A => n3524, ZN => n3523);
   U4346 : OAI222_X1 port map( A1 => n5276, A2 => n3278, B1 => n5244, B2 => 
                           n3279, C1 => n5212, C2 => n421, ZN => n3524);
   U4347 : AOI221_X1 port map( B1 => n3280, B2 => n728, C1 => n3281, C2 => n304
                           , A => n3525, ZN => n3522);
   U4348 : OAI22_X1 port map( A1 => n208, A2 => n413, B1 => n632, B2 => n3283, 
                           ZN => n3525);
   U4349 : AOI221_X1 port map( B1 => n1754, B2 => n6556, C1 => n3285, C2 => 
                           n6588, A => n3526, ZN => n3521);
   U4350 : OAI222_X1 port map( A1 => n5372, A2 => n3287, B1 => n5340, B2 => 
                           n1579, C1 => n5308, C2 => n3288, ZN => n3526);
   U4351 : AOI221_X1 port map( B1 => n3289, B2 => n729, C1 => n3290, C2 => n305
                           , A => n3527, ZN => n3520);
   U4352 : OAI22_X1 port map( A1 => n209, A2 => n414, B1 => n633, B2 => n3292, 
                           ZN => n3527);
   U4353 : NAND4_X1 port map( A1 => n3528, A2 => n3529, A3 => n3530, A4 => 
                           n3531, ZN => n3518);
   U4354 : AOI221_X1 port map( B1 => n3297, B2 => n6300, C1 => n3298, C2 => 
                           n6332, A => n3532, ZN => n3531);
   U4355 : OAI222_X1 port map( A1 => n5084, A2 => n3300, B1 => n5052, B2 => 
                           n3301, C1 => n5020, C2 => n3302, ZN => n3532);
   U4356 : AOI221_X1 port map( B1 => n3303, B2 => n526, C1 => n3304, C2 => n166
                           , A => n3533, ZN => n3530);
   U4357 : OAI22_X1 port map( A1 => n430, A2 => n3306, B1 => n70, B2 => n3307, 
                           ZN => n3533);
   U4358 : AOI221_X1 port map( B1 => n3308, B2 => n6364, C1 => n3309, C2 => 
                           n6396, A => n3534, ZN => n3529);
   U4359 : OAI222_X1 port map( A1 => n5180, A2 => n3311, B1 => n5148, B2 => 
                           n3312, C1 => n5116, C2 => n422, ZN => n3534);
   U4360 : AOI221_X1 port map( B1 => n3313, B2 => n563, C1 => n3314, C2 => n107
                           , A => n3535, ZN => n3528);
   U4361 : OAI22_X1 port map( A1 => n11, A2 => n415, B1 => n467, B2 => n3316, 
                           ZN => n3535);
   U4362 : NAND4_X1 port map( A1 => n3536, A2 => n3537, A3 => n3538, A4 => 
                           n3539, ZN => n3517);
   U4363 : AOI221_X1 port map( B1 => n3321, B2 => n6108, C1 => n3322, C2 => 
                           n6140, A => n3540, ZN => n3539);
   U4364 : OAI222_X1 port map( A1 => n4892, A2 => n3324, B1 => n4860, B2 => 
                           n3325, C1 => n4828, C2 => n423, ZN => n3540);
   U4365 : AOI221_X1 port map( B1 => n3326, B2 => n730, C1 => n3327, C2 => n306
                           , A => n3541, ZN => n3538);
   U4366 : OAI22_X1 port map( A1 => n210, A2 => n3329, B1 => n634, B2 => n3330,
                           ZN => n3541);
   U4367 : AOI221_X1 port map( B1 => n3331, B2 => n6236, C1 => n3332, C2 => 
                           n6268, A => n3542, ZN => n3537);
   U4368 : OAI222_X1 port map( A1 => n4988, A2 => n3334, B1 => n4956, B2 => 
                           n3335, C1 => n4924, C2 => n3336, ZN => n3542);
   U4369 : AOI221_X1 port map( B1 => n3337, B2 => n564, C1 => n3338, C2 => n108
                           , A => n3543, ZN => n3536);
   U4370 : OAI22_X1 port map( A1 => n12, A2 => n3340, B1 => n468, B2 => n3341, 
                           ZN => n3543);
   U4371 : NAND4_X1 port map( A1 => n3544, A2 => n3545, A3 => n3546, A4 => 
                           n3547, ZN => n3516);
   U4372 : AOI221_X1 port map( B1 => n3346, B2 => n5852, C1 => n3347, C2 => 
                           n5884, A => n3548, ZN => n3547);
   U4373 : OAI222_X1 port map( A1 => n4636, A2 => n3349, B1 => n4604, B2 => 
                           n3350, C1 => n4572, C2 => n3351, ZN => n3548);
   U4374 : AOI221_X1 port map( B1 => n3352, B2 => n5916, C1 => n3353, C2 => 
                           n5948, A => n3549, ZN => n3546);
   U4375 : OAI22_X1 port map( A1 => n4700, A2 => n3355, B1 => n4668, B2 => 
                           n3356, ZN => n3549);
   U4376 : AOI221_X1 port map( B1 => n1753, B2 => n5980, C1 => n3358, C2 => 
                           n6012, A => n3550, ZN => n3545);
   U4377 : OAI222_X1 port map( A1 => n4796, A2 => n3360, B1 => n4764, B2 => 
                           n3361, C1 => n4732, C2 => n424, ZN => n3550);
   U4378 : AOI221_X1 port map( B1 => n3362, B2 => n6076, C1 => n3363, C2 => 
                           n6044, A => n3551, ZN => n3544);
   U4379 : OAI22_X1 port map( A1 => n5639, A2 => n3365, B1 => n5638, B2 => 
                           n3366, ZN => n3551);
   U4380 : INV_X1 port map( A => DATAIN(26), ZN => n2204);
   U4381 : OAI21_X1 port map( B1 => n3266, B2 => n1550, A => ENABLE, ZN => 
                           n7598);
   U4382 : OAI222_X1 port map( A1 => n2242, A2 => n3263, B1 => n3552, B2 => 
                           n3265, C1 => n3266, C2 => n1487, ZN => n7597);
   U4383 : NOR4_X1 port map( A1 => n3553, A2 => n3554, A3 => n3555, A4 => n3556
                           , ZN => n3552);
   U4384 : NAND4_X1 port map( A1 => n3557, A2 => n3558, A3 => n3559, A4 => 
                           n3560, ZN => n3556);
   U4385 : AOI221_X1 port map( B1 => n1748, B2 => n6427, C1 => n3276, C2 => 
                           n6459, A => n3561, ZN => n3560);
   U4386 : OAI222_X1 port map( A1 => n5275, A2 => n3278, B1 => n5243, B2 => 
                           n3279, C1 => n5211, C2 => n421, ZN => n3561);
   U4387 : AOI221_X1 port map( B1 => n3280, B2 => n731, C1 => n3281, C2 => n307
                           , A => n3562, ZN => n3559);
   U4388 : OAI22_X1 port map( A1 => n211, A2 => n413, B1 => n635, B2 => n3283, 
                           ZN => n3562);
   U4389 : AOI221_X1 port map( B1 => n1754, B2 => n6555, C1 => n3285, C2 => 
                           n6587, A => n3563, ZN => n3558);
   U4390 : OAI222_X1 port map( A1 => n5371, A2 => n3287, B1 => n5339, B2 => 
                           n1579, C1 => n5307, C2 => n3288, ZN => n3563);
   U4391 : AOI221_X1 port map( B1 => n3289, B2 => n732, C1 => n3290, C2 => n308
                           , A => n3564, ZN => n3557);
   U4392 : OAI22_X1 port map( A1 => n212, A2 => n414, B1 => n636, B2 => n3292, 
                           ZN => n3564);
   U4393 : NAND4_X1 port map( A1 => n3565, A2 => n3566, A3 => n3567, A4 => 
                           n3568, ZN => n3555);
   U4394 : AOI221_X1 port map( B1 => n3297, B2 => n6299, C1 => n3298, C2 => 
                           n6331, A => n3569, ZN => n3568);
   U4395 : OAI222_X1 port map( A1 => n5083, A2 => n3300, B1 => n5051, B2 => 
                           n3301, C1 => n5019, C2 => n3302, ZN => n3569);
   U4396 : AOI221_X1 port map( B1 => n3303, B2 => n527, C1 => n3304, C2 => n167
                           , A => n3570, ZN => n3567);
   U4397 : OAI22_X1 port map( A1 => n431, A2 => n3306, B1 => n71, B2 => n3307, 
                           ZN => n3570);
   U4398 : AOI221_X1 port map( B1 => n3308, B2 => n6363, C1 => n3309, C2 => 
                           n6395, A => n3571, ZN => n3566);
   U4399 : OAI222_X1 port map( A1 => n5179, A2 => n3311, B1 => n5147, B2 => 
                           n3312, C1 => n5115, C2 => n422, ZN => n3571);
   U4400 : AOI221_X1 port map( B1 => n3313, B2 => n565, C1 => n3314, C2 => n109
                           , A => n3572, ZN => n3565);
   U4401 : OAI22_X1 port map( A1 => n13, A2 => n415, B1 => n469, B2 => n3316, 
                           ZN => n3572);
   U4402 : NAND4_X1 port map( A1 => n3573, A2 => n3574, A3 => n3575, A4 => 
                           n3576, ZN => n3554);
   U4403 : AOI221_X1 port map( B1 => n3321, B2 => n6107, C1 => n3322, C2 => 
                           n6139, A => n3577, ZN => n3576);
   U4404 : OAI222_X1 port map( A1 => n4891, A2 => n3324, B1 => n4859, B2 => 
                           n3325, C1 => n4827, C2 => n423, ZN => n3577);
   U4405 : AOI221_X1 port map( B1 => n3326, B2 => n733, C1 => n3327, C2 => n309
                           , A => n3578, ZN => n3575);
   U4406 : OAI22_X1 port map( A1 => n213, A2 => n3329, B1 => n637, B2 => n3330,
                           ZN => n3578);
   U4407 : AOI221_X1 port map( B1 => n3331, B2 => n6235, C1 => n3332, C2 => 
                           n6267, A => n3579, ZN => n3574);
   U4408 : OAI222_X1 port map( A1 => n4987, A2 => n3334, B1 => n4955, B2 => 
                           n3335, C1 => n4923, C2 => n3336, ZN => n3579);
   U4409 : AOI221_X1 port map( B1 => n3337, B2 => n566, C1 => n3338, C2 => n110
                           , A => n3580, ZN => n3573);
   U4410 : OAI22_X1 port map( A1 => n14, A2 => n3340, B1 => n470, B2 => n3341, 
                           ZN => n3580);
   U4411 : NAND4_X1 port map( A1 => n3581, A2 => n3582, A3 => n3583, A4 => 
                           n3584, ZN => n3553);
   U4412 : AOI221_X1 port map( B1 => n3346, B2 => n5851, C1 => n3347, C2 => 
                           n5883, A => n3585, ZN => n3584);
   U4413 : OAI222_X1 port map( A1 => n4635, A2 => n3349, B1 => n4603, B2 => 
                           n3350, C1 => n4571, C2 => n3351, ZN => n3585);
   U4414 : AOI221_X1 port map( B1 => n3352, B2 => n5915, C1 => n3353, C2 => 
                           n5947, A => n3586, ZN => n3583);
   U4415 : OAI22_X1 port map( A1 => n4699, A2 => n3355, B1 => n4667, B2 => 
                           n3356, ZN => n3586);
   U4416 : AOI221_X1 port map( B1 => n1753, B2 => n5979, C1 => n3358, C2 => 
                           n6011, A => n3587, ZN => n3582);
   U4417 : OAI222_X1 port map( A1 => n4795, A2 => n3360, B1 => n4763, B2 => 
                           n3361, C1 => n4731, C2 => n424, ZN => n3587);
   U4418 : AOI221_X1 port map( B1 => n3362, B2 => n6075, C1 => n3363, C2 => 
                           n6043, A => n3588, ZN => n3581);
   U4419 : OAI22_X1 port map( A1 => n5629, A2 => n3365, B1 => n5628, B2 => 
                           n3366, ZN => n3588);
   U4420 : INV_X1 port map( A => DATAIN(25), ZN => n2242);
   U4421 : OAI21_X1 port map( B1 => n3266, B2 => n1551, A => ENABLE, ZN => 
                           n7596);
   U4422 : OAI222_X1 port map( A1 => n2280, A2 => n3263, B1 => n3589, B2 => 
                           n3265, C1 => n3266, C2 => n1488, ZN => n7595);
   U4423 : NOR4_X1 port map( A1 => n3590, A2 => n3591, A3 => n3592, A4 => n3593
                           , ZN => n3589);
   U4424 : NAND4_X1 port map( A1 => n3594, A2 => n3595, A3 => n3596, A4 => 
                           n3597, ZN => n3593);
   U4425 : AOI221_X1 port map( B1 => n3275, B2 => n6426, C1 => n3276, C2 => 
                           n6458, A => n3598, ZN => n3597);
   U4426 : OAI222_X1 port map( A1 => n5274, A2 => n3278, B1 => n5242, B2 => 
                           n3279, C1 => n5210, C2 => n421, ZN => n3598);
   U4427 : AOI221_X1 port map( B1 => n3280, B2 => n734, C1 => n3281, C2 => n310
                           , A => n3599, ZN => n3596);
   U4428 : OAI22_X1 port map( A1 => n214, A2 => n413, B1 => n638, B2 => n3283, 
                           ZN => n3599);
   U4429 : AOI221_X1 port map( B1 => n3284, B2 => n6554, C1 => n3285, C2 => 
                           n6586, A => n3600, ZN => n3595);
   U4430 : OAI222_X1 port map( A1 => n5370, A2 => n3287, B1 => n5338, B2 => 
                           n1579, C1 => n5306, C2 => n3288, ZN => n3600);
   U4431 : AOI221_X1 port map( B1 => n3289, B2 => n735, C1 => n3290, C2 => n311
                           , A => n3601, ZN => n3594);
   U4432 : OAI22_X1 port map( A1 => n215, A2 => n414, B1 => n639, B2 => n3292, 
                           ZN => n3601);
   U4433 : NAND4_X1 port map( A1 => n3602, A2 => n3603, A3 => n3604, A4 => 
                           n3605, ZN => n3592);
   U4434 : AOI221_X1 port map( B1 => n3297, B2 => n6298, C1 => n3298, C2 => 
                           n6330, A => n3606, ZN => n3605);
   U4435 : OAI222_X1 port map( A1 => n5082, A2 => n3300, B1 => n5050, B2 => 
                           n3301, C1 => n5018, C2 => n3302, ZN => n3606);
   U4436 : AOI221_X1 port map( B1 => n3303, B2 => n528, C1 => n3304, C2 => n168
                           , A => n3607, ZN => n3604);
   U4437 : OAI22_X1 port map( A1 => n432, A2 => n3306, B1 => n72, B2 => n3307, 
                           ZN => n3607);
   U4438 : AOI221_X1 port map( B1 => n3308, B2 => n6362, C1 => n3309, C2 => 
                           n6394, A => n3608, ZN => n3603);
   U4439 : OAI222_X1 port map( A1 => n5178, A2 => n3311, B1 => n5146, B2 => 
                           n3312, C1 => n5114, C2 => n422, ZN => n3608);
   U4440 : AOI221_X1 port map( B1 => n3313, B2 => n567, C1 => n3314, C2 => n111
                           , A => n3609, ZN => n3602);
   U4441 : OAI22_X1 port map( A1 => n15, A2 => n415, B1 => n471, B2 => n3316, 
                           ZN => n3609);
   U4442 : NAND4_X1 port map( A1 => n3610, A2 => n3611, A3 => n3612, A4 => 
                           n3613, ZN => n3591);
   U4443 : AOI221_X1 port map( B1 => n3321, B2 => n6106, C1 => n3322, C2 => 
                           n6138, A => n3614, ZN => n3613);
   U4444 : OAI222_X1 port map( A1 => n4890, A2 => n3324, B1 => n4858, B2 => 
                           n3325, C1 => n4826, C2 => n423, ZN => n3614);
   U4445 : AOI221_X1 port map( B1 => n3326, B2 => n736, C1 => n3327, C2 => n312
                           , A => n3615, ZN => n3612);
   U4446 : OAI22_X1 port map( A1 => n216, A2 => n3329, B1 => n640, B2 => n3330,
                           ZN => n3615);
   U4447 : AOI221_X1 port map( B1 => n3331, B2 => n6234, C1 => n3332, C2 => 
                           n6266, A => n3616, ZN => n3611);
   U4448 : OAI222_X1 port map( A1 => n4986, A2 => n3334, B1 => n4954, B2 => 
                           n3335, C1 => n4922, C2 => n3336, ZN => n3616);
   U4449 : AOI221_X1 port map( B1 => n3337, B2 => n568, C1 => n3338, C2 => n112
                           , A => n3617, ZN => n3610);
   U4450 : OAI22_X1 port map( A1 => n16, A2 => n3340, B1 => n472, B2 => n3341, 
                           ZN => n3617);
   U4451 : NAND4_X1 port map( A1 => n3618, A2 => n3619, A3 => n3620, A4 => 
                           n3621, ZN => n3590);
   U4452 : AOI221_X1 port map( B1 => n3346, B2 => n5850, C1 => n3347, C2 => 
                           n5882, A => n3622, ZN => n3621);
   U4453 : OAI222_X1 port map( A1 => n4634, A2 => n3349, B1 => n4602, B2 => 
                           n3350, C1 => n4570, C2 => n3351, ZN => n3622);
   U4454 : AOI221_X1 port map( B1 => n3352, B2 => n5914, C1 => n3353, C2 => 
                           n5946, A => n3623, ZN => n3620);
   U4455 : OAI22_X1 port map( A1 => n4698, A2 => n3355, B1 => n4666, B2 => 
                           n3356, ZN => n3623);
   U4456 : AOI221_X1 port map( B1 => n3357, B2 => n5978, C1 => n3358, C2 => 
                           n6010, A => n3624, ZN => n3619);
   U4457 : OAI222_X1 port map( A1 => n4794, A2 => n3360, B1 => n4762, B2 => 
                           n3361, C1 => n4730, C2 => n424, ZN => n3624);
   U4458 : AOI221_X1 port map( B1 => n3362, B2 => n6074, C1 => n3363, C2 => 
                           n6042, A => n3625, ZN => n3618);
   U4459 : OAI22_X1 port map( A1 => n5619, A2 => n3365, B1 => n5618, B2 => 
                           n3366, ZN => n3625);
   U4460 : INV_X1 port map( A => DATAIN(24), ZN => n2280);
   U4461 : OAI21_X1 port map( B1 => n3266, B2 => n1552, A => ENABLE, ZN => 
                           n7594);
   U4462 : OAI222_X1 port map( A1 => n2318, A2 => n3263, B1 => n3626, B2 => 
                           n3265, C1 => n3266, C2 => n1489, ZN => n7593);
   U4463 : NOR4_X1 port map( A1 => n3627, A2 => n3628, A3 => n3629, A4 => n3630
                           , ZN => n3626);
   U4464 : NAND4_X1 port map( A1 => n3631, A2 => n3632, A3 => n3633, A4 => 
                           n3634, ZN => n3630);
   U4465 : AOI221_X1 port map( B1 => n3275, B2 => n6425, C1 => n3276, C2 => 
                           n6457, A => n3635, ZN => n3634);
   U4466 : OAI222_X1 port map( A1 => n5273, A2 => n3278, B1 => n5241, B2 => 
                           n3279, C1 => n5209, C2 => n421, ZN => n3635);
   U4467 : AOI221_X1 port map( B1 => n3280, B2 => n737, C1 => n3281, C2 => n313
                           , A => n3636, ZN => n3633);
   U4468 : OAI22_X1 port map( A1 => n217, A2 => n413, B1 => n641, B2 => n3283, 
                           ZN => n3636);
   U4469 : AOI221_X1 port map( B1 => n3284, B2 => n6553, C1 => n3285, C2 => 
                           n6585, A => n3637, ZN => n3632);
   U4470 : OAI222_X1 port map( A1 => n5369, A2 => n3287, B1 => n5337, B2 => 
                           n1579, C1 => n5305, C2 => n3288, ZN => n3637);
   U4471 : AOI221_X1 port map( B1 => n3289, B2 => n738, C1 => n3290, C2 => n314
                           , A => n3638, ZN => n3631);
   U4472 : OAI22_X1 port map( A1 => n218, A2 => n414, B1 => n642, B2 => n3292, 
                           ZN => n3638);
   U4473 : NAND4_X1 port map( A1 => n3639, A2 => n3640, A3 => n3641, A4 => 
                           n3642, ZN => n3629);
   U4474 : AOI221_X1 port map( B1 => n3297, B2 => n6297, C1 => n3298, C2 => 
                           n6329, A => n3643, ZN => n3642);
   U4475 : OAI222_X1 port map( A1 => n5081, A2 => n3300, B1 => n5049, B2 => 
                           n3301, C1 => n5017, C2 => n3302, ZN => n3643);
   U4476 : AOI221_X1 port map( B1 => n3303, B2 => n529, C1 => n3304, C2 => n169
                           , A => n3644, ZN => n3641);
   U4477 : OAI22_X1 port map( A1 => n433, A2 => n3306, B1 => n73, B2 => n3307, 
                           ZN => n3644);
   U4478 : AOI221_X1 port map( B1 => n3308, B2 => n6361, C1 => n3309, C2 => 
                           n6393, A => n3645, ZN => n3640);
   U4479 : OAI222_X1 port map( A1 => n5177, A2 => n3311, B1 => n5145, B2 => 
                           n3312, C1 => n5113, C2 => n422, ZN => n3645);
   U4480 : AOI221_X1 port map( B1 => n3313, B2 => n569, C1 => n3314, C2 => n113
                           , A => n3646, ZN => n3639);
   U4481 : OAI22_X1 port map( A1 => n17, A2 => n415, B1 => n473, B2 => n3316, 
                           ZN => n3646);
   U4482 : NAND4_X1 port map( A1 => n3647, A2 => n3648, A3 => n3649, A4 => 
                           n3650, ZN => n3628);
   U4483 : AOI221_X1 port map( B1 => n3321, B2 => n6105, C1 => n3322, C2 => 
                           n6137, A => n3651, ZN => n3650);
   U4484 : OAI222_X1 port map( A1 => n4889, A2 => n3324, B1 => n4857, B2 => 
                           n3325, C1 => n4825, C2 => n423, ZN => n3651);
   U4485 : AOI221_X1 port map( B1 => n3326, B2 => n739, C1 => n3327, C2 => n315
                           , A => n3652, ZN => n3649);
   U4486 : OAI22_X1 port map( A1 => n219, A2 => n3329, B1 => n643, B2 => n3330,
                           ZN => n3652);
   U4487 : AOI221_X1 port map( B1 => n3331, B2 => n6233, C1 => n3332, C2 => 
                           n6265, A => n3653, ZN => n3648);
   U4488 : OAI222_X1 port map( A1 => n4985, A2 => n3334, B1 => n4953, B2 => 
                           n3335, C1 => n4921, C2 => n3336, ZN => n3653);
   U4489 : AOI221_X1 port map( B1 => n3337, B2 => n570, C1 => n3338, C2 => n114
                           , A => n3654, ZN => n3647);
   U4490 : OAI22_X1 port map( A1 => n18, A2 => n3340, B1 => n474, B2 => n3341, 
                           ZN => n3654);
   U4491 : NAND4_X1 port map( A1 => n3655, A2 => n3656, A3 => n3657, A4 => 
                           n3658, ZN => n3627);
   U4492 : AOI221_X1 port map( B1 => n3346, B2 => n5849, C1 => n3347, C2 => 
                           n5881, A => n3659, ZN => n3658);
   U4493 : OAI222_X1 port map( A1 => n4633, A2 => n3349, B1 => n4601, B2 => 
                           n3350, C1 => n4569, C2 => n3351, ZN => n3659);
   U4494 : AOI221_X1 port map( B1 => n3352, B2 => n5913, C1 => n3353, C2 => 
                           n5945, A => n3660, ZN => n3657);
   U4495 : OAI22_X1 port map( A1 => n4697, A2 => n3355, B1 => n4665, B2 => 
                           n3356, ZN => n3660);
   U4496 : AOI221_X1 port map( B1 => n3357, B2 => n5977, C1 => n3358, C2 => 
                           n6009, A => n3661, ZN => n3656);
   U4497 : OAI222_X1 port map( A1 => n4793, A2 => n3360, B1 => n4761, B2 => 
                           n3361, C1 => n4729, C2 => n424, ZN => n3661);
   U4498 : AOI221_X1 port map( B1 => n3362, B2 => n6073, C1 => n3363, C2 => 
                           n6041, A => n3662, ZN => n3655);
   U4499 : OAI22_X1 port map( A1 => n5609, A2 => n3365, B1 => n5608, B2 => 
                           n3366, ZN => n3662);
   U4500 : INV_X1 port map( A => DATAIN(23), ZN => n2318);
   U4501 : OAI21_X1 port map( B1 => n3266, B2 => n1553, A => ENABLE, ZN => 
                           n7592);
   U4502 : OAI222_X1 port map( A1 => n2356, A2 => n3263, B1 => n3663, B2 => 
                           n3265, C1 => n3266, C2 => n1490, ZN => n7591);
   U4503 : NOR4_X1 port map( A1 => n3664, A2 => n3665, A3 => n3666, A4 => n3667
                           , ZN => n3663);
   U4504 : NAND4_X1 port map( A1 => n3668, A2 => n3669, A3 => n3670, A4 => 
                           n3671, ZN => n3667);
   U4505 : AOI221_X1 port map( B1 => n3275, B2 => n6424, C1 => n3276, C2 => 
                           n6456, A => n3672, ZN => n3671);
   U4506 : OAI222_X1 port map( A1 => n5272, A2 => n3278, B1 => n5240, B2 => 
                           n3279, C1 => n5208, C2 => n421, ZN => n3672);
   U4507 : AOI221_X1 port map( B1 => n3280, B2 => n740, C1 => n3281, C2 => n316
                           , A => n3673, ZN => n3670);
   U4508 : OAI22_X1 port map( A1 => n220, A2 => n413, B1 => n644, B2 => n3283, 
                           ZN => n3673);
   U4509 : AOI221_X1 port map( B1 => n3284, B2 => n6552, C1 => n3285, C2 => 
                           n6584, A => n3674, ZN => n3669);
   U4510 : OAI222_X1 port map( A1 => n5368, A2 => n3287, B1 => n5336, B2 => 
                           n1579, C1 => n5304, C2 => n3288, ZN => n3674);
   U4511 : AOI221_X1 port map( B1 => n3289, B2 => n741, C1 => n3290, C2 => n317
                           , A => n3675, ZN => n3668);
   U4512 : OAI22_X1 port map( A1 => n221, A2 => n414, B1 => n645, B2 => n3292, 
                           ZN => n3675);
   U4513 : NAND4_X1 port map( A1 => n3676, A2 => n3677, A3 => n3678, A4 => 
                           n3679, ZN => n3666);
   U4514 : AOI221_X1 port map( B1 => n3297, B2 => n6296, C1 => n3298, C2 => 
                           n6328, A => n3680, ZN => n3679);
   U4515 : OAI222_X1 port map( A1 => n5080, A2 => n3300, B1 => n5048, B2 => 
                           n3301, C1 => n5016, C2 => n3302, ZN => n3680);
   U4516 : AOI221_X1 port map( B1 => n3303, B2 => n530, C1 => n3304, C2 => n170
                           , A => n3681, ZN => n3678);
   U4517 : OAI22_X1 port map( A1 => n434, A2 => n3306, B1 => n74, B2 => n3307, 
                           ZN => n3681);
   U4518 : AOI221_X1 port map( B1 => n3308, B2 => n6360, C1 => n3309, C2 => 
                           n6392, A => n3682, ZN => n3677);
   U4519 : OAI222_X1 port map( A1 => n5176, A2 => n3311, B1 => n5144, B2 => 
                           n3312, C1 => n5112, C2 => n422, ZN => n3682);
   U4520 : AOI221_X1 port map( B1 => n3313, B2 => n571, C1 => n3314, C2 => n115
                           , A => n3683, ZN => n3676);
   U4521 : OAI22_X1 port map( A1 => n19, A2 => n415, B1 => n475, B2 => n3316, 
                           ZN => n3683);
   U4522 : NAND4_X1 port map( A1 => n3684, A2 => n3685, A3 => n3686, A4 => 
                           n3687, ZN => n3665);
   U4523 : AOI221_X1 port map( B1 => n3321, B2 => n6104, C1 => n3322, C2 => 
                           n6136, A => n3688, ZN => n3687);
   U4524 : OAI222_X1 port map( A1 => n4888, A2 => n3324, B1 => n4856, B2 => 
                           n3325, C1 => n4824, C2 => n423, ZN => n3688);
   U4525 : AOI221_X1 port map( B1 => n3326, B2 => n742, C1 => n3327, C2 => n318
                           , A => n3689, ZN => n3686);
   U4526 : OAI22_X1 port map( A1 => n222, A2 => n3329, B1 => n646, B2 => n3330,
                           ZN => n3689);
   U4527 : AOI221_X1 port map( B1 => n3331, B2 => n6232, C1 => n3332, C2 => 
                           n6264, A => n3690, ZN => n3685);
   U4528 : OAI222_X1 port map( A1 => n4984, A2 => n3334, B1 => n4952, B2 => 
                           n3335, C1 => n4920, C2 => n3336, ZN => n3690);
   U4529 : AOI221_X1 port map( B1 => n3337, B2 => n572, C1 => n3338, C2 => n116
                           , A => n3691, ZN => n3684);
   U4530 : OAI22_X1 port map( A1 => n20, A2 => n3340, B1 => n476, B2 => n3341, 
                           ZN => n3691);
   U4531 : NAND4_X1 port map( A1 => n3692, A2 => n3693, A3 => n3694, A4 => 
                           n3695, ZN => n3664);
   U4532 : AOI221_X1 port map( B1 => n3346, B2 => n5848, C1 => n3347, C2 => 
                           n5880, A => n3696, ZN => n3695);
   U4533 : OAI222_X1 port map( A1 => n4632, A2 => n3349, B1 => n4600, B2 => 
                           n3350, C1 => n4568, C2 => n3351, ZN => n3696);
   U4534 : AOI221_X1 port map( B1 => n3352, B2 => n5912, C1 => n3353, C2 => 
                           n5944, A => n3697, ZN => n3694);
   U4535 : OAI22_X1 port map( A1 => n4696, A2 => n3355, B1 => n4664, B2 => 
                           n3356, ZN => n3697);
   U4536 : AOI221_X1 port map( B1 => n3357, B2 => n5976, C1 => n3358, C2 => 
                           n6008, A => n3698, ZN => n3693);
   U4537 : OAI222_X1 port map( A1 => n4792, A2 => n3360, B1 => n4760, B2 => 
                           n3361, C1 => n4728, C2 => n424, ZN => n3698);
   U4538 : AOI221_X1 port map( B1 => n3362, B2 => n6072, C1 => n3363, C2 => 
                           n6040, A => n3699, ZN => n3692);
   U4539 : OAI22_X1 port map( A1 => n5599, A2 => n3365, B1 => n5598, B2 => 
                           n3366, ZN => n3699);
   U4540 : INV_X1 port map( A => DATAIN(22), ZN => n2356);
   U4541 : OAI21_X1 port map( B1 => n3266, B2 => n1554, A => ENABLE, ZN => 
                           n7590);
   U4542 : OAI222_X1 port map( A1 => n2394, A2 => n3263, B1 => n3700, B2 => 
                           n3265, C1 => n3266, C2 => n1491, ZN => n7589);
   U4543 : NOR4_X1 port map( A1 => n3701, A2 => n3702, A3 => n3703, A4 => n3704
                           , ZN => n3700);
   U4544 : NAND4_X1 port map( A1 => n3705, A2 => n3706, A3 => n3707, A4 => 
                           n3708, ZN => n3704);
   U4545 : AOI221_X1 port map( B1 => n3275, B2 => n6423, C1 => n3276, C2 => 
                           n6455, A => n3709, ZN => n3708);
   U4546 : OAI222_X1 port map( A1 => n5271, A2 => n3278, B1 => n5239, B2 => 
                           n3279, C1 => n5207, C2 => n421, ZN => n3709);
   U4547 : AOI221_X1 port map( B1 => n3280, B2 => n743, C1 => n3281, C2 => n319
                           , A => n3710, ZN => n3707);
   U4548 : OAI22_X1 port map( A1 => n223, A2 => n413, B1 => n647, B2 => n3283, 
                           ZN => n3710);
   U4549 : AOI221_X1 port map( B1 => n3284, B2 => n6551, C1 => n3285, C2 => 
                           n6583, A => n3711, ZN => n3706);
   U4550 : OAI222_X1 port map( A1 => n5367, A2 => n3287, B1 => n5335, B2 => 
                           n1579, C1 => n5303, C2 => n3288, ZN => n3711);
   U4551 : AOI221_X1 port map( B1 => n3289, B2 => n744, C1 => n3290, C2 => n320
                           , A => n3712, ZN => n3705);
   U4552 : OAI22_X1 port map( A1 => n224, A2 => n414, B1 => n648, B2 => n3292, 
                           ZN => n3712);
   U4553 : NAND4_X1 port map( A1 => n3713, A2 => n3714, A3 => n3715, A4 => 
                           n3716, ZN => n3703);
   U4554 : AOI221_X1 port map( B1 => n3297, B2 => n6295, C1 => n3298, C2 => 
                           n6327, A => n3717, ZN => n3716);
   U4555 : OAI222_X1 port map( A1 => n5079, A2 => n3300, B1 => n5047, B2 => 
                           n3301, C1 => n5015, C2 => n3302, ZN => n3717);
   U4556 : AOI221_X1 port map( B1 => n3303, B2 => n531, C1 => n3304, C2 => n171
                           , A => n3718, ZN => n3715);
   U4557 : OAI22_X1 port map( A1 => n435, A2 => n3306, B1 => n75, B2 => n3307, 
                           ZN => n3718);
   U4558 : AOI221_X1 port map( B1 => n3308, B2 => n6359, C1 => n3309, C2 => 
                           n6391, A => n3719, ZN => n3714);
   U4559 : OAI222_X1 port map( A1 => n5175, A2 => n3311, B1 => n5143, B2 => 
                           n3312, C1 => n5111, C2 => n422, ZN => n3719);
   U4560 : AOI221_X1 port map( B1 => n3313, B2 => n573, C1 => n3314, C2 => n117
                           , A => n3720, ZN => n3713);
   U4561 : OAI22_X1 port map( A1 => n21, A2 => n415, B1 => n477, B2 => n3316, 
                           ZN => n3720);
   U4562 : NAND4_X1 port map( A1 => n3721, A2 => n3722, A3 => n3723, A4 => 
                           n3724, ZN => n3702);
   U4563 : AOI221_X1 port map( B1 => n3321, B2 => n6103, C1 => n3322, C2 => 
                           n6135, A => n3725, ZN => n3724);
   U4564 : OAI222_X1 port map( A1 => n4887, A2 => n3324, B1 => n4855, B2 => 
                           n3325, C1 => n4823, C2 => n423, ZN => n3725);
   U4565 : AOI221_X1 port map( B1 => n3326, B2 => n745, C1 => n3327, C2 => n321
                           , A => n3726, ZN => n3723);
   U4566 : OAI22_X1 port map( A1 => n225, A2 => n3329, B1 => n649, B2 => n3330,
                           ZN => n3726);
   U4567 : AOI221_X1 port map( B1 => n3331, B2 => n6231, C1 => n3332, C2 => 
                           n6263, A => n3727, ZN => n3722);
   U4568 : OAI222_X1 port map( A1 => n4983, A2 => n3334, B1 => n4951, B2 => 
                           n3335, C1 => n4919, C2 => n3336, ZN => n3727);
   U4569 : AOI221_X1 port map( B1 => n3337, B2 => n574, C1 => n3338, C2 => n118
                           , A => n3728, ZN => n3721);
   U4570 : OAI22_X1 port map( A1 => n22, A2 => n3340, B1 => n478, B2 => n3341, 
                           ZN => n3728);
   U4571 : NAND4_X1 port map( A1 => n3729, A2 => n3730, A3 => n3731, A4 => 
                           n3732, ZN => n3701);
   U4572 : AOI221_X1 port map( B1 => n3346, B2 => n5847, C1 => n3347, C2 => 
                           n5879, A => n3733, ZN => n3732);
   U4573 : OAI222_X1 port map( A1 => n4631, A2 => n3349, B1 => n4599, B2 => 
                           n3350, C1 => n4567, C2 => n3351, ZN => n3733);
   U4574 : AOI221_X1 port map( B1 => n3352, B2 => n5911, C1 => n3353, C2 => 
                           n5943, A => n3734, ZN => n3731);
   U4575 : OAI22_X1 port map( A1 => n4695, A2 => n3355, B1 => n4663, B2 => 
                           n3356, ZN => n3734);
   U4576 : AOI221_X1 port map( B1 => n3357, B2 => n5975, C1 => n3358, C2 => 
                           n6007, A => n3735, ZN => n3730);
   U4577 : OAI222_X1 port map( A1 => n4791, A2 => n3360, B1 => n4759, B2 => 
                           n3361, C1 => n4727, C2 => n424, ZN => n3735);
   U4578 : AOI221_X1 port map( B1 => n3362, B2 => n6071, C1 => n3363, C2 => 
                           n6039, A => n3736, ZN => n3729);
   U4579 : OAI22_X1 port map( A1 => n5589, A2 => n3365, B1 => n5588, B2 => 
                           n3366, ZN => n3736);
   U4580 : INV_X1 port map( A => DATAIN(21), ZN => n2394);
   U4581 : OAI21_X1 port map( B1 => n3266, B2 => n1555, A => ENABLE, ZN => 
                           n7588);
   U4582 : OAI222_X1 port map( A1 => n2432, A2 => n3263, B1 => n3737, B2 => 
                           n3265, C1 => n3266, C2 => n1492, ZN => n7587);
   U4583 : NOR4_X1 port map( A1 => n3738, A2 => n3739, A3 => n3740, A4 => n3741
                           , ZN => n3737);
   U4584 : NAND4_X1 port map( A1 => n3742, A2 => n3743, A3 => n3744, A4 => 
                           n3745, ZN => n3741);
   U4585 : AOI221_X1 port map( B1 => n3275, B2 => n6422, C1 => n3276, C2 => 
                           n6454, A => n3746, ZN => n3745);
   U4586 : OAI222_X1 port map( A1 => n5270, A2 => n3278, B1 => n5238, B2 => 
                           n3279, C1 => n5206, C2 => n421, ZN => n3746);
   U4587 : AOI221_X1 port map( B1 => n3280, B2 => n746, C1 => n3281, C2 => n322
                           , A => n3747, ZN => n3744);
   U4588 : OAI22_X1 port map( A1 => n226, A2 => n413, B1 => n650, B2 => n3283, 
                           ZN => n3747);
   U4589 : AOI221_X1 port map( B1 => n3284, B2 => n6550, C1 => n3285, C2 => 
                           n6582, A => n3748, ZN => n3743);
   U4590 : OAI222_X1 port map( A1 => n5366, A2 => n3287, B1 => n5334, B2 => 
                           n1579, C1 => n5302, C2 => n3288, ZN => n3748);
   U4591 : AOI221_X1 port map( B1 => n3289, B2 => n747, C1 => n3290, C2 => n323
                           , A => n3749, ZN => n3742);
   U4592 : OAI22_X1 port map( A1 => n227, A2 => n414, B1 => n651, B2 => n3292, 
                           ZN => n3749);
   U4593 : NAND4_X1 port map( A1 => n3750, A2 => n3751, A3 => n3752, A4 => 
                           n3753, ZN => n3740);
   U4594 : AOI221_X1 port map( B1 => n3297, B2 => n6294, C1 => n3298, C2 => 
                           n6326, A => n3754, ZN => n3753);
   U4595 : OAI222_X1 port map( A1 => n5078, A2 => n3300, B1 => n5046, B2 => 
                           n3301, C1 => n5014, C2 => n3302, ZN => n3754);
   U4596 : AOI221_X1 port map( B1 => n3303, B2 => n532, C1 => n3304, C2 => n172
                           , A => n3755, ZN => n3752);
   U4597 : OAI22_X1 port map( A1 => n436, A2 => n3306, B1 => n76, B2 => n3307, 
                           ZN => n3755);
   U4598 : AOI221_X1 port map( B1 => n3308, B2 => n6358, C1 => n3309, C2 => 
                           n6390, A => n3756, ZN => n3751);
   U4599 : OAI222_X1 port map( A1 => n5174, A2 => n3311, B1 => n5142, B2 => 
                           n3312, C1 => n5110, C2 => n422, ZN => n3756);
   U4600 : AOI221_X1 port map( B1 => n3313, B2 => n575, C1 => n3314, C2 => n119
                           , A => n3757, ZN => n3750);
   U4601 : OAI22_X1 port map( A1 => n23, A2 => n415, B1 => n479, B2 => n3316, 
                           ZN => n3757);
   U4602 : NAND4_X1 port map( A1 => n3758, A2 => n3759, A3 => n3760, A4 => 
                           n3761, ZN => n3739);
   U4603 : AOI221_X1 port map( B1 => n3321, B2 => n6102, C1 => n3322, C2 => 
                           n6134, A => n3762, ZN => n3761);
   U4604 : OAI222_X1 port map( A1 => n4886, A2 => n3324, B1 => n4854, B2 => 
                           n3325, C1 => n4822, C2 => n423, ZN => n3762);
   U4605 : AOI221_X1 port map( B1 => n3326, B2 => n748, C1 => n3327, C2 => n324
                           , A => n3763, ZN => n3760);
   U4606 : OAI22_X1 port map( A1 => n228, A2 => n3329, B1 => n652, B2 => n3330,
                           ZN => n3763);
   U4607 : AOI221_X1 port map( B1 => n3331, B2 => n6230, C1 => n3332, C2 => 
                           n6262, A => n3764, ZN => n3759);
   U4608 : OAI222_X1 port map( A1 => n4982, A2 => n3334, B1 => n4950, B2 => 
                           n3335, C1 => n4918, C2 => n3336, ZN => n3764);
   U4609 : AOI221_X1 port map( B1 => n3337, B2 => n576, C1 => n3338, C2 => n120
                           , A => n3765, ZN => n3758);
   U4610 : OAI22_X1 port map( A1 => n24, A2 => n3340, B1 => n480, B2 => n3341, 
                           ZN => n3765);
   U4611 : NAND4_X1 port map( A1 => n3766, A2 => n3767, A3 => n3768, A4 => 
                           n3769, ZN => n3738);
   U4612 : AOI221_X1 port map( B1 => n3346, B2 => n5846, C1 => n3347, C2 => 
                           n5878, A => n3770, ZN => n3769);
   U4613 : OAI222_X1 port map( A1 => n4630, A2 => n3349, B1 => n4598, B2 => 
                           n3350, C1 => n4566, C2 => n3351, ZN => n3770);
   U4614 : AOI221_X1 port map( B1 => n3352, B2 => n5910, C1 => n3353, C2 => 
                           n5942, A => n3771, ZN => n3768);
   U4615 : OAI22_X1 port map( A1 => n4694, A2 => n3355, B1 => n4662, B2 => 
                           n3356, ZN => n3771);
   U4616 : AOI221_X1 port map( B1 => n3357, B2 => n5974, C1 => n3358, C2 => 
                           n6006, A => n3772, ZN => n3767);
   U4617 : OAI222_X1 port map( A1 => n4790, A2 => n3360, B1 => n4758, B2 => 
                           n3361, C1 => n4726, C2 => n424, ZN => n3772);
   U4618 : AOI221_X1 port map( B1 => n3362, B2 => n6070, C1 => n3363, C2 => 
                           n6038, A => n3773, ZN => n3766);
   U4619 : OAI22_X1 port map( A1 => n5579, A2 => n3365, B1 => n5578, B2 => 
                           n3366, ZN => n3773);
   U4620 : INV_X1 port map( A => DATAIN(20), ZN => n2432);
   U4621 : OAI21_X1 port map( B1 => n3266, B2 => n1556, A => ENABLE, ZN => 
                           n7586);
   U4622 : OAI222_X1 port map( A1 => n2470, A2 => n3263, B1 => n3774, B2 => 
                           n3265, C1 => n3266, C2 => n1493, ZN => n7585);
   U4623 : NOR4_X1 port map( A1 => n3775, A2 => n3776, A3 => n3777, A4 => n3778
                           , ZN => n3774);
   U4624 : NAND4_X1 port map( A1 => n3779, A2 => n3780, A3 => n3781, A4 => 
                           n3782, ZN => n3778);
   U4625 : AOI221_X1 port map( B1 => n3275, B2 => n6421, C1 => n3276, C2 => 
                           n6453, A => n3783, ZN => n3782);
   U4626 : OAI222_X1 port map( A1 => n5269, A2 => n3278, B1 => n5237, B2 => 
                           n3279, C1 => n5205, C2 => n421, ZN => n3783);
   U4627 : AOI221_X1 port map( B1 => n3280, B2 => n749, C1 => n3281, C2 => n325
                           , A => n3784, ZN => n3781);
   U4628 : OAI22_X1 port map( A1 => n229, A2 => n413, B1 => n653, B2 => n3283, 
                           ZN => n3784);
   U4629 : AOI221_X1 port map( B1 => n3284, B2 => n6549, C1 => n3285, C2 => 
                           n6581, A => n3785, ZN => n3780);
   U4630 : OAI222_X1 port map( A1 => n5365, A2 => n3287, B1 => n5333, B2 => 
                           n1579, C1 => n5301, C2 => n3288, ZN => n3785);
   U4631 : AOI221_X1 port map( B1 => n3289, B2 => n750, C1 => n3290, C2 => n326
                           , A => n3786, ZN => n3779);
   U4632 : OAI22_X1 port map( A1 => n230, A2 => n414, B1 => n654, B2 => n3292, 
                           ZN => n3786);
   U4633 : NAND4_X1 port map( A1 => n3787, A2 => n3788, A3 => n3789, A4 => 
                           n3790, ZN => n3777);
   U4634 : AOI221_X1 port map( B1 => n3297, B2 => n6293, C1 => n3298, C2 => 
                           n6325, A => n3791, ZN => n3790);
   U4635 : OAI222_X1 port map( A1 => n5077, A2 => n3300, B1 => n5045, B2 => 
                           n3301, C1 => n5013, C2 => n3302, ZN => n3791);
   U4636 : AOI221_X1 port map( B1 => n3303, B2 => n533, C1 => n3304, C2 => n173
                           , A => n3792, ZN => n3789);
   U4637 : OAI22_X1 port map( A1 => n437, A2 => n3306, B1 => n77, B2 => n3307, 
                           ZN => n3792);
   U4638 : AOI221_X1 port map( B1 => n3308, B2 => n6357, C1 => n3309, C2 => 
                           n6389, A => n3793, ZN => n3788);
   U4639 : OAI222_X1 port map( A1 => n5173, A2 => n3311, B1 => n5141, B2 => 
                           n3312, C1 => n5109, C2 => n422, ZN => n3793);
   U4640 : AOI221_X1 port map( B1 => n3313, B2 => n577, C1 => n3314, C2 => n121
                           , A => n3794, ZN => n3787);
   U4641 : OAI22_X1 port map( A1 => n25, A2 => n415, B1 => n481, B2 => n3316, 
                           ZN => n3794);
   U4642 : NAND4_X1 port map( A1 => n3795, A2 => n3796, A3 => n3797, A4 => 
                           n3798, ZN => n3776);
   U4643 : AOI221_X1 port map( B1 => n3321, B2 => n6101, C1 => n3322, C2 => 
                           n6133, A => n3799, ZN => n3798);
   U4644 : OAI222_X1 port map( A1 => n4885, A2 => n3324, B1 => n4853, B2 => 
                           n3325, C1 => n4821, C2 => n423, ZN => n3799);
   U4645 : AOI221_X1 port map( B1 => n3326, B2 => n751, C1 => n3327, C2 => n327
                           , A => n3800, ZN => n3797);
   U4646 : OAI22_X1 port map( A1 => n231, A2 => n3329, B1 => n655, B2 => n3330,
                           ZN => n3800);
   U4647 : AOI221_X1 port map( B1 => n3331, B2 => n6229, C1 => n3332, C2 => 
                           n6261, A => n3801, ZN => n3796);
   U4648 : OAI222_X1 port map( A1 => n4981, A2 => n3334, B1 => n4949, B2 => 
                           n3335, C1 => n4917, C2 => n3336, ZN => n3801);
   U4649 : AOI221_X1 port map( B1 => n3337, B2 => n578, C1 => n3338, C2 => n122
                           , A => n3802, ZN => n3795);
   U4650 : OAI22_X1 port map( A1 => n26, A2 => n3340, B1 => n482, B2 => n3341, 
                           ZN => n3802);
   U4651 : NAND4_X1 port map( A1 => n3803, A2 => n3804, A3 => n3805, A4 => 
                           n3806, ZN => n3775);
   U4652 : AOI221_X1 port map( B1 => n3346, B2 => n5845, C1 => n3347, C2 => 
                           n5877, A => n3807, ZN => n3806);
   U4653 : OAI222_X1 port map( A1 => n4629, A2 => n3349, B1 => n4597, B2 => 
                           n3350, C1 => n4565, C2 => n3351, ZN => n3807);
   U4654 : AOI221_X1 port map( B1 => n3352, B2 => n5909, C1 => n3353, C2 => 
                           n5941, A => n3808, ZN => n3805);
   U4655 : OAI22_X1 port map( A1 => n4693, A2 => n3355, B1 => n4661, B2 => 
                           n3356, ZN => n3808);
   U4656 : AOI221_X1 port map( B1 => n3357, B2 => n5973, C1 => n3358, C2 => 
                           n6005, A => n3809, ZN => n3804);
   U4657 : OAI222_X1 port map( A1 => n4789, A2 => n3360, B1 => n4757, B2 => 
                           n3361, C1 => n4725, C2 => n424, ZN => n3809);
   U4658 : AOI221_X1 port map( B1 => n3362, B2 => n6069, C1 => n3363, C2 => 
                           n6037, A => n3810, ZN => n3803);
   U4659 : OAI22_X1 port map( A1 => n5569, A2 => n3365, B1 => n5568, B2 => 
                           n3366, ZN => n3810);
   U4660 : INV_X1 port map( A => DATAIN(19), ZN => n2470);
   U4661 : OAI21_X1 port map( B1 => n3266, B2 => n1557, A => ENABLE, ZN => 
                           n7584);
   U4662 : OAI222_X1 port map( A1 => n2508, A2 => n3263, B1 => n3811, B2 => 
                           n3265, C1 => n3266, C2 => n1494, ZN => n7583);
   U4663 : NOR4_X1 port map( A1 => n3812, A2 => n3813, A3 => n3814, A4 => n3815
                           , ZN => n3811);
   U4664 : NAND4_X1 port map( A1 => n3816, A2 => n3817, A3 => n3818, A4 => 
                           n3819, ZN => n3815);
   U4665 : AOI221_X1 port map( B1 => n3275, B2 => n6420, C1 => n3276, C2 => 
                           n6452, A => n3820, ZN => n3819);
   U4666 : OAI222_X1 port map( A1 => n5268, A2 => n3278, B1 => n5236, B2 => 
                           n3279, C1 => n5204, C2 => n421, ZN => n3820);
   U4667 : AOI221_X1 port map( B1 => n3280, B2 => n752, C1 => n3281, C2 => n328
                           , A => n3821, ZN => n3818);
   U4668 : OAI22_X1 port map( A1 => n232, A2 => n413, B1 => n656, B2 => n3283, 
                           ZN => n3821);
   U4669 : AOI221_X1 port map( B1 => n3284, B2 => n6548, C1 => n3285, C2 => 
                           n6580, A => n3822, ZN => n3817);
   U4670 : OAI222_X1 port map( A1 => n5364, A2 => n3287, B1 => n5332, B2 => 
                           n1579, C1 => n5300, C2 => n3288, ZN => n3822);
   U4671 : AOI221_X1 port map( B1 => n3289, B2 => n753, C1 => n3290, C2 => n329
                           , A => n3823, ZN => n3816);
   U4672 : OAI22_X1 port map( A1 => n233, A2 => n414, B1 => n657, B2 => n3292, 
                           ZN => n3823);
   U4673 : NAND4_X1 port map( A1 => n3824, A2 => n3825, A3 => n3826, A4 => 
                           n3827, ZN => n3814);
   U4674 : AOI221_X1 port map( B1 => n3297, B2 => n6292, C1 => n3298, C2 => 
                           n6324, A => n3828, ZN => n3827);
   U4675 : OAI222_X1 port map( A1 => n5076, A2 => n3300, B1 => n5044, B2 => 
                           n3301, C1 => n5012, C2 => n3302, ZN => n3828);
   U4676 : AOI221_X1 port map( B1 => n3303, B2 => n534, C1 => n3304, C2 => n174
                           , A => n3829, ZN => n3826);
   U4677 : OAI22_X1 port map( A1 => n438, A2 => n3306, B1 => n78, B2 => n3307, 
                           ZN => n3829);
   U4678 : AOI221_X1 port map( B1 => n3308, B2 => n6356, C1 => n3309, C2 => 
                           n6388, A => n3830, ZN => n3825);
   U4679 : OAI222_X1 port map( A1 => n5172, A2 => n3311, B1 => n5140, B2 => 
                           n3312, C1 => n5108, C2 => n422, ZN => n3830);
   U4680 : AOI221_X1 port map( B1 => n3313, B2 => n579, C1 => n3314, C2 => n123
                           , A => n3831, ZN => n3824);
   U4681 : OAI22_X1 port map( A1 => n27, A2 => n415, B1 => n483, B2 => n3316, 
                           ZN => n3831);
   U4682 : NAND4_X1 port map( A1 => n3832, A2 => n3833, A3 => n3834, A4 => 
                           n3835, ZN => n3813);
   U4683 : AOI221_X1 port map( B1 => n3321, B2 => n6100, C1 => n3322, C2 => 
                           n6132, A => n3836, ZN => n3835);
   U4684 : OAI222_X1 port map( A1 => n4884, A2 => n3324, B1 => n4852, B2 => 
                           n3325, C1 => n4820, C2 => n423, ZN => n3836);
   U4685 : AOI221_X1 port map( B1 => n3326, B2 => n754, C1 => n3327, C2 => n330
                           , A => n3837, ZN => n3834);
   U4686 : OAI22_X1 port map( A1 => n234, A2 => n3329, B1 => n658, B2 => n3330,
                           ZN => n3837);
   U4687 : AOI221_X1 port map( B1 => n3331, B2 => n6228, C1 => n3332, C2 => 
                           n6260, A => n3838, ZN => n3833);
   U4688 : OAI222_X1 port map( A1 => n4980, A2 => n3334, B1 => n4948, B2 => 
                           n3335, C1 => n4916, C2 => n3336, ZN => n3838);
   U4689 : AOI221_X1 port map( B1 => n3337, B2 => n580, C1 => n3338, C2 => n124
                           , A => n3839, ZN => n3832);
   U4690 : OAI22_X1 port map( A1 => n28, A2 => n3340, B1 => n484, B2 => n3341, 
                           ZN => n3839);
   U4691 : NAND4_X1 port map( A1 => n3840, A2 => n3841, A3 => n3842, A4 => 
                           n3843, ZN => n3812);
   U4692 : AOI221_X1 port map( B1 => n3346, B2 => n5844, C1 => n3347, C2 => 
                           n5876, A => n3844, ZN => n3843);
   U4693 : OAI222_X1 port map( A1 => n4628, A2 => n3349, B1 => n4596, B2 => 
                           n3350, C1 => n4564, C2 => n3351, ZN => n3844);
   U4694 : AOI221_X1 port map( B1 => n3352, B2 => n5908, C1 => n3353, C2 => 
                           n5940, A => n3845, ZN => n3842);
   U4695 : OAI22_X1 port map( A1 => n4692, A2 => n3355, B1 => n4660, B2 => 
                           n3356, ZN => n3845);
   U4696 : AOI221_X1 port map( B1 => n3357, B2 => n5972, C1 => n3358, C2 => 
                           n6004, A => n3846, ZN => n3841);
   U4697 : OAI222_X1 port map( A1 => n4788, A2 => n3360, B1 => n4756, B2 => 
                           n3361, C1 => n4724, C2 => n424, ZN => n3846);
   U4698 : AOI221_X1 port map( B1 => n3362, B2 => n6068, C1 => n3363, C2 => 
                           n6036, A => n3847, ZN => n3840);
   U4699 : OAI22_X1 port map( A1 => n5559, A2 => n3365, B1 => n5558, B2 => 
                           n3366, ZN => n3847);
   U4700 : INV_X1 port map( A => DATAIN(18), ZN => n2508);
   U4701 : OAI21_X1 port map( B1 => n3266, B2 => n1558, A => ENABLE, ZN => 
                           n7582);
   U4702 : OAI222_X1 port map( A1 => n2546, A2 => n3263, B1 => n3848, B2 => 
                           n3265, C1 => n3266, C2 => n1495, ZN => n7581);
   U4703 : NOR4_X1 port map( A1 => n3849, A2 => n3850, A3 => n3851, A4 => n3852
                           , ZN => n3848);
   U4704 : NAND4_X1 port map( A1 => n3853, A2 => n3854, A3 => n3855, A4 => 
                           n3856, ZN => n3852);
   U4705 : AOI221_X1 port map( B1 => n3275, B2 => n6419, C1 => n3276, C2 => 
                           n6451, A => n3857, ZN => n3856);
   U4706 : OAI222_X1 port map( A1 => n5267, A2 => n3278, B1 => n5235, B2 => 
                           n3279, C1 => n5203, C2 => n421, ZN => n3857);
   U4707 : AOI221_X1 port map( B1 => n3280, B2 => n755, C1 => n3281, C2 => n331
                           , A => n3858, ZN => n3855);
   U4708 : OAI22_X1 port map( A1 => n235, A2 => n413, B1 => n659, B2 => n3283, 
                           ZN => n3858);
   U4709 : AOI221_X1 port map( B1 => n3284, B2 => n6547, C1 => n3285, C2 => 
                           n6579, A => n3859, ZN => n3854);
   U4710 : OAI222_X1 port map( A1 => n5363, A2 => n3287, B1 => n5331, B2 => 
                           n1579, C1 => n5299, C2 => n3288, ZN => n3859);
   U4711 : AOI221_X1 port map( B1 => n3289, B2 => n756, C1 => n3290, C2 => n332
                           , A => n3860, ZN => n3853);
   U4712 : OAI22_X1 port map( A1 => n236, A2 => n414, B1 => n660, B2 => n3292, 
                           ZN => n3860);
   U4713 : NAND4_X1 port map( A1 => n3861, A2 => n3862, A3 => n3863, A4 => 
                           n3864, ZN => n3851);
   U4714 : AOI221_X1 port map( B1 => n3297, B2 => n6291, C1 => n3298, C2 => 
                           n6323, A => n3865, ZN => n3864);
   U4715 : OAI222_X1 port map( A1 => n5075, A2 => n3300, B1 => n5043, B2 => 
                           n3301, C1 => n5011, C2 => n3302, ZN => n3865);
   U4716 : AOI221_X1 port map( B1 => n3303, B2 => n535, C1 => n3304, C2 => n175
                           , A => n3866, ZN => n3863);
   U4717 : OAI22_X1 port map( A1 => n439, A2 => n3306, B1 => n79, B2 => n3307, 
                           ZN => n3866);
   U4718 : AOI221_X1 port map( B1 => n3308, B2 => n6355, C1 => n3309, C2 => 
                           n6387, A => n3867, ZN => n3862);
   U4719 : OAI222_X1 port map( A1 => n5171, A2 => n3311, B1 => n5139, B2 => 
                           n3312, C1 => n5107, C2 => n422, ZN => n3867);
   U4720 : AOI221_X1 port map( B1 => n3313, B2 => n581, C1 => n3314, C2 => n125
                           , A => n3868, ZN => n3861);
   U4721 : OAI22_X1 port map( A1 => n29, A2 => n415, B1 => n485, B2 => n3316, 
                           ZN => n3868);
   U4722 : NAND4_X1 port map( A1 => n3869, A2 => n3870, A3 => n3871, A4 => 
                           n3872, ZN => n3850);
   U4723 : AOI221_X1 port map( B1 => n3321, B2 => n6099, C1 => n3322, C2 => 
                           n6131, A => n3873, ZN => n3872);
   U4724 : OAI222_X1 port map( A1 => n4883, A2 => n3324, B1 => n4851, B2 => 
                           n3325, C1 => n4819, C2 => n423, ZN => n3873);
   U4725 : AOI221_X1 port map( B1 => n3326, B2 => n757, C1 => n3327, C2 => n333
                           , A => n3874, ZN => n3871);
   U4726 : OAI22_X1 port map( A1 => n237, A2 => n3329, B1 => n661, B2 => n3330,
                           ZN => n3874);
   U4727 : AOI221_X1 port map( B1 => n3331, B2 => n6227, C1 => n3332, C2 => 
                           n6259, A => n3875, ZN => n3870);
   U4728 : OAI222_X1 port map( A1 => n4979, A2 => n3334, B1 => n4947, B2 => 
                           n3335, C1 => n4915, C2 => n3336, ZN => n3875);
   U4729 : AOI221_X1 port map( B1 => n3337, B2 => n582, C1 => n3338, C2 => n126
                           , A => n3876, ZN => n3869);
   U4730 : OAI22_X1 port map( A1 => n30, A2 => n3340, B1 => n486, B2 => n3341, 
                           ZN => n3876);
   U4731 : NAND4_X1 port map( A1 => n3877, A2 => n3878, A3 => n3879, A4 => 
                           n3880, ZN => n3849);
   U4732 : AOI221_X1 port map( B1 => n3346, B2 => n5843, C1 => n3347, C2 => 
                           n5875, A => n3881, ZN => n3880);
   U4733 : OAI222_X1 port map( A1 => n4627, A2 => n3349, B1 => n4595, B2 => 
                           n3350, C1 => n4563, C2 => n3351, ZN => n3881);
   U4734 : AOI221_X1 port map( B1 => n3352, B2 => n5907, C1 => n3353, C2 => 
                           n5939, A => n3882, ZN => n3879);
   U4735 : OAI22_X1 port map( A1 => n4691, A2 => n3355, B1 => n4659, B2 => 
                           n3356, ZN => n3882);
   U4736 : AOI221_X1 port map( B1 => n3357, B2 => n5971, C1 => n3358, C2 => 
                           n6003, A => n3883, ZN => n3878);
   U4737 : OAI222_X1 port map( A1 => n4787, A2 => n3360, B1 => n4755, B2 => 
                           n3361, C1 => n4723, C2 => n424, ZN => n3883);
   U4738 : AOI221_X1 port map( B1 => n3362, B2 => n6067, C1 => n3363, C2 => 
                           n6035, A => n3884, ZN => n3877);
   U4739 : OAI22_X1 port map( A1 => n5549, A2 => n3365, B1 => n5548, B2 => 
                           n3366, ZN => n3884);
   U4740 : INV_X1 port map( A => DATAIN(17), ZN => n2546);
   U4741 : OAI21_X1 port map( B1 => n3266, B2 => n1559, A => ENABLE, ZN => 
                           n7580);
   U4742 : OAI222_X1 port map( A1 => n2584, A2 => n3263, B1 => n3885, B2 => 
                           n3265, C1 => n3266, C2 => n1496, ZN => n7579);
   U4743 : NOR4_X1 port map( A1 => n3886, A2 => n3887, A3 => n3888, A4 => n3889
                           , ZN => n3885);
   U4744 : NAND4_X1 port map( A1 => n3890, A2 => n3891, A3 => n3892, A4 => 
                           n3893, ZN => n3889);
   U4745 : AOI221_X1 port map( B1 => n3275, B2 => n6418, C1 => n3276, C2 => 
                           n6450, A => n3894, ZN => n3893);
   U4746 : OAI222_X1 port map( A1 => n5266, A2 => n3278, B1 => n5234, B2 => 
                           n3279, C1 => n5202, C2 => n421, ZN => n3894);
   U4747 : AOI221_X1 port map( B1 => n3280, B2 => n758, C1 => n3281, C2 => n334
                           , A => n3895, ZN => n3892);
   U4748 : OAI22_X1 port map( A1 => n238, A2 => n413, B1 => n662, B2 => n3283, 
                           ZN => n3895);
   U4749 : AOI221_X1 port map( B1 => n3284, B2 => n6546, C1 => n3285, C2 => 
                           n6578, A => n3896, ZN => n3891);
   U4750 : OAI222_X1 port map( A1 => n5362, A2 => n3287, B1 => n5330, B2 => 
                           n1579, C1 => n5298, C2 => n3288, ZN => n3896);
   U4751 : AOI221_X1 port map( B1 => n3289, B2 => n759, C1 => n3290, C2 => n335
                           , A => n3897, ZN => n3890);
   U4752 : OAI22_X1 port map( A1 => n239, A2 => n414, B1 => n663, B2 => n3292, 
                           ZN => n3897);
   U4753 : NAND4_X1 port map( A1 => n3898, A2 => n3899, A3 => n3900, A4 => 
                           n3901, ZN => n3888);
   U4754 : AOI221_X1 port map( B1 => n3297, B2 => n6290, C1 => n3298, C2 => 
                           n6322, A => n3902, ZN => n3901);
   U4755 : OAI222_X1 port map( A1 => n5074, A2 => n3300, B1 => n5042, B2 => 
                           n3301, C1 => n5010, C2 => n3302, ZN => n3902);
   U4756 : AOI221_X1 port map( B1 => n3303, B2 => n536, C1 => n3304, C2 => n176
                           , A => n3903, ZN => n3900);
   U4757 : OAI22_X1 port map( A1 => n440, A2 => n3306, B1 => n80, B2 => n3307, 
                           ZN => n3903);
   U4758 : AOI221_X1 port map( B1 => n3308, B2 => n6354, C1 => n3309, C2 => 
                           n6386, A => n3904, ZN => n3899);
   U4759 : OAI222_X1 port map( A1 => n5170, A2 => n3311, B1 => n5138, B2 => 
                           n3312, C1 => n5106, C2 => n422, ZN => n3904);
   U4760 : AOI221_X1 port map( B1 => n3313, B2 => n583, C1 => n3314, C2 => n127
                           , A => n3905, ZN => n3898);
   U4761 : OAI22_X1 port map( A1 => n31, A2 => n415, B1 => n487, B2 => n3316, 
                           ZN => n3905);
   U4762 : NAND4_X1 port map( A1 => n3906, A2 => n3907, A3 => n3908, A4 => 
                           n3909, ZN => n3887);
   U4763 : AOI221_X1 port map( B1 => n3321, B2 => n6098, C1 => n3322, C2 => 
                           n6130, A => n3910, ZN => n3909);
   U4764 : OAI222_X1 port map( A1 => n4882, A2 => n3324, B1 => n4850, B2 => 
                           n3325, C1 => n4818, C2 => n423, ZN => n3910);
   U4765 : AOI221_X1 port map( B1 => n3326, B2 => n760, C1 => n3327, C2 => n336
                           , A => n3911, ZN => n3908);
   U4766 : OAI22_X1 port map( A1 => n240, A2 => n3329, B1 => n664, B2 => n3330,
                           ZN => n3911);
   U4767 : AOI221_X1 port map( B1 => n3331, B2 => n6226, C1 => n3332, C2 => 
                           n6258, A => n3912, ZN => n3907);
   U4768 : OAI222_X1 port map( A1 => n4978, A2 => n3334, B1 => n4946, B2 => 
                           n3335, C1 => n4914, C2 => n3336, ZN => n3912);
   U4769 : AOI221_X1 port map( B1 => n3337, B2 => n584, C1 => n3338, C2 => n128
                           , A => n3913, ZN => n3906);
   U4770 : OAI22_X1 port map( A1 => n32, A2 => n3340, B1 => n488, B2 => n3341, 
                           ZN => n3913);
   U4771 : NAND4_X1 port map( A1 => n3914, A2 => n3915, A3 => n3916, A4 => 
                           n3917, ZN => n3886);
   U4772 : AOI221_X1 port map( B1 => n3346, B2 => n5842, C1 => n3347, C2 => 
                           n5874, A => n3918, ZN => n3917);
   U4773 : OAI222_X1 port map( A1 => n4626, A2 => n3349, B1 => n4594, B2 => 
                           n3350, C1 => n4562, C2 => n3351, ZN => n3918);
   U4774 : AOI221_X1 port map( B1 => n3352, B2 => n5906, C1 => n3353, C2 => 
                           n5938, A => n3919, ZN => n3916);
   U4775 : OAI22_X1 port map( A1 => n4690, A2 => n3355, B1 => n4658, B2 => 
                           n3356, ZN => n3919);
   U4776 : AOI221_X1 port map( B1 => n3357, B2 => n5970, C1 => n3358, C2 => 
                           n6002, A => n3920, ZN => n3915);
   U4777 : OAI222_X1 port map( A1 => n4786, A2 => n3360, B1 => n4754, B2 => 
                           n3361, C1 => n4722, C2 => n424, ZN => n3920);
   U4778 : AOI221_X1 port map( B1 => n3362, B2 => n6066, C1 => n3363, C2 => 
                           n6034, A => n3921, ZN => n3914);
   U4779 : OAI22_X1 port map( A1 => n5539, A2 => n3365, B1 => n5538, B2 => 
                           n3366, ZN => n3921);
   U4780 : INV_X1 port map( A => DATAIN(16), ZN => n2584);
   U4781 : OAI21_X1 port map( B1 => n3266, B2 => n1560, A => ENABLE, ZN => 
                           n7578);
   U4782 : OAI222_X1 port map( A1 => n2622, A2 => n3263, B1 => n3922, B2 => 
                           n3265, C1 => n3266, C2 => n1497, ZN => n7577);
   U4783 : NOR4_X1 port map( A1 => n3923, A2 => n3924, A3 => n3925, A4 => n3926
                           , ZN => n3922);
   U4784 : NAND4_X1 port map( A1 => n3927, A2 => n3928, A3 => n3929, A4 => 
                           n3930, ZN => n3926);
   U4785 : AOI221_X1 port map( B1 => n3275, B2 => n6417, C1 => n3276, C2 => 
                           n6449, A => n3931, ZN => n3930);
   U4786 : OAI222_X1 port map( A1 => n5265, A2 => n3278, B1 => n5233, B2 => 
                           n3279, C1 => n5201, C2 => n421, ZN => n3931);
   U4787 : AOI221_X1 port map( B1 => n3280, B2 => n761, C1 => n3281, C2 => n337
                           , A => n3932, ZN => n3929);
   U4788 : OAI22_X1 port map( A1 => n241, A2 => n413, B1 => n665, B2 => n3283, 
                           ZN => n3932);
   U4789 : AOI221_X1 port map( B1 => n3284, B2 => n6545, C1 => n3285, C2 => 
                           n6577, A => n3933, ZN => n3928);
   U4790 : OAI222_X1 port map( A1 => n5361, A2 => n3287, B1 => n5329, B2 => 
                           n1579, C1 => n5297, C2 => n3288, ZN => n3933);
   U4791 : AOI221_X1 port map( B1 => n3289, B2 => n762, C1 => n3290, C2 => n338
                           , A => n3934, ZN => n3927);
   U4792 : OAI22_X1 port map( A1 => n242, A2 => n414, B1 => n666, B2 => n3292, 
                           ZN => n3934);
   U4793 : NAND4_X1 port map( A1 => n3935, A2 => n3936, A3 => n3937, A4 => 
                           n3938, ZN => n3925);
   U4794 : AOI221_X1 port map( B1 => n3297, B2 => n6289, C1 => n3298, C2 => 
                           n6321, A => n3939, ZN => n3938);
   U4795 : OAI222_X1 port map( A1 => n5073, A2 => n3300, B1 => n5041, B2 => 
                           n3301, C1 => n5009, C2 => n3302, ZN => n3939);
   U4796 : AOI221_X1 port map( B1 => n3303, B2 => n537, C1 => n3304, C2 => n177
                           , A => n3940, ZN => n3937);
   U4797 : OAI22_X1 port map( A1 => n441, A2 => n3306, B1 => n81, B2 => n3307, 
                           ZN => n3940);
   U4798 : AOI221_X1 port map( B1 => n3308, B2 => n6353, C1 => n3309, C2 => 
                           n6385, A => n3941, ZN => n3936);
   U4799 : OAI222_X1 port map( A1 => n5169, A2 => n3311, B1 => n5137, B2 => 
                           n3312, C1 => n5105, C2 => n422, ZN => n3941);
   U4800 : AOI221_X1 port map( B1 => n3313, B2 => n585, C1 => n3314, C2 => n129
                           , A => n3942, ZN => n3935);
   U4801 : OAI22_X1 port map( A1 => n33, A2 => n415, B1 => n489, B2 => n3316, 
                           ZN => n3942);
   U4802 : NAND4_X1 port map( A1 => n3943, A2 => n3944, A3 => n3945, A4 => 
                           n3946, ZN => n3924);
   U4803 : AOI221_X1 port map( B1 => n3321, B2 => n6097, C1 => n3322, C2 => 
                           n6129, A => n3947, ZN => n3946);
   U4804 : OAI222_X1 port map( A1 => n4881, A2 => n3324, B1 => n4849, B2 => 
                           n3325, C1 => n4817, C2 => n423, ZN => n3947);
   U4805 : AOI221_X1 port map( B1 => n3326, B2 => n763, C1 => n3327, C2 => n339
                           , A => n3948, ZN => n3945);
   U4806 : OAI22_X1 port map( A1 => n243, A2 => n3329, B1 => n667, B2 => n3330,
                           ZN => n3948);
   U4807 : AOI221_X1 port map( B1 => n3331, B2 => n6225, C1 => n3332, C2 => 
                           n6257, A => n3949, ZN => n3944);
   U4808 : OAI222_X1 port map( A1 => n4977, A2 => n3334, B1 => n4945, B2 => 
                           n3335, C1 => n4913, C2 => n3336, ZN => n3949);
   U4809 : AOI221_X1 port map( B1 => n3337, B2 => n586, C1 => n3338, C2 => n130
                           , A => n3950, ZN => n3943);
   U4810 : OAI22_X1 port map( A1 => n34, A2 => n3340, B1 => n490, B2 => n3341, 
                           ZN => n3950);
   U4811 : NAND4_X1 port map( A1 => n3951, A2 => n3952, A3 => n3953, A4 => 
                           n3954, ZN => n3923);
   U4812 : AOI221_X1 port map( B1 => n3346, B2 => n5841, C1 => n3347, C2 => 
                           n5873, A => n3955, ZN => n3954);
   U4813 : OAI222_X1 port map( A1 => n4625, A2 => n3349, B1 => n4593, B2 => 
                           n3350, C1 => n4561, C2 => n3351, ZN => n3955);
   U4814 : AOI221_X1 port map( B1 => n3352, B2 => n5905, C1 => n3353, C2 => 
                           n5937, A => n3956, ZN => n3953);
   U4815 : OAI22_X1 port map( A1 => n4689, A2 => n3355, B1 => n4657, B2 => 
                           n3356, ZN => n3956);
   U4816 : AOI221_X1 port map( B1 => n3357, B2 => n5969, C1 => n3358, C2 => 
                           n6001, A => n3957, ZN => n3952);
   U4817 : OAI222_X1 port map( A1 => n4785, A2 => n3360, B1 => n4753, B2 => 
                           n3361, C1 => n4721, C2 => n424, ZN => n3957);
   U4818 : AOI221_X1 port map( B1 => n3362, B2 => n6065, C1 => n3363, C2 => 
                           n6033, A => n3958, ZN => n3951);
   U4819 : OAI22_X1 port map( A1 => n5529, A2 => n3365, B1 => n5528, B2 => 
                           n3366, ZN => n3958);
   U4820 : INV_X1 port map( A => DATAIN(15), ZN => n2622);
   U4821 : OAI21_X1 port map( B1 => n3266, B2 => n1561, A => ENABLE, ZN => 
                           n7576);
   U4822 : OAI222_X1 port map( A1 => n2660, A2 => n3263, B1 => n3959, B2 => 
                           n3265, C1 => n3266, C2 => n1498, ZN => n7575);
   U4823 : NOR4_X1 port map( A1 => n3960, A2 => n3961, A3 => n3962, A4 => n3963
                           , ZN => n3959);
   U4824 : NAND4_X1 port map( A1 => n3964, A2 => n3965, A3 => n3966, A4 => 
                           n3967, ZN => n3963);
   U4825 : AOI221_X1 port map( B1 => n3275, B2 => n6416, C1 => n3276, C2 => 
                           n6448, A => n3968, ZN => n3967);
   U4826 : OAI222_X1 port map( A1 => n5264, A2 => n3278, B1 => n5232, B2 => 
                           n3279, C1 => n5200, C2 => n421, ZN => n3968);
   U4827 : AOI221_X1 port map( B1 => n3280, B2 => n764, C1 => n3281, C2 => n340
                           , A => n3969, ZN => n3966);
   U4828 : OAI22_X1 port map( A1 => n244, A2 => n413, B1 => n668, B2 => n3283, 
                           ZN => n3969);
   U4829 : AOI221_X1 port map( B1 => n3284, B2 => n6544, C1 => n3285, C2 => 
                           n6576, A => n3970, ZN => n3965);
   U4830 : OAI222_X1 port map( A1 => n5360, A2 => n3287, B1 => n5328, B2 => 
                           n1579, C1 => n5296, C2 => n3288, ZN => n3970);
   U4831 : AOI221_X1 port map( B1 => n3289, B2 => n765, C1 => n3290, C2 => n341
                           , A => n3971, ZN => n3964);
   U4832 : OAI22_X1 port map( A1 => n245, A2 => n414, B1 => n669, B2 => n3292, 
                           ZN => n3971);
   U4833 : NAND4_X1 port map( A1 => n3972, A2 => n3973, A3 => n3974, A4 => 
                           n3975, ZN => n3962);
   U4834 : AOI221_X1 port map( B1 => n3297, B2 => n6288, C1 => n3298, C2 => 
                           n6320, A => n3976, ZN => n3975);
   U4835 : OAI222_X1 port map( A1 => n5072, A2 => n3300, B1 => n5040, B2 => 
                           n3301, C1 => n5008, C2 => n3302, ZN => n3976);
   U4836 : AOI221_X1 port map( B1 => n3303, B2 => n538, C1 => n3304, C2 => n178
                           , A => n3977, ZN => n3974);
   U4837 : OAI22_X1 port map( A1 => n442, A2 => n3306, B1 => n82, B2 => n3307, 
                           ZN => n3977);
   U4838 : AOI221_X1 port map( B1 => n3308, B2 => n6352, C1 => n3309, C2 => 
                           n6384, A => n3978, ZN => n3973);
   U4839 : OAI222_X1 port map( A1 => n5168, A2 => n3311, B1 => n5136, B2 => 
                           n3312, C1 => n5104, C2 => n422, ZN => n3978);
   U4840 : AOI221_X1 port map( B1 => n3313, B2 => n587, C1 => n3314, C2 => n131
                           , A => n3979, ZN => n3972);
   U4841 : OAI22_X1 port map( A1 => n35, A2 => n415, B1 => n491, B2 => n3316, 
                           ZN => n3979);
   U4842 : NAND4_X1 port map( A1 => n3980, A2 => n3981, A3 => n3982, A4 => 
                           n3983, ZN => n3961);
   U4843 : AOI221_X1 port map( B1 => n3321, B2 => n6096, C1 => n3322, C2 => 
                           n6128, A => n3984, ZN => n3983);
   U4844 : OAI222_X1 port map( A1 => n4880, A2 => n3324, B1 => n4848, B2 => 
                           n3325, C1 => n4816, C2 => n423, ZN => n3984);
   U4845 : AOI221_X1 port map( B1 => n3326, B2 => n766, C1 => n3327, C2 => n342
                           , A => n3985, ZN => n3982);
   U4846 : OAI22_X1 port map( A1 => n246, A2 => n3329, B1 => n670, B2 => n3330,
                           ZN => n3985);
   U4847 : AOI221_X1 port map( B1 => n3331, B2 => n6224, C1 => n3332, C2 => 
                           n6256, A => n3986, ZN => n3981);
   U4848 : OAI222_X1 port map( A1 => n4976, A2 => n3334, B1 => n4944, B2 => 
                           n3335, C1 => n4912, C2 => n3336, ZN => n3986);
   U4849 : AOI221_X1 port map( B1 => n3337, B2 => n588, C1 => n3338, C2 => n132
                           , A => n3987, ZN => n3980);
   U4850 : OAI22_X1 port map( A1 => n36, A2 => n3340, B1 => n492, B2 => n3341, 
                           ZN => n3987);
   U4851 : NAND4_X1 port map( A1 => n3988, A2 => n3989, A3 => n3990, A4 => 
                           n3991, ZN => n3960);
   U4852 : AOI221_X1 port map( B1 => n3346, B2 => n5840, C1 => n3347, C2 => 
                           n5872, A => n3992, ZN => n3991);
   U4853 : OAI222_X1 port map( A1 => n4624, A2 => n3349, B1 => n4592, B2 => 
                           n3350, C1 => n4560, C2 => n3351, ZN => n3992);
   U4854 : AOI221_X1 port map( B1 => n3352, B2 => n5904, C1 => n3353, C2 => 
                           n5936, A => n3993, ZN => n3990);
   U4855 : OAI22_X1 port map( A1 => n4688, A2 => n3355, B1 => n4656, B2 => 
                           n3356, ZN => n3993);
   U4856 : AOI221_X1 port map( B1 => n3357, B2 => n5968, C1 => n3358, C2 => 
                           n6000, A => n3994, ZN => n3989);
   U4857 : OAI222_X1 port map( A1 => n4784, A2 => n3360, B1 => n4752, B2 => 
                           n3361, C1 => n4720, C2 => n424, ZN => n3994);
   U4858 : AOI221_X1 port map( B1 => n3362, B2 => n6064, C1 => n3363, C2 => 
                           n6032, A => n3995, ZN => n3988);
   U4859 : OAI22_X1 port map( A1 => n5519, A2 => n3365, B1 => n5518, B2 => 
                           n3366, ZN => n3995);
   U4860 : INV_X1 port map( A => DATAIN(14), ZN => n2660);
   U4861 : OAI21_X1 port map( B1 => n3266, B2 => n1562, A => ENABLE, ZN => 
                           n7574);
   U4862 : OAI222_X1 port map( A1 => n2698, A2 => n3263, B1 => n3996, B2 => 
                           n3265, C1 => n3266, C2 => n1499, ZN => n7573);
   U4863 : NOR4_X1 port map( A1 => n3997, A2 => n3998, A3 => n3999, A4 => n4000
                           , ZN => n3996);
   U4864 : NAND4_X1 port map( A1 => n4001, A2 => n4002, A3 => n4003, A4 => 
                           n4004, ZN => n4000);
   U4865 : AOI221_X1 port map( B1 => n3275, B2 => n6415, C1 => n3276, C2 => 
                           n6447, A => n4005, ZN => n4004);
   U4866 : OAI222_X1 port map( A1 => n5263, A2 => n3278, B1 => n5231, B2 => 
                           n3279, C1 => n5199, C2 => n421, ZN => n4005);
   U4867 : AOI221_X1 port map( B1 => n3280, B2 => n767, C1 => n3281, C2 => n343
                           , A => n4006, ZN => n4003);
   U4868 : OAI22_X1 port map( A1 => n247, A2 => n413, B1 => n671, B2 => n3283, 
                           ZN => n4006);
   U4869 : AOI221_X1 port map( B1 => n3284, B2 => n6543, C1 => n3285, C2 => 
                           n6575, A => n4007, ZN => n4002);
   U4870 : OAI222_X1 port map( A1 => n5359, A2 => n3287, B1 => n5327, B2 => 
                           n1579, C1 => n5295, C2 => n3288, ZN => n4007);
   U4871 : AOI221_X1 port map( B1 => n3289, B2 => n768, C1 => n3290, C2 => n344
                           , A => n4008, ZN => n4001);
   U4872 : OAI22_X1 port map( A1 => n248, A2 => n414, B1 => n672, B2 => n3292, 
                           ZN => n4008);
   U4873 : NAND4_X1 port map( A1 => n4009, A2 => n4010, A3 => n4011, A4 => 
                           n4012, ZN => n3999);
   U4874 : AOI221_X1 port map( B1 => n3297, B2 => n6287, C1 => n3298, C2 => 
                           n6319, A => n4013, ZN => n4012);
   U4875 : OAI222_X1 port map( A1 => n5071, A2 => n3300, B1 => n5039, B2 => 
                           n3301, C1 => n5007, C2 => n3302, ZN => n4013);
   U4876 : AOI221_X1 port map( B1 => n3303, B2 => n539, C1 => n3304, C2 => n179
                           , A => n4014, ZN => n4011);
   U4877 : OAI22_X1 port map( A1 => n443, A2 => n3306, B1 => n83, B2 => n3307, 
                           ZN => n4014);
   U4878 : AOI221_X1 port map( B1 => n3308, B2 => n6351, C1 => n3309, C2 => 
                           n6383, A => n4015, ZN => n4010);
   U4879 : OAI222_X1 port map( A1 => n5167, A2 => n3311, B1 => n5135, B2 => 
                           n3312, C1 => n5103, C2 => n422, ZN => n4015);
   U4880 : AOI221_X1 port map( B1 => n3313, B2 => n589, C1 => n3314, C2 => n133
                           , A => n4016, ZN => n4009);
   U4881 : OAI22_X1 port map( A1 => n37, A2 => n415, B1 => n493, B2 => n3316, 
                           ZN => n4016);
   U4882 : NAND4_X1 port map( A1 => n4017, A2 => n4018, A3 => n4019, A4 => 
                           n4020, ZN => n3998);
   U4883 : AOI221_X1 port map( B1 => n3321, B2 => n6095, C1 => n3322, C2 => 
                           n6127, A => n4021, ZN => n4020);
   U4884 : OAI222_X1 port map( A1 => n4879, A2 => n3324, B1 => n4847, B2 => 
                           n3325, C1 => n4815, C2 => n423, ZN => n4021);
   U4885 : AOI221_X1 port map( B1 => n3326, B2 => n769, C1 => n3327, C2 => n345
                           , A => n4022, ZN => n4019);
   U4886 : OAI22_X1 port map( A1 => n249, A2 => n3329, B1 => n673, B2 => n3330,
                           ZN => n4022);
   U4887 : AOI221_X1 port map( B1 => n3331, B2 => n6223, C1 => n3332, C2 => 
                           n6255, A => n4023, ZN => n4018);
   U4888 : OAI222_X1 port map( A1 => n4975, A2 => n3334, B1 => n4943, B2 => 
                           n3335, C1 => n4911, C2 => n3336, ZN => n4023);
   U4889 : AOI221_X1 port map( B1 => n3337, B2 => n590, C1 => n3338, C2 => n134
                           , A => n4024, ZN => n4017);
   U4890 : OAI22_X1 port map( A1 => n38, A2 => n3340, B1 => n494, B2 => n3341, 
                           ZN => n4024);
   U4891 : NAND4_X1 port map( A1 => n4025, A2 => n4026, A3 => n4027, A4 => 
                           n4028, ZN => n3997);
   U4892 : AOI221_X1 port map( B1 => n3346, B2 => n5839, C1 => n3347, C2 => 
                           n5871, A => n4029, ZN => n4028);
   U4893 : OAI222_X1 port map( A1 => n4623, A2 => n3349, B1 => n4591, B2 => 
                           n3350, C1 => n4559, C2 => n3351, ZN => n4029);
   U4894 : AOI221_X1 port map( B1 => n3352, B2 => n5903, C1 => n3353, C2 => 
                           n5935, A => n4030, ZN => n4027);
   U4895 : OAI22_X1 port map( A1 => n4687, A2 => n3355, B1 => n4655, B2 => 
                           n3356, ZN => n4030);
   U4896 : AOI221_X1 port map( B1 => n3357, B2 => n5967, C1 => n3358, C2 => 
                           n5999, A => n4031, ZN => n4026);
   U4897 : OAI222_X1 port map( A1 => n4783, A2 => n3360, B1 => n4751, B2 => 
                           n3361, C1 => n4719, C2 => n424, ZN => n4031);
   U4898 : AOI221_X1 port map( B1 => n3362, B2 => n6063, C1 => n3363, C2 => 
                           n6031, A => n4032, ZN => n4025);
   U4899 : OAI22_X1 port map( A1 => n5509, A2 => n3365, B1 => n5508, B2 => 
                           n3366, ZN => n4032);
   U4900 : INV_X1 port map( A => DATAIN(13), ZN => n2698);
   U4901 : OAI21_X1 port map( B1 => n3266, B2 => n1563, A => ENABLE, ZN => 
                           n7572);
   U4902 : OAI222_X1 port map( A1 => n2736, A2 => n3263, B1 => n4033, B2 => 
                           n3265, C1 => n3266, C2 => n1500, ZN => n7571);
   U4903 : NOR4_X1 port map( A1 => n4034, A2 => n4035, A3 => n4036, A4 => n4037
                           , ZN => n4033);
   U4904 : NAND4_X1 port map( A1 => n4038, A2 => n4039, A3 => n4040, A4 => 
                           n4041, ZN => n4037);
   U4905 : AOI221_X1 port map( B1 => n3275, B2 => n6414, C1 => n3276, C2 => 
                           n6446, A => n4042, ZN => n4041);
   U4906 : OAI222_X1 port map( A1 => n5262, A2 => n3278, B1 => n5230, B2 => 
                           n3279, C1 => n5198, C2 => n421, ZN => n4042);
   U4907 : AOI221_X1 port map( B1 => n3280, B2 => n770, C1 => n3281, C2 => n346
                           , A => n4043, ZN => n4040);
   U4908 : OAI22_X1 port map( A1 => n250, A2 => n413, B1 => n674, B2 => n3283, 
                           ZN => n4043);
   U4909 : AOI221_X1 port map( B1 => n3284, B2 => n6542, C1 => n3285, C2 => 
                           n6574, A => n4044, ZN => n4039);
   U4910 : OAI222_X1 port map( A1 => n5358, A2 => n3287, B1 => n5326, B2 => 
                           n1579, C1 => n5294, C2 => n3288, ZN => n4044);
   U4911 : AOI221_X1 port map( B1 => n3289, B2 => n771, C1 => n3290, C2 => n347
                           , A => n4045, ZN => n4038);
   U4912 : OAI22_X1 port map( A1 => n251, A2 => n414, B1 => n675, B2 => n3292, 
                           ZN => n4045);
   U4913 : NAND4_X1 port map( A1 => n4046, A2 => n4047, A3 => n4048, A4 => 
                           n4049, ZN => n4036);
   U4914 : AOI221_X1 port map( B1 => n3297, B2 => n6286, C1 => n3298, C2 => 
                           n6318, A => n4050, ZN => n4049);
   U4915 : OAI222_X1 port map( A1 => n5070, A2 => n3300, B1 => n5038, B2 => 
                           n3301, C1 => n5006, C2 => n3302, ZN => n4050);
   U4916 : AOI221_X1 port map( B1 => n3303, B2 => n540, C1 => n3304, C2 => n180
                           , A => n4051, ZN => n4048);
   U4917 : OAI22_X1 port map( A1 => n444, A2 => n3306, B1 => n84, B2 => n3307, 
                           ZN => n4051);
   U4918 : AOI221_X1 port map( B1 => n3308, B2 => n6350, C1 => n3309, C2 => 
                           n6382, A => n4052, ZN => n4047);
   U4919 : OAI222_X1 port map( A1 => n5166, A2 => n3311, B1 => n5134, B2 => 
                           n3312, C1 => n5102, C2 => n422, ZN => n4052);
   U4920 : AOI221_X1 port map( B1 => n3313, B2 => n591, C1 => n3314, C2 => n135
                           , A => n4053, ZN => n4046);
   U4921 : OAI22_X1 port map( A1 => n39, A2 => n415, B1 => n495, B2 => n3316, 
                           ZN => n4053);
   U4922 : NAND4_X1 port map( A1 => n4054, A2 => n4055, A3 => n4056, A4 => 
                           n4057, ZN => n4035);
   U4923 : AOI221_X1 port map( B1 => n3321, B2 => n6094, C1 => n3322, C2 => 
                           n6126, A => n4058, ZN => n4057);
   U4924 : OAI222_X1 port map( A1 => n4878, A2 => n3324, B1 => n4846, B2 => 
                           n3325, C1 => n4814, C2 => n423, ZN => n4058);
   U4925 : AOI221_X1 port map( B1 => n3326, B2 => n772, C1 => n3327, C2 => n348
                           , A => n4059, ZN => n4056);
   U4926 : OAI22_X1 port map( A1 => n252, A2 => n3329, B1 => n676, B2 => n3330,
                           ZN => n4059);
   U4927 : AOI221_X1 port map( B1 => n3331, B2 => n6222, C1 => n3332, C2 => 
                           n6254, A => n4060, ZN => n4055);
   U4928 : OAI222_X1 port map( A1 => n4974, A2 => n3334, B1 => n4942, B2 => 
                           n3335, C1 => n4910, C2 => n3336, ZN => n4060);
   U4929 : AOI221_X1 port map( B1 => n3337, B2 => n592, C1 => n3338, C2 => n136
                           , A => n4061, ZN => n4054);
   U4930 : OAI22_X1 port map( A1 => n40, A2 => n3340, B1 => n496, B2 => n3341, 
                           ZN => n4061);
   U4931 : NAND4_X1 port map( A1 => n4062, A2 => n4063, A3 => n4064, A4 => 
                           n4065, ZN => n4034);
   U4932 : AOI221_X1 port map( B1 => n3346, B2 => n5838, C1 => n3347, C2 => 
                           n5870, A => n4066, ZN => n4065);
   U4933 : OAI222_X1 port map( A1 => n4622, A2 => n3349, B1 => n4590, B2 => 
                           n3350, C1 => n4558, C2 => n3351, ZN => n4066);
   U4934 : AOI221_X1 port map( B1 => n3352, B2 => n5902, C1 => n3353, C2 => 
                           n5934, A => n4067, ZN => n4064);
   U4935 : OAI22_X1 port map( A1 => n4686, A2 => n3355, B1 => n4654, B2 => 
                           n3356, ZN => n4067);
   U4936 : AOI221_X1 port map( B1 => n3357, B2 => n5966, C1 => n3358, C2 => 
                           n5998, A => n4068, ZN => n4063);
   U4937 : OAI222_X1 port map( A1 => n4782, A2 => n3360, B1 => n4750, B2 => 
                           n3361, C1 => n4718, C2 => n424, ZN => n4068);
   U4938 : AOI221_X1 port map( B1 => n3362, B2 => n6062, C1 => n3363, C2 => 
                           n6030, A => n4069, ZN => n4062);
   U4939 : OAI22_X1 port map( A1 => n5499, A2 => n3365, B1 => n5498, B2 => 
                           n3366, ZN => n4069);
   U4940 : INV_X1 port map( A => DATAIN(12), ZN => n2736);
   U4941 : OAI21_X1 port map( B1 => n3266, B2 => n1564, A => ENABLE, ZN => 
                           n7570);
   U4942 : OAI222_X1 port map( A1 => n2774, A2 => n3263, B1 => n4070, B2 => 
                           n3265, C1 => n3266, C2 => n1501, ZN => n7569);
   U4943 : NOR4_X1 port map( A1 => n4071, A2 => n4072, A3 => n4073, A4 => n4074
                           , ZN => n4070);
   U4944 : NAND4_X1 port map( A1 => n4075, A2 => n4076, A3 => n4077, A4 => 
                           n4078, ZN => n4074);
   U4945 : AOI221_X1 port map( B1 => n3275, B2 => n6413, C1 => n3276, C2 => 
                           n6445, A => n4079, ZN => n4078);
   U4946 : OAI222_X1 port map( A1 => n5261, A2 => n3278, B1 => n5229, B2 => 
                           n3279, C1 => n5197, C2 => n421, ZN => n4079);
   U4947 : AOI221_X1 port map( B1 => n3280, B2 => n773, C1 => n3281, C2 => n349
                           , A => n4080, ZN => n4077);
   U4948 : OAI22_X1 port map( A1 => n253, A2 => n413, B1 => n677, B2 => n3283, 
                           ZN => n4080);
   U4949 : AOI221_X1 port map( B1 => n3284, B2 => n6541, C1 => n3285, C2 => 
                           n6573, A => n4081, ZN => n4076);
   U4950 : OAI222_X1 port map( A1 => n5357, A2 => n3287, B1 => n5325, B2 => 
                           n1579, C1 => n5293, C2 => n3288, ZN => n4081);
   U4951 : AOI221_X1 port map( B1 => n3289, B2 => n774, C1 => n3290, C2 => n350
                           , A => n4082, ZN => n4075);
   U4952 : OAI22_X1 port map( A1 => n254, A2 => n414, B1 => n678, B2 => n3292, 
                           ZN => n4082);
   U4953 : NAND4_X1 port map( A1 => n4083, A2 => n4084, A3 => n4085, A4 => 
                           n4086, ZN => n4073);
   U4954 : AOI221_X1 port map( B1 => n3297, B2 => n6285, C1 => n3298, C2 => 
                           n6317, A => n4087, ZN => n4086);
   U4955 : OAI222_X1 port map( A1 => n5069, A2 => n3300, B1 => n5037, B2 => 
                           n3301, C1 => n5005, C2 => n3302, ZN => n4087);
   U4956 : AOI221_X1 port map( B1 => n3303, B2 => n541, C1 => n3304, C2 => n181
                           , A => n4088, ZN => n4085);
   U4957 : OAI22_X1 port map( A1 => n445, A2 => n3306, B1 => n85, B2 => n3307, 
                           ZN => n4088);
   U4958 : AOI221_X1 port map( B1 => n3308, B2 => n6349, C1 => n3309, C2 => 
                           n6381, A => n4089, ZN => n4084);
   U4959 : OAI222_X1 port map( A1 => n5165, A2 => n3311, B1 => n5133, B2 => 
                           n3312, C1 => n5101, C2 => n422, ZN => n4089);
   U4960 : AOI221_X1 port map( B1 => n3313, B2 => n593, C1 => n3314, C2 => n137
                           , A => n4090, ZN => n4083);
   U4961 : OAI22_X1 port map( A1 => n41, A2 => n415, B1 => n497, B2 => n3316, 
                           ZN => n4090);
   U4962 : NAND4_X1 port map( A1 => n4091, A2 => n4092, A3 => n4093, A4 => 
                           n4094, ZN => n4072);
   U4963 : AOI221_X1 port map( B1 => n3321, B2 => n6093, C1 => n3322, C2 => 
                           n6125, A => n4095, ZN => n4094);
   U4964 : OAI222_X1 port map( A1 => n4877, A2 => n3324, B1 => n4845, B2 => 
                           n3325, C1 => n4813, C2 => n423, ZN => n4095);
   U4965 : AOI221_X1 port map( B1 => n3326, B2 => n775, C1 => n3327, C2 => n351
                           , A => n4096, ZN => n4093);
   U4966 : OAI22_X1 port map( A1 => n255, A2 => n3329, B1 => n679, B2 => n3330,
                           ZN => n4096);
   U4967 : AOI221_X1 port map( B1 => n3331, B2 => n6221, C1 => n3332, C2 => 
                           n6253, A => n4097, ZN => n4092);
   U4968 : OAI222_X1 port map( A1 => n4973, A2 => n3334, B1 => n4941, B2 => 
                           n3335, C1 => n4909, C2 => n3336, ZN => n4097);
   U4969 : AOI221_X1 port map( B1 => n3337, B2 => n594, C1 => n3338, C2 => n138
                           , A => n4098, ZN => n4091);
   U4970 : OAI22_X1 port map( A1 => n42, A2 => n3340, B1 => n498, B2 => n3341, 
                           ZN => n4098);
   U4971 : NAND4_X1 port map( A1 => n4099, A2 => n4100, A3 => n4101, A4 => 
                           n4102, ZN => n4071);
   U4972 : AOI221_X1 port map( B1 => n3346, B2 => n5837, C1 => n3347, C2 => 
                           n5869, A => n4103, ZN => n4102);
   U4973 : OAI222_X1 port map( A1 => n4621, A2 => n3349, B1 => n4589, B2 => 
                           n3350, C1 => n4557, C2 => n3351, ZN => n4103);
   U4974 : AOI221_X1 port map( B1 => n3352, B2 => n5901, C1 => n3353, C2 => 
                           n5933, A => n4104, ZN => n4101);
   U4975 : OAI22_X1 port map( A1 => n4685, A2 => n3355, B1 => n4653, B2 => 
                           n3356, ZN => n4104);
   U4976 : AOI221_X1 port map( B1 => n3357, B2 => n5965, C1 => n3358, C2 => 
                           n5997, A => n4105, ZN => n4100);
   U4977 : OAI222_X1 port map( A1 => n4781, A2 => n3360, B1 => n4749, B2 => 
                           n3361, C1 => n4717, C2 => n424, ZN => n4105);
   U4978 : AOI221_X1 port map( B1 => n3362, B2 => n6061, C1 => n3363, C2 => 
                           n6029, A => n4106, ZN => n4099);
   U4979 : OAI22_X1 port map( A1 => n5489, A2 => n3365, B1 => n5488, B2 => 
                           n3366, ZN => n4106);
   U4980 : INV_X1 port map( A => DATAIN(11), ZN => n2774);
   U4981 : OAI21_X1 port map( B1 => n3266, B2 => n1565, A => ENABLE, ZN => 
                           n7568);
   U4982 : OAI222_X1 port map( A1 => n2812, A2 => n3263, B1 => n4107, B2 => 
                           n3265, C1 => n3266, C2 => n1502, ZN => n7567);
   U4983 : NOR4_X1 port map( A1 => n4108, A2 => n4109, A3 => n4110, A4 => n4111
                           , ZN => n4107);
   U4984 : NAND4_X1 port map( A1 => n4112, A2 => n4113, A3 => n4114, A4 => 
                           n4115, ZN => n4111);
   U4985 : AOI221_X1 port map( B1 => n3275, B2 => n6412, C1 => n3276, C2 => 
                           n6444, A => n4116, ZN => n4115);
   U4986 : OAI222_X1 port map( A1 => n5260, A2 => n3278, B1 => n5228, B2 => 
                           n3279, C1 => n5196, C2 => n421, ZN => n4116);
   U4987 : AOI221_X1 port map( B1 => n3280, B2 => n776, C1 => n3281, C2 => n352
                           , A => n4117, ZN => n4114);
   U4988 : OAI22_X1 port map( A1 => n256, A2 => n413, B1 => n680, B2 => n3283, 
                           ZN => n4117);
   U4989 : AOI221_X1 port map( B1 => n3284, B2 => n6540, C1 => n3285, C2 => 
                           n6572, A => n4118, ZN => n4113);
   U4990 : OAI222_X1 port map( A1 => n5356, A2 => n3287, B1 => n5324, B2 => 
                           n1579, C1 => n5292, C2 => n3288, ZN => n4118);
   U4991 : AOI221_X1 port map( B1 => n3289, B2 => n777, C1 => n3290, C2 => n353
                           , A => n4119, ZN => n4112);
   U4992 : OAI22_X1 port map( A1 => n257, A2 => n414, B1 => n681, B2 => n3292, 
                           ZN => n4119);
   U4993 : NAND4_X1 port map( A1 => n4120, A2 => n4121, A3 => n4122, A4 => 
                           n4123, ZN => n4110);
   U4994 : AOI221_X1 port map( B1 => n3297, B2 => n6284, C1 => n3298, C2 => 
                           n6316, A => n4124, ZN => n4123);
   U4995 : OAI222_X1 port map( A1 => n5068, A2 => n3300, B1 => n5036, B2 => 
                           n3301, C1 => n5004, C2 => n3302, ZN => n4124);
   U4996 : AOI221_X1 port map( B1 => n3303, B2 => n542, C1 => n3304, C2 => n182
                           , A => n4125, ZN => n4122);
   U4997 : OAI22_X1 port map( A1 => n446, A2 => n3306, B1 => n86, B2 => n3307, 
                           ZN => n4125);
   U4998 : AOI221_X1 port map( B1 => n3308, B2 => n6348, C1 => n3309, C2 => 
                           n6380, A => n4126, ZN => n4121);
   U4999 : OAI222_X1 port map( A1 => n5164, A2 => n3311, B1 => n5132, B2 => 
                           n3312, C1 => n5100, C2 => n422, ZN => n4126);
   U5000 : AOI221_X1 port map( B1 => n3313, B2 => n595, C1 => n3314, C2 => n139
                           , A => n4127, ZN => n4120);
   U5001 : OAI22_X1 port map( A1 => n43, A2 => n415, B1 => n499, B2 => n3316, 
                           ZN => n4127);
   U5002 : NAND4_X1 port map( A1 => n4128, A2 => n4129, A3 => n4130, A4 => 
                           n4131, ZN => n4109);
   U5003 : AOI221_X1 port map( B1 => n3321, B2 => n6092, C1 => n3322, C2 => 
                           n6124, A => n4132, ZN => n4131);
   U5004 : OAI222_X1 port map( A1 => n4876, A2 => n3324, B1 => n4844, B2 => 
                           n3325, C1 => n4812, C2 => n423, ZN => n4132);
   U5005 : AOI221_X1 port map( B1 => n3326, B2 => n778, C1 => n3327, C2 => n354
                           , A => n4133, ZN => n4130);
   U5006 : OAI22_X1 port map( A1 => n258, A2 => n3329, B1 => n682, B2 => n3330,
                           ZN => n4133);
   U5007 : AOI221_X1 port map( B1 => n3331, B2 => n6220, C1 => n3332, C2 => 
                           n6252, A => n4134, ZN => n4129);
   U5008 : OAI222_X1 port map( A1 => n4972, A2 => n3334, B1 => n4940, B2 => 
                           n3335, C1 => n4908, C2 => n3336, ZN => n4134);
   U5009 : AOI221_X1 port map( B1 => n3337, B2 => n596, C1 => n3338, C2 => n140
                           , A => n4135, ZN => n4128);
   U5010 : OAI22_X1 port map( A1 => n44, A2 => n3340, B1 => n500, B2 => n3341, 
                           ZN => n4135);
   U5011 : NAND4_X1 port map( A1 => n4136, A2 => n4137, A3 => n4138, A4 => 
                           n4139, ZN => n4108);
   U5012 : AOI221_X1 port map( B1 => n3346, B2 => n5836, C1 => n3347, C2 => 
                           n5868, A => n4140, ZN => n4139);
   U5013 : OAI222_X1 port map( A1 => n4620, A2 => n3349, B1 => n4588, B2 => 
                           n3350, C1 => n4556, C2 => n3351, ZN => n4140);
   U5014 : AOI221_X1 port map( B1 => n3352, B2 => n5900, C1 => n3353, C2 => 
                           n5932, A => n4141, ZN => n4138);
   U5015 : OAI22_X1 port map( A1 => n4684, A2 => n3355, B1 => n4652, B2 => 
                           n3356, ZN => n4141);
   U5016 : AOI221_X1 port map( B1 => n3357, B2 => n5964, C1 => n3358, C2 => 
                           n5996, A => n4142, ZN => n4137);
   U5017 : OAI222_X1 port map( A1 => n4780, A2 => n3360, B1 => n4748, B2 => 
                           n3361, C1 => n4716, C2 => n424, ZN => n4142);
   U5018 : AOI221_X1 port map( B1 => n3362, B2 => n6060, C1 => n3363, C2 => 
                           n6028, A => n4143, ZN => n4136);
   U5019 : OAI22_X1 port map( A1 => n5479, A2 => n3365, B1 => n5478, B2 => 
                           n3366, ZN => n4143);
   U5020 : INV_X1 port map( A => DATAIN(10), ZN => n2812);
   U5021 : OAI21_X1 port map( B1 => n3266, B2 => n1566, A => ENABLE, ZN => 
                           n7566);
   U5022 : OAI222_X1 port map( A1 => n2850, A2 => n3263, B1 => n4144, B2 => 
                           n3265, C1 => n3266, C2 => n1503, ZN => n7565);
   U5023 : NOR4_X1 port map( A1 => n4145, A2 => n4146, A3 => n4147, A4 => n4148
                           , ZN => n4144);
   U5024 : NAND4_X1 port map( A1 => n4149, A2 => n4150, A3 => n4151, A4 => 
                           n4152, ZN => n4148);
   U5025 : AOI221_X1 port map( B1 => n3275, B2 => n6411, C1 => n3276, C2 => 
                           n6443, A => n4153, ZN => n4152);
   U5026 : OAI222_X1 port map( A1 => n5259, A2 => n3278, B1 => n5227, B2 => 
                           n3279, C1 => n5195, C2 => n421, ZN => n4153);
   U5027 : AOI221_X1 port map( B1 => n3280, B2 => n779, C1 => n3281, C2 => n355
                           , A => n4154, ZN => n4151);
   U5028 : OAI22_X1 port map( A1 => n259, A2 => n413, B1 => n683, B2 => n3283, 
                           ZN => n4154);
   U5029 : AOI221_X1 port map( B1 => n3284, B2 => n6539, C1 => n3285, C2 => 
                           n6571, A => n4155, ZN => n4150);
   U5030 : OAI222_X1 port map( A1 => n5355, A2 => n3287, B1 => n5323, B2 => 
                           n1579, C1 => n5291, C2 => n3288, ZN => n4155);
   U5031 : AOI221_X1 port map( B1 => n3289, B2 => n780, C1 => n3290, C2 => n356
                           , A => n4156, ZN => n4149);
   U5032 : OAI22_X1 port map( A1 => n260, A2 => n414, B1 => n684, B2 => n3292, 
                           ZN => n4156);
   U5033 : NAND4_X1 port map( A1 => n4157, A2 => n4158, A3 => n4159, A4 => 
                           n4160, ZN => n4147);
   U5034 : AOI221_X1 port map( B1 => n3297, B2 => n6283, C1 => n3298, C2 => 
                           n6315, A => n4161, ZN => n4160);
   U5035 : OAI222_X1 port map( A1 => n5067, A2 => n3300, B1 => n5035, B2 => 
                           n3301, C1 => n5003, C2 => n3302, ZN => n4161);
   U5036 : AOI221_X1 port map( B1 => n3303, B2 => n543, C1 => n3304, C2 => n183
                           , A => n4162, ZN => n4159);
   U5037 : OAI22_X1 port map( A1 => n447, A2 => n3306, B1 => n87, B2 => n3307, 
                           ZN => n4162);
   U5038 : AOI221_X1 port map( B1 => n3308, B2 => n6347, C1 => n3309, C2 => 
                           n6379, A => n4163, ZN => n4158);
   U5039 : OAI222_X1 port map( A1 => n5163, A2 => n3311, B1 => n5131, B2 => 
                           n3312, C1 => n5099, C2 => n422, ZN => n4163);
   U5040 : AOI221_X1 port map( B1 => n3313, B2 => n597, C1 => n3314, C2 => n141
                           , A => n4164, ZN => n4157);
   U5041 : OAI22_X1 port map( A1 => n45, A2 => n415, B1 => n501, B2 => n3316, 
                           ZN => n4164);
   U5042 : NAND4_X1 port map( A1 => n4165, A2 => n4166, A3 => n4167, A4 => 
                           n4168, ZN => n4146);
   U5043 : AOI221_X1 port map( B1 => n3321, B2 => n6091, C1 => n3322, C2 => 
                           n6123, A => n4169, ZN => n4168);
   U5044 : OAI222_X1 port map( A1 => n4875, A2 => n3324, B1 => n4843, B2 => 
                           n3325, C1 => n4811, C2 => n423, ZN => n4169);
   U5045 : AOI221_X1 port map( B1 => n3326, B2 => n781, C1 => n3327, C2 => n357
                           , A => n4170, ZN => n4167);
   U5046 : OAI22_X1 port map( A1 => n261, A2 => n3329, B1 => n685, B2 => n3330,
                           ZN => n4170);
   U5047 : AOI221_X1 port map( B1 => n3331, B2 => n6219, C1 => n3332, C2 => 
                           n6251, A => n4171, ZN => n4166);
   U5048 : OAI222_X1 port map( A1 => n4971, A2 => n3334, B1 => n4939, B2 => 
                           n3335, C1 => n4907, C2 => n3336, ZN => n4171);
   U5049 : AOI221_X1 port map( B1 => n3337, B2 => n598, C1 => n3338, C2 => n142
                           , A => n4172, ZN => n4165);
   U5050 : OAI22_X1 port map( A1 => n46, A2 => n3340, B1 => n502, B2 => n3341, 
                           ZN => n4172);
   U5051 : NAND4_X1 port map( A1 => n4173, A2 => n4174, A3 => n4175, A4 => 
                           n4176, ZN => n4145);
   U5052 : AOI221_X1 port map( B1 => n3346, B2 => n5835, C1 => n3347, C2 => 
                           n5867, A => n4177, ZN => n4176);
   U5053 : OAI222_X1 port map( A1 => n4619, A2 => n3349, B1 => n4587, B2 => 
                           n3350, C1 => n4555, C2 => n3351, ZN => n4177);
   U5054 : AOI221_X1 port map( B1 => n3352, B2 => n5899, C1 => n3353, C2 => 
                           n5931, A => n4178, ZN => n4175);
   U5055 : OAI22_X1 port map( A1 => n4683, A2 => n3355, B1 => n4651, B2 => 
                           n3356, ZN => n4178);
   U5056 : AOI221_X1 port map( B1 => n3357, B2 => n5963, C1 => n3358, C2 => 
                           n5995, A => n4179, ZN => n4174);
   U5057 : OAI222_X1 port map( A1 => n4779, A2 => n3360, B1 => n4747, B2 => 
                           n3361, C1 => n4715, C2 => n424, ZN => n4179);
   U5058 : AOI221_X1 port map( B1 => n3362, B2 => n6059, C1 => n3363, C2 => 
                           n6027, A => n4180, ZN => n4173);
   U5059 : OAI22_X1 port map( A1 => n5469, A2 => n3365, B1 => n5468, B2 => 
                           n3366, ZN => n4180);
   U5060 : INV_X1 port map( A => DATAIN(9), ZN => n2850);
   U5061 : OAI21_X1 port map( B1 => n3266, B2 => n1567, A => ENABLE, ZN => 
                           n7564);
   U5062 : OAI222_X1 port map( A1 => n2888, A2 => n3263, B1 => n4181, B2 => 
                           n3265, C1 => n3266, C2 => n1504, ZN => n7563);
   U5063 : NOR4_X1 port map( A1 => n4182, A2 => n4183, A3 => n4184, A4 => n4185
                           , ZN => n4181);
   U5064 : NAND4_X1 port map( A1 => n4186, A2 => n4187, A3 => n4188, A4 => 
                           n4189, ZN => n4185);
   U5065 : AOI221_X1 port map( B1 => n3275, B2 => n6410, C1 => n3276, C2 => 
                           n6442, A => n4190, ZN => n4189);
   U5066 : OAI222_X1 port map( A1 => n5258, A2 => n3278, B1 => n5226, B2 => 
                           n3279, C1 => n5194, C2 => n421, ZN => n4190);
   U5067 : AOI221_X1 port map( B1 => n3280, B2 => n782, C1 => n3281, C2 => n358
                           , A => n4191, ZN => n4188);
   U5068 : OAI22_X1 port map( A1 => n262, A2 => n413, B1 => n686, B2 => n3283, 
                           ZN => n4191);
   U5069 : AOI221_X1 port map( B1 => n3284, B2 => n6538, C1 => n3285, C2 => 
                           n6570, A => n4192, ZN => n4187);
   U5070 : OAI222_X1 port map( A1 => n5354, A2 => n3287, B1 => n5322, B2 => 
                           n1579, C1 => n5290, C2 => n3288, ZN => n4192);
   U5071 : AOI221_X1 port map( B1 => n3289, B2 => n783, C1 => n3290, C2 => n359
                           , A => n4193, ZN => n4186);
   U5072 : OAI22_X1 port map( A1 => n263, A2 => n414, B1 => n687, B2 => n3292, 
                           ZN => n4193);
   U5073 : NAND4_X1 port map( A1 => n4194, A2 => n4195, A3 => n4196, A4 => 
                           n4197, ZN => n4184);
   U5074 : AOI221_X1 port map( B1 => n3297, B2 => n6282, C1 => n3298, C2 => 
                           n6314, A => n4198, ZN => n4197);
   U5075 : OAI222_X1 port map( A1 => n5066, A2 => n3300, B1 => n5034, B2 => 
                           n3301, C1 => n5002, C2 => n3302, ZN => n4198);
   U5076 : AOI221_X1 port map( B1 => n3303, B2 => n544, C1 => n3304, C2 => n184
                           , A => n4199, ZN => n4196);
   U5077 : OAI22_X1 port map( A1 => n448, A2 => n3306, B1 => n88, B2 => n3307, 
                           ZN => n4199);
   U5078 : AOI221_X1 port map( B1 => n3308, B2 => n6346, C1 => n3309, C2 => 
                           n6378, A => n4200, ZN => n4195);
   U5079 : OAI222_X1 port map( A1 => n5162, A2 => n3311, B1 => n5130, B2 => 
                           n3312, C1 => n5098, C2 => n422, ZN => n4200);
   U5080 : AOI221_X1 port map( B1 => n3313, B2 => n599, C1 => n3314, C2 => n143
                           , A => n4201, ZN => n4194);
   U5081 : OAI22_X1 port map( A1 => n47, A2 => n415, B1 => n503, B2 => n3316, 
                           ZN => n4201);
   U5082 : NAND4_X1 port map( A1 => n4202, A2 => n4203, A3 => n4204, A4 => 
                           n4205, ZN => n4183);
   U5083 : AOI221_X1 port map( B1 => n3321, B2 => n6090, C1 => n3322, C2 => 
                           n6122, A => n4206, ZN => n4205);
   U5084 : OAI222_X1 port map( A1 => n4874, A2 => n3324, B1 => n4842, B2 => 
                           n3325, C1 => n4810, C2 => n423, ZN => n4206);
   U5085 : AOI221_X1 port map( B1 => n3326, B2 => n784, C1 => n3327, C2 => n360
                           , A => n4207, ZN => n4204);
   U5086 : OAI22_X1 port map( A1 => n264, A2 => n3329, B1 => n688, B2 => n3330,
                           ZN => n4207);
   U5087 : AOI221_X1 port map( B1 => n3331, B2 => n6218, C1 => n3332, C2 => 
                           n6250, A => n4208, ZN => n4203);
   U5088 : OAI222_X1 port map( A1 => n4970, A2 => n3334, B1 => n4938, B2 => 
                           n3335, C1 => n4906, C2 => n3336, ZN => n4208);
   U5089 : AOI221_X1 port map( B1 => n3337, B2 => n600, C1 => n3338, C2 => n144
                           , A => n4209, ZN => n4202);
   U5090 : OAI22_X1 port map( A1 => n48, A2 => n3340, B1 => n504, B2 => n3341, 
                           ZN => n4209);
   U5091 : NAND4_X1 port map( A1 => n4210, A2 => n4211, A3 => n4212, A4 => 
                           n4213, ZN => n4182);
   U5092 : AOI221_X1 port map( B1 => n3346, B2 => n5834, C1 => n3347, C2 => 
                           n5866, A => n4214, ZN => n4213);
   U5093 : OAI222_X1 port map( A1 => n4618, A2 => n3349, B1 => n4586, B2 => 
                           n3350, C1 => n4554, C2 => n3351, ZN => n4214);
   U5094 : AOI221_X1 port map( B1 => n3352, B2 => n5898, C1 => n3353, C2 => 
                           n5930, A => n4215, ZN => n4212);
   U5095 : OAI22_X1 port map( A1 => n4682, A2 => n3355, B1 => n4650, B2 => 
                           n3356, ZN => n4215);
   U5096 : AOI221_X1 port map( B1 => n3357, B2 => n5962, C1 => n3358, C2 => 
                           n5994, A => n4216, ZN => n4211);
   U5097 : OAI222_X1 port map( A1 => n4778, A2 => n3360, B1 => n4746, B2 => 
                           n3361, C1 => n4714, C2 => n424, ZN => n4216);
   U5098 : AOI221_X1 port map( B1 => n3362, B2 => n6058, C1 => n3363, C2 => 
                           n6026, A => n4217, ZN => n4210);
   U5099 : OAI22_X1 port map( A1 => n5459, A2 => n3365, B1 => n5458, B2 => 
                           n3366, ZN => n4217);
   U5100 : INV_X1 port map( A => DATAIN(8), ZN => n2888);
   U5101 : OAI21_X1 port map( B1 => n3266, B2 => n1568, A => ENABLE, ZN => 
                           n7562);
   U5102 : OAI222_X1 port map( A1 => n2926, A2 => n3263, B1 => n4218, B2 => 
                           n3265, C1 => n3266, C2 => n1505, ZN => n7561);
   U5103 : NOR4_X1 port map( A1 => n4219, A2 => n4220, A3 => n4221, A4 => n4222
                           , ZN => n4218);
   U5104 : NAND4_X1 port map( A1 => n4223, A2 => n4224, A3 => n4225, A4 => 
                           n4226, ZN => n4222);
   U5105 : AOI221_X1 port map( B1 => n3275, B2 => n6409, C1 => n3276, C2 => 
                           n6441, A => n4227, ZN => n4226);
   U5106 : OAI222_X1 port map( A1 => n5257, A2 => n3278, B1 => n5225, B2 => 
                           n3279, C1 => n5193, C2 => n421, ZN => n4227);
   U5107 : AOI221_X1 port map( B1 => n3280, B2 => n785, C1 => n3281, C2 => n361
                           , A => n4228, ZN => n4225);
   U5108 : OAI22_X1 port map( A1 => n265, A2 => n413, B1 => n689, B2 => n3283, 
                           ZN => n4228);
   U5109 : AOI221_X1 port map( B1 => n3284, B2 => n6537, C1 => n3285, C2 => 
                           n6569, A => n4229, ZN => n4224);
   U5110 : OAI222_X1 port map( A1 => n5353, A2 => n3287, B1 => n5321, B2 => 
                           n1579, C1 => n5289, C2 => n3288, ZN => n4229);
   U5111 : AOI221_X1 port map( B1 => n3289, B2 => n786, C1 => n3290, C2 => n362
                           , A => n4230, ZN => n4223);
   U5112 : OAI22_X1 port map( A1 => n266, A2 => n414, B1 => n690, B2 => n3292, 
                           ZN => n4230);
   U5113 : NAND4_X1 port map( A1 => n4231, A2 => n4232, A3 => n4233, A4 => 
                           n4234, ZN => n4221);
   U5114 : AOI221_X1 port map( B1 => n3297, B2 => n6281, C1 => n3298, C2 => 
                           n6313, A => n4235, ZN => n4234);
   U5115 : OAI222_X1 port map( A1 => n5065, A2 => n3300, B1 => n5033, B2 => 
                           n3301, C1 => n5001, C2 => n3302, ZN => n4235);
   U5116 : AOI221_X1 port map( B1 => n3303, B2 => n545, C1 => n3304, C2 => n185
                           , A => n4236, ZN => n4233);
   U5117 : OAI22_X1 port map( A1 => n449, A2 => n3306, B1 => n89, B2 => n3307, 
                           ZN => n4236);
   U5118 : AOI221_X1 port map( B1 => n3308, B2 => n6345, C1 => n3309, C2 => 
                           n6377, A => n4237, ZN => n4232);
   U5119 : OAI222_X1 port map( A1 => n5161, A2 => n3311, B1 => n5129, B2 => 
                           n3312, C1 => n5097, C2 => n422, ZN => n4237);
   U5120 : AOI221_X1 port map( B1 => n3313, B2 => n601, C1 => n3314, C2 => n145
                           , A => n4238, ZN => n4231);
   U5121 : OAI22_X1 port map( A1 => n49, A2 => n415, B1 => n505, B2 => n3316, 
                           ZN => n4238);
   U5122 : NAND4_X1 port map( A1 => n4239, A2 => n4240, A3 => n4241, A4 => 
                           n4242, ZN => n4220);
   U5123 : AOI221_X1 port map( B1 => n3321, B2 => n6089, C1 => n3322, C2 => 
                           n6121, A => n4243, ZN => n4242);
   U5124 : OAI222_X1 port map( A1 => n4873, A2 => n3324, B1 => n4841, B2 => 
                           n3325, C1 => n4809, C2 => n423, ZN => n4243);
   U5125 : AOI221_X1 port map( B1 => n3326, B2 => n787, C1 => n3327, C2 => n363
                           , A => n4244, ZN => n4241);
   U5126 : OAI22_X1 port map( A1 => n267, A2 => n3329, B1 => n691, B2 => n3330,
                           ZN => n4244);
   U5127 : AOI221_X1 port map( B1 => n3331, B2 => n6217, C1 => n3332, C2 => 
                           n6249, A => n4245, ZN => n4240);
   U5128 : OAI222_X1 port map( A1 => n4969, A2 => n3334, B1 => n4937, B2 => 
                           n3335, C1 => n4905, C2 => n3336, ZN => n4245);
   U5129 : AOI221_X1 port map( B1 => n3337, B2 => n602, C1 => n3338, C2 => n146
                           , A => n4246, ZN => n4239);
   U5130 : OAI22_X1 port map( A1 => n50, A2 => n3340, B1 => n506, B2 => n3341, 
                           ZN => n4246);
   U5131 : NAND4_X1 port map( A1 => n4247, A2 => n4248, A3 => n4249, A4 => 
                           n4250, ZN => n4219);
   U5132 : AOI221_X1 port map( B1 => n3346, B2 => n5833, C1 => n3347, C2 => 
                           n5865, A => n4251, ZN => n4250);
   U5133 : OAI222_X1 port map( A1 => n4617, A2 => n3349, B1 => n4585, B2 => 
                           n3350, C1 => n4553, C2 => n3351, ZN => n4251);
   U5134 : AOI221_X1 port map( B1 => n3352, B2 => n5897, C1 => n3353, C2 => 
                           n5929, A => n4252, ZN => n4249);
   U5135 : OAI22_X1 port map( A1 => n4681, A2 => n3355, B1 => n4649, B2 => 
                           n3356, ZN => n4252);
   U5136 : AOI221_X1 port map( B1 => n3357, B2 => n5961, C1 => n3358, C2 => 
                           n5993, A => n4253, ZN => n4248);
   U5137 : OAI222_X1 port map( A1 => n4777, A2 => n3360, B1 => n4745, B2 => 
                           n3361, C1 => n4713, C2 => n424, ZN => n4253);
   U5138 : AOI221_X1 port map( B1 => n3362, B2 => n6057, C1 => n3363, C2 => 
                           n6025, A => n4254, ZN => n4247);
   U5139 : OAI22_X1 port map( A1 => n5449, A2 => n3365, B1 => n5448, B2 => 
                           n3366, ZN => n4254);
   U5140 : INV_X1 port map( A => DATAIN(7), ZN => n2926);
   U5141 : OAI21_X1 port map( B1 => n3266, B2 => n1569, A => ENABLE, ZN => 
                           n7560);
   U5142 : OAI222_X1 port map( A1 => n2964, A2 => n3263, B1 => n4255, B2 => 
                           n3265, C1 => n3266, C2 => n1506, ZN => n7559);
   U5143 : NOR4_X1 port map( A1 => n4256, A2 => n4257, A3 => n4258, A4 => n4259
                           , ZN => n4255);
   U5144 : NAND4_X1 port map( A1 => n4260, A2 => n4261, A3 => n4262, A4 => 
                           n4263, ZN => n4259);
   U5145 : AOI221_X1 port map( B1 => n3275, B2 => n6408, C1 => n3276, C2 => 
                           n6440, A => n4264, ZN => n4263);
   U5146 : OAI222_X1 port map( A1 => n5256, A2 => n3278, B1 => n5224, B2 => 
                           n3279, C1 => n5192, C2 => n421, ZN => n4264);
   U5147 : AOI221_X1 port map( B1 => n3280, B2 => n788, C1 => n3281, C2 => n364
                           , A => n4265, ZN => n4262);
   U5148 : OAI22_X1 port map( A1 => n268, A2 => n413, B1 => n692, B2 => n3283, 
                           ZN => n4265);
   U5149 : AOI221_X1 port map( B1 => n3284, B2 => n6536, C1 => n3285, C2 => 
                           n6568, A => n4266, ZN => n4261);
   U5150 : OAI222_X1 port map( A1 => n5352, A2 => n3287, B1 => n5320, B2 => 
                           n1579, C1 => n5288, C2 => n3288, ZN => n4266);
   U5151 : AOI221_X1 port map( B1 => n3289, B2 => n789, C1 => n3290, C2 => n365
                           , A => n4267, ZN => n4260);
   U5152 : OAI22_X1 port map( A1 => n269, A2 => n414, B1 => n693, B2 => n3292, 
                           ZN => n4267);
   U5153 : NAND4_X1 port map( A1 => n4268, A2 => n4269, A3 => n4270, A4 => 
                           n4271, ZN => n4258);
   U5154 : AOI221_X1 port map( B1 => n3297, B2 => n6280, C1 => n3298, C2 => 
                           n6312, A => n4272, ZN => n4271);
   U5155 : OAI222_X1 port map( A1 => n5064, A2 => n3300, B1 => n5032, B2 => 
                           n3301, C1 => n5000, C2 => n3302, ZN => n4272);
   U5156 : AOI221_X1 port map( B1 => n3303, B2 => n546, C1 => n3304, C2 => n186
                           , A => n4273, ZN => n4270);
   U5157 : OAI22_X1 port map( A1 => n450, A2 => n3306, B1 => n90, B2 => n3307, 
                           ZN => n4273);
   U5158 : AOI221_X1 port map( B1 => n3308, B2 => n6344, C1 => n3309, C2 => 
                           n6376, A => n4274, ZN => n4269);
   U5159 : OAI222_X1 port map( A1 => n5160, A2 => n3311, B1 => n5128, B2 => 
                           n3312, C1 => n5096, C2 => n422, ZN => n4274);
   U5160 : AOI221_X1 port map( B1 => n3313, B2 => n603, C1 => n3314, C2 => n147
                           , A => n4275, ZN => n4268);
   U5161 : OAI22_X1 port map( A1 => n51, A2 => n415, B1 => n507, B2 => n3316, 
                           ZN => n4275);
   U5162 : NAND4_X1 port map( A1 => n4276, A2 => n4277, A3 => n4278, A4 => 
                           n4279, ZN => n4257);
   U5163 : AOI221_X1 port map( B1 => n3321, B2 => n6088, C1 => n3322, C2 => 
                           n6120, A => n4280, ZN => n4279);
   U5164 : OAI222_X1 port map( A1 => n4872, A2 => n3324, B1 => n4840, B2 => 
                           n3325, C1 => n4808, C2 => n423, ZN => n4280);
   U5165 : AOI221_X1 port map( B1 => n3326, B2 => n790, C1 => n3327, C2 => n366
                           , A => n4281, ZN => n4278);
   U5166 : OAI22_X1 port map( A1 => n270, A2 => n3329, B1 => n694, B2 => n3330,
                           ZN => n4281);
   U5167 : AOI221_X1 port map( B1 => n3331, B2 => n6216, C1 => n3332, C2 => 
                           n6248, A => n4282, ZN => n4277);
   U5168 : OAI222_X1 port map( A1 => n4968, A2 => n3334, B1 => n4936, B2 => 
                           n3335, C1 => n4904, C2 => n3336, ZN => n4282);
   U5169 : AOI221_X1 port map( B1 => n3337, B2 => n604, C1 => n3338, C2 => n148
                           , A => n4283, ZN => n4276);
   U5170 : OAI22_X1 port map( A1 => n52, A2 => n3340, B1 => n508, B2 => n3341, 
                           ZN => n4283);
   U5171 : NAND4_X1 port map( A1 => n4284, A2 => n4285, A3 => n4286, A4 => 
                           n4287, ZN => n4256);
   U5172 : AOI221_X1 port map( B1 => n3346, B2 => n5832, C1 => n3347, C2 => 
                           n5864, A => n4288, ZN => n4287);
   U5173 : OAI222_X1 port map( A1 => n4616, A2 => n3349, B1 => n4584, B2 => 
                           n3350, C1 => n4552, C2 => n3351, ZN => n4288);
   U5174 : AOI221_X1 port map( B1 => n3352, B2 => n5896, C1 => n3353, C2 => 
                           n5928, A => n4289, ZN => n4286);
   U5175 : OAI22_X1 port map( A1 => n4680, A2 => n3355, B1 => n4648, B2 => 
                           n3356, ZN => n4289);
   U5176 : AOI221_X1 port map( B1 => n3357, B2 => n5960, C1 => n3358, C2 => 
                           n5992, A => n4290, ZN => n4285);
   U5177 : OAI222_X1 port map( A1 => n4776, A2 => n3360, B1 => n4744, B2 => 
                           n3361, C1 => n4712, C2 => n424, ZN => n4290);
   U5178 : AOI221_X1 port map( B1 => n3362, B2 => n6056, C1 => n3363, C2 => 
                           n6024, A => n4291, ZN => n4284);
   U5179 : OAI22_X1 port map( A1 => n5439, A2 => n3365, B1 => n5438, B2 => 
                           n3366, ZN => n4291);
   U5180 : INV_X1 port map( A => DATAIN(6), ZN => n2964);
   U5181 : OAI21_X1 port map( B1 => n3266, B2 => n1570, A => ENABLE, ZN => 
                           n7558);
   U5182 : OAI222_X1 port map( A1 => n3002, A2 => n3263, B1 => n4292, B2 => 
                           n3265, C1 => n3266, C2 => n1507, ZN => n7557);
   U5183 : NOR4_X1 port map( A1 => n4293, A2 => n4294, A3 => n4295, A4 => n4296
                           , ZN => n4292);
   U5184 : NAND4_X1 port map( A1 => n4297, A2 => n4298, A3 => n4299, A4 => 
                           n4300, ZN => n4296);
   U5185 : AOI221_X1 port map( B1 => n3275, B2 => n6407, C1 => n3276, C2 => 
                           n6439, A => n4301, ZN => n4300);
   U5186 : OAI222_X1 port map( A1 => n5255, A2 => n3278, B1 => n5223, B2 => 
                           n3279, C1 => n5191, C2 => n421, ZN => n4301);
   U5187 : AOI221_X1 port map( B1 => n3280, B2 => n791, C1 => n3281, C2 => n367
                           , A => n4302, ZN => n4299);
   U5188 : OAI22_X1 port map( A1 => n271, A2 => n413, B1 => n695, B2 => n3283, 
                           ZN => n4302);
   U5189 : AOI221_X1 port map( B1 => n3284, B2 => n6535, C1 => n3285, C2 => 
                           n6567, A => n4303, ZN => n4298);
   U5190 : OAI222_X1 port map( A1 => n5351, A2 => n3287, B1 => n5319, B2 => 
                           n1579, C1 => n5287, C2 => n3288, ZN => n4303);
   U5191 : AOI221_X1 port map( B1 => n3289, B2 => n792, C1 => n3290, C2 => n368
                           , A => n4304, ZN => n4297);
   U5192 : OAI22_X1 port map( A1 => n272, A2 => n414, B1 => n696, B2 => n3292, 
                           ZN => n4304);
   U5193 : NAND4_X1 port map( A1 => n4305, A2 => n4306, A3 => n4307, A4 => 
                           n4308, ZN => n4295);
   U5194 : AOI221_X1 port map( B1 => n3297, B2 => n6279, C1 => n3298, C2 => 
                           n6311, A => n4309, ZN => n4308);
   U5195 : OAI222_X1 port map( A1 => n5063, A2 => n3300, B1 => n5031, B2 => 
                           n3301, C1 => n4999, C2 => n3302, ZN => n4309);
   U5196 : AOI221_X1 port map( B1 => n3303, B2 => n547, C1 => n3304, C2 => n187
                           , A => n4310, ZN => n4307);
   U5197 : OAI22_X1 port map( A1 => n451, A2 => n3306, B1 => n91, B2 => n3307, 
                           ZN => n4310);
   U5198 : AOI221_X1 port map( B1 => n3308, B2 => n6343, C1 => n3309, C2 => 
                           n6375, A => n4311, ZN => n4306);
   U5199 : OAI222_X1 port map( A1 => n5159, A2 => n3311, B1 => n5127, B2 => 
                           n3312, C1 => n5095, C2 => n422, ZN => n4311);
   U5200 : AOI221_X1 port map( B1 => n3313, B2 => n605, C1 => n3314, C2 => n149
                           , A => n4312, ZN => n4305);
   U5201 : OAI22_X1 port map( A1 => n53, A2 => n415, B1 => n509, B2 => n3316, 
                           ZN => n4312);
   U5202 : NAND4_X1 port map( A1 => n4313, A2 => n4314, A3 => n4315, A4 => 
                           n4316, ZN => n4294);
   U5203 : AOI221_X1 port map( B1 => n3321, B2 => n6087, C1 => n3322, C2 => 
                           n6119, A => n4317, ZN => n4316);
   U5204 : OAI222_X1 port map( A1 => n4871, A2 => n3324, B1 => n4839, B2 => 
                           n3325, C1 => n4807, C2 => n423, ZN => n4317);
   U5205 : AOI221_X1 port map( B1 => n3326, B2 => n793, C1 => n3327, C2 => n369
                           , A => n4318, ZN => n4315);
   U5206 : OAI22_X1 port map( A1 => n273, A2 => n3329, B1 => n697, B2 => n3330,
                           ZN => n4318);
   U5207 : AOI221_X1 port map( B1 => n3331, B2 => n6215, C1 => n3332, C2 => 
                           n6247, A => n4319, ZN => n4314);
   U5208 : OAI222_X1 port map( A1 => n4967, A2 => n3334, B1 => n4935, B2 => 
                           n3335, C1 => n4903, C2 => n3336, ZN => n4319);
   U5209 : AOI221_X1 port map( B1 => n3337, B2 => n606, C1 => n3338, C2 => n150
                           , A => n4320, ZN => n4313);
   U5210 : OAI22_X1 port map( A1 => n54, A2 => n3340, B1 => n510, B2 => n3341, 
                           ZN => n4320);
   U5211 : NAND4_X1 port map( A1 => n4321, A2 => n4322, A3 => n4323, A4 => 
                           n4324, ZN => n4293);
   U5212 : AOI221_X1 port map( B1 => n3346, B2 => n5831, C1 => n3347, C2 => 
                           n5863, A => n4325, ZN => n4324);
   U5213 : OAI222_X1 port map( A1 => n4615, A2 => n3349, B1 => n4583, B2 => 
                           n3350, C1 => n4551, C2 => n3351, ZN => n4325);
   U5214 : AOI221_X1 port map( B1 => n3352, B2 => n5895, C1 => n3353, C2 => 
                           n5927, A => n4326, ZN => n4323);
   U5215 : OAI22_X1 port map( A1 => n4679, A2 => n3355, B1 => n4647, B2 => 
                           n3356, ZN => n4326);
   U5216 : AOI221_X1 port map( B1 => n3357, B2 => n5959, C1 => n3358, C2 => 
                           n5991, A => n4327, ZN => n4322);
   U5217 : OAI222_X1 port map( A1 => n4775, A2 => n3360, B1 => n4743, B2 => 
                           n3361, C1 => n4711, C2 => n424, ZN => n4327);
   U5218 : AOI221_X1 port map( B1 => n3362, B2 => n6055, C1 => n3363, C2 => 
                           n6023, A => n4328, ZN => n4321);
   U5219 : OAI22_X1 port map( A1 => n5429, A2 => n3365, B1 => n5428, B2 => 
                           n3366, ZN => n4328);
   U5220 : INV_X1 port map( A => DATAIN(5), ZN => n3002);
   U5221 : OAI21_X1 port map( B1 => n3266, B2 => n1571, A => ENABLE, ZN => 
                           n7556);
   U5222 : OAI222_X1 port map( A1 => n3040, A2 => n3263, B1 => n4329, B2 => 
                           n3265, C1 => n3266, C2 => n1508, ZN => n7555);
   U5223 : NOR4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => n4333
                           , ZN => n4329);
   U5224 : NAND4_X1 port map( A1 => n4334, A2 => n4335, A3 => n4336, A4 => 
                           n4337, ZN => n4333);
   U5225 : AOI221_X1 port map( B1 => n3275, B2 => n6406, C1 => n3276, C2 => 
                           n6438, A => n4338, ZN => n4337);
   U5226 : OAI222_X1 port map( A1 => n5254, A2 => n3278, B1 => n5222, B2 => 
                           n3279, C1 => n5190, C2 => n421, ZN => n4338);
   U5227 : AOI221_X1 port map( B1 => n3280, B2 => n794, C1 => n3281, C2 => n370
                           , A => n4339, ZN => n4336);
   U5228 : OAI22_X1 port map( A1 => n274, A2 => n413, B1 => n698, B2 => n3283, 
                           ZN => n4339);
   U5229 : AOI221_X1 port map( B1 => n3284, B2 => n6534, C1 => n3285, C2 => 
                           n6566, A => n4340, ZN => n4335);
   U5230 : OAI222_X1 port map( A1 => n5350, A2 => n3287, B1 => n5318, B2 => 
                           n1579, C1 => n5286, C2 => n3288, ZN => n4340);
   U5231 : AOI221_X1 port map( B1 => n3289, B2 => n795, C1 => n3290, C2 => n371
                           , A => n4341, ZN => n4334);
   U5232 : OAI22_X1 port map( A1 => n275, A2 => n414, B1 => n699, B2 => n3292, 
                           ZN => n4341);
   U5233 : NAND4_X1 port map( A1 => n4342, A2 => n4343, A3 => n4344, A4 => 
                           n4345, ZN => n4332);
   U5234 : AOI221_X1 port map( B1 => n3297, B2 => n6278, C1 => n3298, C2 => 
                           n6310, A => n4346, ZN => n4345);
   U5235 : OAI222_X1 port map( A1 => n5062, A2 => n3300, B1 => n5030, B2 => 
                           n3301, C1 => n4998, C2 => n3302, ZN => n4346);
   U5236 : AOI221_X1 port map( B1 => n3303, B2 => n548, C1 => n3304, C2 => n188
                           , A => n4347, ZN => n4344);
   U5237 : OAI22_X1 port map( A1 => n452, A2 => n3306, B1 => n92, B2 => n3307, 
                           ZN => n4347);
   U5238 : AOI221_X1 port map( B1 => n3308, B2 => n6342, C1 => n3309, C2 => 
                           n6374, A => n4348, ZN => n4343);
   U5239 : OAI222_X1 port map( A1 => n5158, A2 => n3311, B1 => n5126, B2 => 
                           n3312, C1 => n5094, C2 => n422, ZN => n4348);
   U5240 : AOI221_X1 port map( B1 => n3313, B2 => n607, C1 => n3314, C2 => n151
                           , A => n4349, ZN => n4342);
   U5241 : OAI22_X1 port map( A1 => n55, A2 => n415, B1 => n511, B2 => n3316, 
                           ZN => n4349);
   U5242 : NAND4_X1 port map( A1 => n4350, A2 => n4351, A3 => n4352, A4 => 
                           n4353, ZN => n4331);
   U5243 : AOI221_X1 port map( B1 => n3321, B2 => n6086, C1 => n3322, C2 => 
                           n6118, A => n4354, ZN => n4353);
   U5244 : OAI222_X1 port map( A1 => n4870, A2 => n3324, B1 => n4838, B2 => 
                           n3325, C1 => n4806, C2 => n423, ZN => n4354);
   U5245 : AOI221_X1 port map( B1 => n3326, B2 => n796, C1 => n3327, C2 => n372
                           , A => n4355, ZN => n4352);
   U5246 : OAI22_X1 port map( A1 => n276, A2 => n3329, B1 => n700, B2 => n3330,
                           ZN => n4355);
   U5247 : AOI221_X1 port map( B1 => n3331, B2 => n6214, C1 => n3332, C2 => 
                           n6246, A => n4356, ZN => n4351);
   U5248 : OAI222_X1 port map( A1 => n4966, A2 => n3334, B1 => n4934, B2 => 
                           n3335, C1 => n4902, C2 => n3336, ZN => n4356);
   U5249 : AOI221_X1 port map( B1 => n3337, B2 => n608, C1 => n3338, C2 => n152
                           , A => n4357, ZN => n4350);
   U5250 : OAI22_X1 port map( A1 => n56, A2 => n3340, B1 => n512, B2 => n3341, 
                           ZN => n4357);
   U5251 : NAND4_X1 port map( A1 => n4358, A2 => n4359, A3 => n4360, A4 => 
                           n4361, ZN => n4330);
   U5252 : AOI221_X1 port map( B1 => n3346, B2 => n5830, C1 => n3347, C2 => 
                           n5862, A => n4362, ZN => n4361);
   U5253 : OAI222_X1 port map( A1 => n4614, A2 => n3349, B1 => n4582, B2 => 
                           n3350, C1 => n4550, C2 => n3351, ZN => n4362);
   U5254 : AOI221_X1 port map( B1 => n3352, B2 => n5894, C1 => n3353, C2 => 
                           n5926, A => n4363, ZN => n4360);
   U5255 : OAI22_X1 port map( A1 => n4678, A2 => n3355, B1 => n4646, B2 => 
                           n3356, ZN => n4363);
   U5256 : AOI221_X1 port map( B1 => n3357, B2 => n5958, C1 => n3358, C2 => 
                           n5990, A => n4364, ZN => n4359);
   U5257 : OAI222_X1 port map( A1 => n4774, A2 => n3360, B1 => n4742, B2 => 
                           n3361, C1 => n4710, C2 => n424, ZN => n4364);
   U5258 : AOI221_X1 port map( B1 => n3362, B2 => n6054, C1 => n3363, C2 => 
                           n6022, A => n4365, ZN => n4358);
   U5259 : OAI22_X1 port map( A1 => n5419, A2 => n3365, B1 => n5418, B2 => 
                           n3366, ZN => n4365);
   U5260 : INV_X1 port map( A => DATAIN(4), ZN => n3040);
   U5261 : OAI21_X1 port map( B1 => n3266, B2 => n1572, A => ENABLE, ZN => 
                           n7554);
   U5262 : OAI222_X1 port map( A1 => n3078, A2 => n3263, B1 => n4366, B2 => 
                           n3265, C1 => n3266, C2 => n1509, ZN => n7553);
   U5263 : NOR4_X1 port map( A1 => n4367, A2 => n4368, A3 => n4369, A4 => n4370
                           , ZN => n4366);
   U5264 : NAND4_X1 port map( A1 => n4371, A2 => n4372, A3 => n4373, A4 => 
                           n4374, ZN => n4370);
   U5265 : AOI221_X1 port map( B1 => n3275, B2 => n6405, C1 => n3276, C2 => 
                           n6437, A => n4375, ZN => n4374);
   U5266 : OAI222_X1 port map( A1 => n5253, A2 => n3278, B1 => n5221, B2 => 
                           n3279, C1 => n5189, C2 => n421, ZN => n4375);
   U5267 : AOI221_X1 port map( B1 => n3280, B2 => n797, C1 => n3281, C2 => n373
                           , A => n4376, ZN => n4373);
   U5268 : OAI22_X1 port map( A1 => n277, A2 => n413, B1 => n701, B2 => n3283, 
                           ZN => n4376);
   U5269 : AOI221_X1 port map( B1 => n3284, B2 => n6533, C1 => n3285, C2 => 
                           n6565, A => n4377, ZN => n4372);
   U5270 : OAI222_X1 port map( A1 => n5349, A2 => n3287, B1 => n5317, B2 => 
                           n1579, C1 => n5285, C2 => n3288, ZN => n4377);
   U5271 : AOI221_X1 port map( B1 => n3289, B2 => n798, C1 => n3290, C2 => n374
                           , A => n4378, ZN => n4371);
   U5272 : OAI22_X1 port map( A1 => n278, A2 => n414, B1 => n702, B2 => n3292, 
                           ZN => n4378);
   U5273 : NAND4_X1 port map( A1 => n4379, A2 => n4380, A3 => n4381, A4 => 
                           n4382, ZN => n4369);
   U5274 : AOI221_X1 port map( B1 => n3297, B2 => n6277, C1 => n3298, C2 => 
                           n6309, A => n4383, ZN => n4382);
   U5275 : OAI222_X1 port map( A1 => n5061, A2 => n3300, B1 => n5029, B2 => 
                           n3301, C1 => n4997, C2 => n3302, ZN => n4383);
   U5276 : AOI221_X1 port map( B1 => n3303, B2 => n549, C1 => n3304, C2 => n189
                           , A => n4384, ZN => n4381);
   U5277 : OAI22_X1 port map( A1 => n453, A2 => n3306, B1 => n93, B2 => n3307, 
                           ZN => n4384);
   U5278 : AOI221_X1 port map( B1 => n3308, B2 => n6341, C1 => n3309, C2 => 
                           n6373, A => n4385, ZN => n4380);
   U5279 : OAI222_X1 port map( A1 => n5157, A2 => n3311, B1 => n5125, B2 => 
                           n3312, C1 => n5093, C2 => n422, ZN => n4385);
   U5280 : AOI221_X1 port map( B1 => n3313, B2 => n609, C1 => n3314, C2 => n153
                           , A => n4386, ZN => n4379);
   U5281 : OAI22_X1 port map( A1 => n57, A2 => n415, B1 => n513, B2 => n3316, 
                           ZN => n4386);
   U5282 : NAND4_X1 port map( A1 => n4387, A2 => n4388, A3 => n4389, A4 => 
                           n4390, ZN => n4368);
   U5283 : AOI221_X1 port map( B1 => n3321, B2 => n6085, C1 => n3322, C2 => 
                           n6117, A => n4391, ZN => n4390);
   U5284 : OAI222_X1 port map( A1 => n4869, A2 => n3324, B1 => n4837, B2 => 
                           n3325, C1 => n4805, C2 => n423, ZN => n4391);
   U5285 : AOI221_X1 port map( B1 => n3326, B2 => n799, C1 => n3327, C2 => n375
                           , A => n4392, ZN => n4389);
   U5286 : OAI22_X1 port map( A1 => n279, A2 => n3329, B1 => n703, B2 => n3330,
                           ZN => n4392);
   U5287 : AOI221_X1 port map( B1 => n3331, B2 => n6213, C1 => n3332, C2 => 
                           n6245, A => n4393, ZN => n4388);
   U5288 : OAI222_X1 port map( A1 => n4965, A2 => n3334, B1 => n4933, B2 => 
                           n3335, C1 => n4901, C2 => n3336, ZN => n4393);
   U5289 : AOI221_X1 port map( B1 => n3337, B2 => n610, C1 => n3338, C2 => n154
                           , A => n4394, ZN => n4387);
   U5290 : OAI22_X1 port map( A1 => n58, A2 => n3340, B1 => n514, B2 => n3341, 
                           ZN => n4394);
   U5291 : NAND4_X1 port map( A1 => n4395, A2 => n4396, A3 => n4397, A4 => 
                           n4398, ZN => n4367);
   U5292 : AOI221_X1 port map( B1 => n3346, B2 => n5829, C1 => n3347, C2 => 
                           n5861, A => n4399, ZN => n4398);
   U5293 : OAI222_X1 port map( A1 => n4613, A2 => n3349, B1 => n4581, B2 => 
                           n3350, C1 => n4549, C2 => n3351, ZN => n4399);
   U5294 : AOI221_X1 port map( B1 => n3352, B2 => n5893, C1 => n3353, C2 => 
                           n5925, A => n4400, ZN => n4397);
   U5295 : OAI22_X1 port map( A1 => n4677, A2 => n3355, B1 => n4645, B2 => 
                           n3356, ZN => n4400);
   U5296 : AOI221_X1 port map( B1 => n3357, B2 => n5957, C1 => n3358, C2 => 
                           n5989, A => n4401, ZN => n4396);
   U5297 : OAI222_X1 port map( A1 => n4773, A2 => n3360, B1 => n4741, B2 => 
                           n3361, C1 => n4709, C2 => n424, ZN => n4401);
   U5298 : AOI221_X1 port map( B1 => n3362, B2 => n6053, C1 => n3363, C2 => 
                           n6021, A => n4402, ZN => n4395);
   U5299 : OAI22_X1 port map( A1 => n5409, A2 => n3365, B1 => n5408, B2 => 
                           n3366, ZN => n4402);
   U5300 : INV_X1 port map( A => DATAIN(3), ZN => n3078);
   U5301 : OAI21_X1 port map( B1 => n3266, B2 => n1573, A => ENABLE, ZN => 
                           n7552);
   U5302 : OAI222_X1 port map( A1 => n3116, A2 => n3263, B1 => n4403, B2 => 
                           n3265, C1 => n3266, C2 => n1510, ZN => n7551);
   U5303 : NOR4_X1 port map( A1 => n4404, A2 => n4405, A3 => n4406, A4 => n4407
                           , ZN => n4403);
   U5304 : NAND4_X1 port map( A1 => n4408, A2 => n4409, A3 => n4410, A4 => 
                           n4411, ZN => n4407);
   U5305 : AOI221_X1 port map( B1 => n3275, B2 => n6404, C1 => n3276, C2 => 
                           n6436, A => n4412, ZN => n4411);
   U5306 : OAI222_X1 port map( A1 => n5252, A2 => n3278, B1 => n5220, B2 => 
                           n3279, C1 => n5188, C2 => n421, ZN => n4412);
   U5307 : AOI221_X1 port map( B1 => n3280, B2 => n800, C1 => n3281, C2 => n376
                           , A => n4413, ZN => n4410);
   U5308 : OAI22_X1 port map( A1 => n280, A2 => n413, B1 => n704, B2 => n3283, 
                           ZN => n4413);
   U5309 : AOI221_X1 port map( B1 => n3284, B2 => n6532, C1 => n3285, C2 => 
                           n6564, A => n4414, ZN => n4409);
   U5310 : OAI222_X1 port map( A1 => n5348, A2 => n3287, B1 => n5316, B2 => 
                           n1579, C1 => n5284, C2 => n3288, ZN => n4414);
   U5311 : AOI221_X1 port map( B1 => n3289, B2 => n801, C1 => n3290, C2 => n377
                           , A => n4415, ZN => n4408);
   U5312 : OAI22_X1 port map( A1 => n281, A2 => n414, B1 => n705, B2 => n3292, 
                           ZN => n4415);
   U5313 : NAND4_X1 port map( A1 => n4416, A2 => n4417, A3 => n4418, A4 => 
                           n4419, ZN => n4406);
   U5314 : AOI221_X1 port map( B1 => n3297, B2 => n6276, C1 => n3298, C2 => 
                           n6308, A => n4420, ZN => n4419);
   U5315 : OAI222_X1 port map( A1 => n5060, A2 => n3300, B1 => n5028, B2 => 
                           n3301, C1 => n4996, C2 => n3302, ZN => n4420);
   U5316 : AOI221_X1 port map( B1 => n3303, B2 => n550, C1 => n3304, C2 => n190
                           , A => n4421, ZN => n4418);
   U5317 : OAI22_X1 port map( A1 => n454, A2 => n3306, B1 => n94, B2 => n3307, 
                           ZN => n4421);
   U5318 : AOI221_X1 port map( B1 => n3308, B2 => n6340, C1 => n3309, C2 => 
                           n6372, A => n4422, ZN => n4417);
   U5319 : OAI222_X1 port map( A1 => n5156, A2 => n3311, B1 => n5124, B2 => 
                           n3312, C1 => n5092, C2 => n422, ZN => n4422);
   U5320 : AOI221_X1 port map( B1 => n3313, B2 => n611, C1 => n3314, C2 => n155
                           , A => n4423, ZN => n4416);
   U5321 : OAI22_X1 port map( A1 => n59, A2 => n415, B1 => n515, B2 => n3316, 
                           ZN => n4423);
   U5322 : NAND4_X1 port map( A1 => n4424, A2 => n4425, A3 => n4426, A4 => 
                           n4427, ZN => n4405);
   U5323 : AOI221_X1 port map( B1 => n3321, B2 => n6084, C1 => n3322, C2 => 
                           n6116, A => n4428, ZN => n4427);
   U5324 : OAI222_X1 port map( A1 => n4868, A2 => n3324, B1 => n4836, B2 => 
                           n3325, C1 => n4804, C2 => n423, ZN => n4428);
   U5325 : AOI221_X1 port map( B1 => n3326, B2 => n802, C1 => n3327, C2 => n378
                           , A => n4429, ZN => n4426);
   U5326 : OAI22_X1 port map( A1 => n282, A2 => n3329, B1 => n706, B2 => n3330,
                           ZN => n4429);
   U5327 : AOI221_X1 port map( B1 => n3331, B2 => n6212, C1 => n3332, C2 => 
                           n6244, A => n4430, ZN => n4425);
   U5328 : OAI222_X1 port map( A1 => n4964, A2 => n3334, B1 => n4932, B2 => 
                           n3335, C1 => n4900, C2 => n3336, ZN => n4430);
   U5329 : AOI221_X1 port map( B1 => n3337, B2 => n612, C1 => n3338, C2 => n156
                           , A => n4431, ZN => n4424);
   U5330 : OAI22_X1 port map( A1 => n60, A2 => n3340, B1 => n516, B2 => n3341, 
                           ZN => n4431);
   U5331 : NAND4_X1 port map( A1 => n4432, A2 => n4433, A3 => n4434, A4 => 
                           n4435, ZN => n4404);
   U5332 : AOI221_X1 port map( B1 => n3346, B2 => n5828, C1 => n3347, C2 => 
                           n5860, A => n4436, ZN => n4435);
   U5333 : OAI222_X1 port map( A1 => n4612, A2 => n3349, B1 => n4580, B2 => 
                           n3350, C1 => n4548, C2 => n3351, ZN => n4436);
   U5334 : AOI221_X1 port map( B1 => n3352, B2 => n5892, C1 => n3353, C2 => 
                           n5924, A => n4437, ZN => n4434);
   U5335 : OAI22_X1 port map( A1 => n4676, A2 => n3355, B1 => n4644, B2 => 
                           n3356, ZN => n4437);
   U5336 : AOI221_X1 port map( B1 => n3357, B2 => n5956, C1 => n3358, C2 => 
                           n5988, A => n4438, ZN => n4433);
   U5337 : OAI222_X1 port map( A1 => n4772, A2 => n3360, B1 => n4740, B2 => 
                           n3361, C1 => n4708, C2 => n424, ZN => n4438);
   U5338 : AOI221_X1 port map( B1 => n3362, B2 => n6052, C1 => n3363, C2 => 
                           n6020, A => n4439, ZN => n4432);
   U5339 : OAI22_X1 port map( A1 => n5399, A2 => n3365, B1 => n5398, B2 => 
                           n3366, ZN => n4439);
   U5340 : INV_X1 port map( A => DATAIN(2), ZN => n3116);
   U5341 : OAI21_X1 port map( B1 => n3266, B2 => n1574, A => ENABLE, ZN => 
                           n7550);
   U5342 : OAI222_X1 port map( A1 => n3154, A2 => n3263, B1 => n4440, B2 => 
                           n3265, C1 => n3266, C2 => n1511, ZN => n7549);
   U5343 : NOR4_X1 port map( A1 => n4441, A2 => n4442, A3 => n4443, A4 => n4444
                           , ZN => n4440);
   U5344 : NAND4_X1 port map( A1 => n4445, A2 => n4446, A3 => n4447, A4 => 
                           n4448, ZN => n4444);
   U5345 : AOI221_X1 port map( B1 => n3275, B2 => n6403, C1 => n3276, C2 => 
                           n6435, A => n4449, ZN => n4448);
   U5346 : OAI222_X1 port map( A1 => n5251, A2 => n3278, B1 => n5219, B2 => 
                           n3279, C1 => n5187, C2 => n421, ZN => n4449);
   U5347 : AOI221_X1 port map( B1 => n3280, B2 => n803, C1 => n3281, C2 => n379
                           , A => n4450, ZN => n4447);
   U5348 : OAI22_X1 port map( A1 => n283, A2 => n413, B1 => n707, B2 => n3283, 
                           ZN => n4450);
   U5349 : AOI221_X1 port map( B1 => n3284, B2 => n6531, C1 => n3285, C2 => 
                           n6563, A => n4451, ZN => n4446);
   U5350 : OAI222_X1 port map( A1 => n5347, A2 => n3287, B1 => n5315, B2 => 
                           n1579, C1 => n5283, C2 => n3288, ZN => n4451);
   U5351 : AOI221_X1 port map( B1 => n3289, B2 => n804, C1 => n3290, C2 => n380
                           , A => n4452, ZN => n4445);
   U5352 : OAI22_X1 port map( A1 => n284, A2 => n414, B1 => n708, B2 => n3292, 
                           ZN => n4452);
   U5353 : NAND4_X1 port map( A1 => n4453, A2 => n4454, A3 => n4455, A4 => 
                           n4456, ZN => n4443);
   U5354 : AOI221_X1 port map( B1 => n3297, B2 => n6275, C1 => n3298, C2 => 
                           n6307, A => n4457, ZN => n4456);
   U5355 : OAI222_X1 port map( A1 => n5059, A2 => n3300, B1 => n5027, B2 => 
                           n3301, C1 => n4995, C2 => n3302, ZN => n4457);
   U5356 : AOI221_X1 port map( B1 => n3303, B2 => n551, C1 => n3304, C2 => n191
                           , A => n4458, ZN => n4455);
   U5357 : OAI22_X1 port map( A1 => n455, A2 => n3306, B1 => n95, B2 => n3307, 
                           ZN => n4458);
   U5358 : AOI221_X1 port map( B1 => n3308, B2 => n6339, C1 => n3309, C2 => 
                           n6371, A => n4459, ZN => n4454);
   U5359 : OAI222_X1 port map( A1 => n5155, A2 => n3311, B1 => n5123, B2 => 
                           n3312, C1 => n5091, C2 => n422, ZN => n4459);
   U5360 : AOI221_X1 port map( B1 => n3313, B2 => n613, C1 => n3314, C2 => n157
                           , A => n4460, ZN => n4453);
   U5361 : OAI22_X1 port map( A1 => n61, A2 => n415, B1 => n517, B2 => n3316, 
                           ZN => n4460);
   U5362 : NAND4_X1 port map( A1 => n4461, A2 => n4462, A3 => n4463, A4 => 
                           n4464, ZN => n4442);
   U5363 : AOI221_X1 port map( B1 => n3321, B2 => n6083, C1 => n3322, C2 => 
                           n6115, A => n4465, ZN => n4464);
   U5364 : OAI222_X1 port map( A1 => n4867, A2 => n3324, B1 => n4835, B2 => 
                           n3325, C1 => n4803, C2 => n423, ZN => n4465);
   U5365 : AOI221_X1 port map( B1 => n3326, B2 => n805, C1 => n3327, C2 => n381
                           , A => n4466, ZN => n4463);
   U5366 : OAI22_X1 port map( A1 => n285, A2 => n3329, B1 => n709, B2 => n3330,
                           ZN => n4466);
   U5367 : AOI221_X1 port map( B1 => n3331, B2 => n6211, C1 => n3332, C2 => 
                           n6243, A => n4467, ZN => n4462);
   U5368 : OAI222_X1 port map( A1 => n4963, A2 => n3334, B1 => n4931, B2 => 
                           n3335, C1 => n4899, C2 => n3336, ZN => n4467);
   U5369 : AOI221_X1 port map( B1 => n3337, B2 => n614, C1 => n3338, C2 => n158
                           , A => n4468, ZN => n4461);
   U5370 : OAI22_X1 port map( A1 => n62, A2 => n3340, B1 => n518, B2 => n3341, 
                           ZN => n4468);
   U5371 : NAND4_X1 port map( A1 => n4469, A2 => n4470, A3 => n4471, A4 => 
                           n4472, ZN => n4441);
   U5372 : AOI221_X1 port map( B1 => n3346, B2 => n5827, C1 => n3347, C2 => 
                           n5859, A => n4473, ZN => n4472);
   U5373 : OAI222_X1 port map( A1 => n4611, A2 => n3349, B1 => n4579, B2 => 
                           n3350, C1 => n4547, C2 => n3351, ZN => n4473);
   U5374 : AOI221_X1 port map( B1 => n3352, B2 => n5891, C1 => n3353, C2 => 
                           n5923, A => n4474, ZN => n4471);
   U5375 : OAI22_X1 port map( A1 => n4675, A2 => n3355, B1 => n4643, B2 => 
                           n3356, ZN => n4474);
   U5376 : AOI221_X1 port map( B1 => n3357, B2 => n5955, C1 => n3358, C2 => 
                           n5987, A => n4475, ZN => n4470);
   U5377 : OAI222_X1 port map( A1 => n4771, A2 => n3360, B1 => n4739, B2 => 
                           n3361, C1 => n4707, C2 => n424, ZN => n4475);
   U5378 : AOI221_X1 port map( B1 => n3362, B2 => n6051, C1 => n3363, C2 => 
                           n6019, A => n4476, ZN => n4469);
   U5379 : OAI22_X1 port map( A1 => n5389, A2 => n3365, B1 => n5388, B2 => 
                           n3366, ZN => n4476);
   U5380 : INV_X1 port map( A => DATAIN(1), ZN => n3154);
   U5381 : OAI21_X1 port map( B1 => n3266, B2 => n1575, A => ENABLE, ZN => 
                           n7548);
   U5382 : OAI222_X1 port map( A1 => n3192, A2 => n3263, B1 => n4477, B2 => 
                           n3265, C1 => n3266, C2 => n1512, ZN => n7547);
   U5383 : NOR4_X1 port map( A1 => n4478, A2 => n4479, A3 => n4480, A4 => n4481
                           , ZN => n4477);
   U5384 : NAND4_X1 port map( A1 => n4482, A2 => n4483, A3 => n4484, A4 => 
                           n4485, ZN => n4481);
   U5385 : AOI221_X1 port map( B1 => n3275, B2 => n6402, C1 => n3276, C2 => 
                           n6434, A => n4486, ZN => n4485);
   U5386 : OAI222_X1 port map( A1 => n5250, A2 => n3278, B1 => n5218, B2 => 
                           n3279, C1 => n5186, C2 => n421, ZN => n4486);
   U5387 : AND2_X1 port map( A1 => n4490, A2 => n4493, ZN => n3275);
   U5388 : AOI221_X1 port map( B1 => n3280, B2 => n806, C1 => n3281, C2 => n382
                           , A => n4494, ZN => n4484);
   U5389 : OAI22_X1 port map( A1 => n286, A2 => n413, B1 => n710, B2 => n3283, 
                           ZN => n4494);
   U5390 : AOI221_X1 port map( B1 => n3284, B2 => n6530, C1 => n3285, C2 => 
                           n6562, A => n4498, ZN => n4483);
   U5391 : OAI222_X1 port map( A1 => n5346, A2 => n3287, B1 => n5314, B2 => 
                           n1579, C1 => n5282, C2 => n3288, ZN => n4498);
   U5392 : AND2_X1 port map( A1 => n4500, A2 => n4492, ZN => n3284);
   U5393 : AOI221_X1 port map( B1 => n3289, B2 => n807, C1 => n3290, C2 => n383
                           , A => n4501, ZN => n4482);
   U5394 : OAI22_X1 port map( A1 => n287, A2 => n414, B1 => n711, B2 => n3292, 
                           ZN => n4501);
   U5395 : NAND4_X1 port map( A1 => n4502, A2 => n4503, A3 => n4504, A4 => 
                           n4505, ZN => n4480);
   U5396 : AOI221_X1 port map( B1 => n3297, B2 => n6274, C1 => n3298, C2 => 
                           n6306, A => n4506, ZN => n4505);
   U5397 : OAI222_X1 port map( A1 => n5058, A2 => n3300, B1 => n5026, B2 => 
                           n3301, C1 => n4994, C2 => n3302, ZN => n4506);
   U5398 : AOI221_X1 port map( B1 => n3303, B2 => n552, C1 => n3304, C2 => n192
                           , A => n4509, ZN => n4504);
   U5399 : OAI22_X1 port map( A1 => n456, A2 => n3306, B1 => n96, B2 => n3307, 
                           ZN => n4509);
   U5400 : AOI221_X1 port map( B1 => n3308, B2 => n6338, C1 => n3309, C2 => 
                           n6370, A => n4510, ZN => n4503);
   U5401 : OAI222_X1 port map( A1 => n5154, A2 => n3311, B1 => n5122, B2 => 
                           n3312, C1 => n5090, C2 => n422, ZN => n4510);
   U5402 : AOI221_X1 port map( B1 => n3313, B2 => n615, C1 => n3314, C2 => n159
                           , A => n4512, ZN => n4502);
   U5403 : OAI22_X1 port map( A1 => n63, A2 => n415, B1 => n519, B2 => n3316, 
                           ZN => n4512);
   U5404 : NAND4_X1 port map( A1 => n4513, A2 => n4514, A3 => n4515, A4 => 
                           n4516, ZN => n4479);
   U5405 : AOI221_X1 port map( B1 => n3321, B2 => n6082, C1 => n3322, C2 => 
                           n6114, A => n4517, ZN => n4516);
   U5406 : OAI222_X1 port map( A1 => n4866, A2 => n3324, B1 => n4834, B2 => 
                           n3325, C1 => n4802, C2 => n423, ZN => n4517);
   U5407 : AOI221_X1 port map( B1 => n3326, B2 => n808, C1 => n3327, C2 => n384
                           , A => n4519, ZN => n4515);
   U5408 : OAI22_X1 port map( A1 => n288, A2 => n3329, B1 => n712, B2 => n3330,
                           ZN => n4519);
   U5409 : AOI221_X1 port map( B1 => n3331, B2 => n6210, C1 => n3332, C2 => 
                           n6242, A => n4521, ZN => n4514);
   U5410 : OAI222_X1 port map( A1 => n4962, A2 => n3334, B1 => n4930, B2 => 
                           n3335, C1 => n4898, C2 => n3336, ZN => n4521);
   U5411 : AOI221_X1 port map( B1 => n3337, B2 => n616, C1 => n3338, C2 => n160
                           , A => n4523, ZN => n4513);
   U5412 : OAI22_X1 port map( A1 => n64, A2 => n3340, B1 => n520, B2 => n3341, 
                           ZN => n4523);
   U5413 : NAND4_X1 port map( A1 => n4524, A2 => n4525, A3 => n4526, A4 => 
                           n4527, ZN => n4478);
   U5414 : AOI221_X1 port map( B1 => n3346, B2 => n5826, C1 => n3347, C2 => 
                           n5858, A => n4528, ZN => n4527);
   U5415 : OAI222_X1 port map( A1 => n4610, A2 => n3349, B1 => n4578, B2 => 
                           n3350, C1 => n4546, C2 => n3351, ZN => n4528);
   U5416 : AOI221_X1 port map( B1 => n3352, B2 => n5890, C1 => n3353, C2 => 
                           n5922, A => n4529, ZN => n4526);
   U5417 : OAI22_X1 port map( A1 => n4674, A2 => n3355, B1 => n4642, B2 => 
                           n3356, ZN => n4529);
   U5418 : AOI221_X1 port map( B1 => n3357, B2 => n5954, C1 => n3358, C2 => 
                           n5986, A => n4531, ZN => n4525);
   U5419 : OAI222_X1 port map( A1 => n4770, A2 => n3360, B1 => n4738, B2 => 
                           n3361, C1 => n4706, C2 => n424, ZN => n4531);
   U5420 : AND2_X1 port map( A1 => n4530, A2 => n4497, ZN => n3357);
   U5421 : AOI221_X1 port map( B1 => n3362, B2 => n6050, C1 => n3363, C2 => 
                           n6018, A => n4535, ZN => n4524);
   U5422 : OAI22_X1 port map( A1 => n5379, A2 => n3365, B1 => n5378, B2 => 
                           n3366, ZN => n4535);
   U5423 : INV_X1 port map( A => ADD_RD2(2), ZN => n4533);
   U5424 : INV_X1 port map( A => ADD_RD2(1), ZN => n4534);
   U5425 : INV_X1 port map( A => ADD_RD2(0), ZN => n4532);
   U5426 : INV_X1 port map( A => ADD_RD2(5), ZN => n4522);
   U5427 : INV_X1 port map( A => ADD_RD2(3), ZN => n4499);
   U5428 : INV_X1 port map( A => ADD_RD2(4), ZN => n4511);
   U5429 : NOR4_X1 port map( A1 => n4540, A2 => n4541, A3 => n4542, A4 => n4543
                           , ZN => n4539);
   U5430 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD2(6), Z => n4543);
   U5431 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD2(5), Z => n4542);
   U5432 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD2(4), Z => n4541);
   U5433 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD2(3), Z => n4540);
   U5434 : NOR3_X1 port map( A1 => n4544, A2 => n3261, A3 => n4545, ZN => n4538
                           );
   U5435 : INV_X1 port map( A => WR, ZN => n3261);
   U5436 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD2(0), Z => n4544);
   U5437 : XOR2_X1 port map( A => n1943, B => ADD_RD2(1), Z => n4537);
   U5438 : INV_X1 port map( A => ADD_WR(1), ZN => n1943);
   U5439 : XOR2_X1 port map( A => n1915, B => ADD_RD2(2), Z => n4536);
   U5440 : INV_X1 port map( A => ADD_WR(2), ZN => n1915);
   U5441 : INV_X1 port map( A => DATAIN(0), ZN => n3192);
   U5442 : OAI21_X1 port map( B1 => n3266, B2 => n1576, A => ENABLE, ZN => 
                           n7546);
   U5443 : INV_X1 port map( A => RD2, ZN => n4545);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5.all;

entity 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  cwp : in std_logic_vector
         (3 downto 0);  add_wr_out, add_rd1_out, add_rd2_out : out 
         std_logic_vector (6 downto 0));

end translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7;

architecture SYN_beh of 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N49, N50, N97, N98, N127, N128, r31_B_AS_3_port, r31_B_AS_4_port, 
      r31_B_AS_5_port, r31_carry_3_port, r31_carry_4_port, r31_carry_5_port, 
      r186_B_AS_3_port, r186_B_AS_4_port, r186_B_AS_5_port, r186_carry_3_port, 
      r186_carry_4_port, r186_carry_5_port, r32_B_AS_3_port, r32_B_AS_4_port, 
      r32_B_AS_5_port, r32_carry_3_port, r32_carry_4_port, r32_carry_5_port, n1
      , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17 
      : std_logic;

begin
   
   r31_U1_3 : FA_X1 port map( A => add_rd2(3), B => r31_B_AS_3_port, CI => 
                           r31_carry_3_port, CO => r31_carry_4_port, S => N127)
                           ;
   r31_U1_4 : FA_X1 port map( A => add_rd2(4), B => r31_B_AS_4_port, CI => 
                           r31_carry_4_port, CO => r31_carry_5_port, S => N128)
                           ;
   r186_U1_3 : FA_X1 port map( A => add_wr(3), B => r186_B_AS_3_port, CI => 
                           r186_carry_3_port, CO => r186_carry_4_port, S => N49
                           );
   r186_U1_4 : FA_X1 port map( A => add_wr(4), B => r186_B_AS_4_port, CI => 
                           r186_carry_4_port, CO => r186_carry_5_port, S => N50
                           );
   r32_U1_3 : FA_X1 port map( A => add_rd1(3), B => r32_B_AS_3_port, CI => 
                           r32_carry_3_port, CO => r32_carry_4_port, S => N97);
   r32_U1_4 : FA_X1 port map( A => add_rd1(4), B => r32_B_AS_4_port, CI => 
                           r32_carry_4_port, CO => r32_carry_5_port, S => N98);
   U3 : NAND2_X1 port map( A1 => r31_B_AS_5_port, A2 => r31_carry_5_port, ZN =>
                           n7);
   U4 : NAND2_X1 port map( A1 => r32_B_AS_5_port, A2 => r32_carry_5_port, ZN =>
                           n9);
   U5 : NAND2_X1 port map( A1 => r186_B_AS_5_port, A2 => r186_carry_5_port, ZN 
                           => n8);
   U6 : XNOR2_X1 port map( A => r31_carry_3_port, B => n7, ZN => n1);
   U7 : XNOR2_X1 port map( A => r32_carry_3_port, B => n9, ZN => n2);
   U8 : XNOR2_X1 port map( A => r186_carry_3_port, B => n8, ZN => n3);
   U9 : XOR2_X1 port map( A => r31_B_AS_5_port, B => r31_carry_5_port, Z => n4)
                           ;
   U10 : XOR2_X1 port map( A => r32_B_AS_5_port, B => r32_carry_5_port, Z => n5
                           );
   U11 : XOR2_X1 port map( A => r186_B_AS_5_port, B => r186_carry_5_port, Z => 
                           n6);
   U12 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => r32_B_AS_5_port);
   U13 : AND3_X1 port map( A1 => cwp(0), A2 => n12, A3 => n11, ZN => 
                           r32_B_AS_4_port);
   U14 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => r32_B_AS_3_port);
   U15 : NAND2_X1 port map( A1 => n10, A2 => n13, ZN => r31_B_AS_5_port);
   U16 : AND3_X1 port map( A1 => cwp(0), A2 => n14, A3 => n13, ZN => 
                           r31_B_AS_4_port);
   U17 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => r31_B_AS_3_port);
   U18 : NAND2_X1 port map( A1 => n10, A2 => n15, ZN => r186_B_AS_5_port);
   U19 : INV_X1 port map( A => cwp(1), ZN => n10);
   U20 : AND3_X1 port map( A1 => cwp(0), A2 => n16, A3 => n15, ZN => 
                           r186_B_AS_4_port);
   U21 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => r186_B_AS_3_port);
   U22 : AND2_X1 port map( A1 => enable, A2 => n3, ZN => add_wr_out(6));
   U23 : AND2_X1 port map( A1 => n6, A2 => enable, ZN => add_wr_out(5));
   U24 : AND2_X1 port map( A1 => N50, A2 => enable, ZN => add_wr_out(4));
   U25 : AND2_X1 port map( A1 => N49, A2 => enable, ZN => add_wr_out(3));
   U26 : AND2_X1 port map( A1 => add_wr(2), A2 => enable, ZN => add_wr_out(2));
   U27 : AND2_X1 port map( A1 => add_wr(1), A2 => enable, ZN => add_wr_out(1));
   U28 : AND2_X1 port map( A1 => add_wr(0), A2 => enable, ZN => add_wr_out(0));
   U29 : AND2_X1 port map( A1 => n1, A2 => enable, ZN => add_rd2_out(6));
   U30 : AND2_X1 port map( A1 => n4, A2 => enable, ZN => add_rd2_out(5));
   U31 : AND2_X1 port map( A1 => N128, A2 => enable, ZN => add_rd2_out(4));
   U32 : AND2_X1 port map( A1 => N127, A2 => enable, ZN => add_rd2_out(3));
   U33 : AND2_X1 port map( A1 => add_rd2(2), A2 => enable, ZN => add_rd2_out(2)
                           );
   U34 : AND2_X1 port map( A1 => add_rd2(1), A2 => enable, ZN => add_rd2_out(1)
                           );
   U35 : AND2_X1 port map( A1 => add_rd2(0), A2 => enable, ZN => add_rd2_out(0)
                           );
   U36 : AND2_X1 port map( A1 => n2, A2 => enable, ZN => add_rd1_out(6));
   U37 : AND2_X1 port map( A1 => n5, A2 => enable, ZN => add_rd1_out(5));
   U38 : AND2_X1 port map( A1 => N98, A2 => enable, ZN => add_rd1_out(4));
   U39 : AND2_X1 port map( A1 => N97, A2 => enable, ZN => add_rd1_out(3));
   U40 : AND2_X1 port map( A1 => add_rd1(2), A2 => enable, ZN => add_rd1_out(2)
                           );
   U41 : AND2_X1 port map( A1 => add_rd1(1), A2 => enable, ZN => add_rd1_out(1)
                           );
   U42 : AND2_X1 port map( A1 => add_rd1(0), A2 => enable, ZN => add_rd1_out(0)
                           );
   U43 : INV_X1 port map( A => n14, ZN => r31_carry_3_port);
   U44 : NAND3_X1 port map( A1 => n17, A2 => n13, A3 => add_rd2(4), ZN => n14);
   U45 : NAND2_X1 port map( A1 => add_rd2(3), A2 => add_rd2(4), ZN => n13);
   U46 : INV_X1 port map( A => n12, ZN => r32_carry_3_port);
   U47 : NAND3_X1 port map( A1 => add_rd1(4), A2 => n11, A3 => n17, ZN => n12);
   U48 : NAND2_X1 port map( A1 => add_rd1(4), A2 => add_rd1(3), ZN => n11);
   U49 : INV_X1 port map( A => n16, ZN => r186_carry_3_port);
   U50 : NAND3_X1 port map( A1 => n17, A2 => n15, A3 => add_wr(4), ZN => n16);
   U51 : NAND2_X1 port map( A1 => add_wr(4), A2 => add_wr(3), ZN => n15);
   U52 : AND2_X1 port map( A1 => cwp(0), A2 => cwp(1), ZN => n17);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5.all;

entity controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
         std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, spill
         : out std_logic;  MMUStrobe : in std_logic;  dataACK : out std_logic);

end controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5;

architecture SYN_beh of 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0
      port( A : in std_logic_vector (31 downto 0);  INC_DEC : in std_logic;  
            SUM : out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port, 
      swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port, 
      need_to_fill_0_port, need_to_spill_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, cansaveNext_3_port, 
      cansaveNext_2_port, cansaveNext_1_port, cansaveNext_0_port, 
      canrestoreNext_3_port, canrestoreNext_2_port, canrestoreNext_1_port, 
      canrestoreNext_0_port, actual_round_31_port, actual_round_30_port, 
      actual_round_29_port, actual_round_28_port, actual_round_27_port, 
      actual_round_26_port, actual_round_25_port, actual_round_24_port, 
      actual_round_23_port, actual_round_22_port, actual_round_21_port, 
      actual_round_20_port, actual_round_19_port, actual_round_18_port, 
      actual_round_17_port, actual_round_16_port, actual_round_15_port, 
      actual_round_14_port, actual_round_13_port, actual_round_12_port, 
      actual_round_11_port, actual_round_10_port, actual_round_9_port, 
      actual_round_8_port, actual_round_7_port, actual_round_6_port, 
      actual_round_5_port, actual_round_4_port, actual_round_3_port, 
      actual_round_2_port, actual_round_1_port, actual_round_0_port, N436, N437
      , N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
      N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, 
      N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, 
      N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, 
      N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, 
      n51, n53, n54, n63, n65, n66, n70, n71, n72, n73, n220, n221, n222, n223,
      n224, n225, n226, n227, n228, n229, n230, n234, n235, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n52, n55, n56, n57, n58, n59, n60, n61, n62, n64, n67, n68, n69, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n_2090, n_2091, n_2092 : std_logic;

begin
   cwpOut <= ( cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port );
   swpOut <= ( swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port );
   
   cansave_reg_0_inst : DFF_X1 port map( D => n230, CK => clk, Q => n1, QN => 
                           n73);
   cansaveNext_reg_2_inst : DLH_X1 port map( G => N442, D => N445, Q => 
                           cansaveNext_2_port);
   cansave_reg_2_inst : DFF_X1 port map( D => n228, CK => clk, Q => n_2090, QN 
                           => n71);
   cansaveNext_reg_3_inst : DLH_X1 port map( G => N442, D => N446, Q => 
                           cansaveNext_3_port);
   cansave_reg_3_inst : DFF_X1 port map( D => n227, CK => clk, Q => n8, QN => 
                           n70);
   nextState_reg_1_inst : DLH_X1 port map( G => N447, D => N449, Q => 
                           nextState_1_port);
   currentState_reg_1_inst : DFF_X1 port map( D => n225, CK => clk, Q => n5, QN
                           => n65);
   nextState_reg_0_inst : DLH_X1 port map( G => N447, D => N448, Q => 
                           nextState_0_port);
   currentState_reg_0_inst : DFF_X1 port map( D => n226, CK => clk, Q => n2, QN
                           => n66);
   nextState_reg_2_inst : DLH_X1 port map( G => N447, D => N450, Q => 
                           nextState_2_port);
   currentState_reg_2_inst : DFF_X1 port map( D => n224, CK => clk, Q => n_2091
                           , QN => n63);
   swp_reg_0_inst : DLH_X1 port map( G => N460, D => N461, Q => swpOut_0_port);
   swp_reg_1_inst : DLH_X1 port map( G => N460, D => N462, Q => swpOut_1_port);
   actual_round_reg_31_inst : DLH_X1 port map( G => n11, D => N497, Q => 
                           actual_round_31_port);
   actual_round_reg_0_inst : DLH_X1 port map( G => n11, D => N466, Q => 
                           actual_round_0_port);
   actual_round_reg_1_inst : DLH_X1 port map( G => n11, D => N467, Q => 
                           actual_round_1_port);
   actual_round_reg_2_inst : DLH_X1 port map( G => n11, D => N468, Q => 
                           actual_round_2_port);
   actual_round_reg_3_inst : DLH_X1 port map( G => n11, D => N469, Q => 
                           actual_round_3_port);
   actual_round_reg_4_inst : DLH_X1 port map( G => n11, D => N470, Q => 
                           actual_round_4_port);
   actual_round_reg_5_inst : DLH_X1 port map( G => n11, D => N471, Q => 
                           actual_round_5_port);
   actual_round_reg_6_inst : DLH_X1 port map( G => n11, D => N472, Q => 
                           actual_round_6_port);
   actual_round_reg_7_inst : DLH_X1 port map( G => n11, D => N473, Q => 
                           actual_round_7_port);
   actual_round_reg_8_inst : DLH_X1 port map( G => n11, D => N474, Q => 
                           actual_round_8_port);
   actual_round_reg_9_inst : DLH_X1 port map( G => n11, D => N475, Q => 
                           actual_round_9_port);
   actual_round_reg_10_inst : DLH_X1 port map( G => n11, D => N476, Q => 
                           actual_round_10_port);
   actual_round_reg_11_inst : DLH_X1 port map( G => n11, D => N477, Q => 
                           actual_round_11_port);
   actual_round_reg_12_inst : DLH_X1 port map( G => n11, D => N478, Q => 
                           actual_round_12_port);
   actual_round_reg_13_inst : DLH_X1 port map( G => n11, D => N479, Q => 
                           actual_round_13_port);
   actual_round_reg_14_inst : DLH_X1 port map( G => n11, D => N480, Q => 
                           actual_round_14_port);
   actual_round_reg_15_inst : DLH_X1 port map( G => n11, D => N481, Q => 
                           actual_round_15_port);
   actual_round_reg_16_inst : DLH_X1 port map( G => n11, D => N482, Q => 
                           actual_round_16_port);
   actual_round_reg_17_inst : DLH_X1 port map( G => n11, D => N483, Q => 
                           actual_round_17_port);
   actual_round_reg_18_inst : DLH_X1 port map( G => n11, D => N484, Q => 
                           actual_round_18_port);
   actual_round_reg_19_inst : DLH_X1 port map( G => n11, D => N485, Q => 
                           actual_round_19_port);
   actual_round_reg_20_inst : DLH_X1 port map( G => n11, D => N486, Q => 
                           actual_round_20_port);
   actual_round_reg_21_inst : DLH_X1 port map( G => n11, D => N487, Q => 
                           actual_round_21_port);
   actual_round_reg_22_inst : DLH_X1 port map( G => n11, D => N488, Q => 
                           actual_round_22_port);
   actual_round_reg_23_inst : DLH_X1 port map( G => n11, D => N489, Q => 
                           actual_round_23_port);
   actual_round_reg_24_inst : DLH_X1 port map( G => n11, D => N490, Q => 
                           actual_round_24_port);
   actual_round_reg_25_inst : DLH_X1 port map( G => n11, D => N491, Q => 
                           actual_round_25_port);
   actual_round_reg_26_inst : DLH_X1 port map( G => n11, D => N492, Q => 
                           actual_round_26_port);
   actual_round_reg_27_inst : DLH_X1 port map( G => n11, D => N493, Q => 
                           actual_round_27_port);
   actual_round_reg_28_inst : DLH_X1 port map( G => n11, D => N494, Q => 
                           actual_round_28_port);
   actual_round_reg_29_inst : DLH_X1 port map( G => n11, D => N495, Q => 
                           actual_round_29_port);
   actual_round_reg_30_inst : DLH_X1 port map( G => n11, D => N496, Q => 
                           actual_round_30_port);
   swp_reg_2_inst : DLH_X1 port map( G => N460, D => N463, Q => swpOut_2_port);
   swp_reg_3_inst : DLH_X1 port map( G => N460, D => N464, Q => swpOut_3_port);
   need_to_spill_reg_0_inst : DLH_X1 port map( G => N438, D => N439, Q => 
                           need_to_spill_0_port);
   canrestoreNext_reg_0_inst : DLH_X1 port map( G => N442, D => N451, Q => 
                           canrestoreNext_0_port);
   canrestore_reg_0_inst : DFF_X1 port map( D => n223, CK => clk, Q => n9, QN 
                           => n54);
   canrestoreNext_reg_2_inst : DLH_X1 port map( G => N442, D => N453, Q => 
                           canrestoreNext_2_port);
   canrestore_reg_2_inst : DFF_X1 port map( D => n221, CK => clk, Q => n174, QN
                           => n4);
   canrestoreNext_reg_3_inst : DLH_X1 port map( G => N442, D => N454, Q => 
                           canrestoreNext_3_port);
   canrestore_reg_3_inst : DFF_X1 port map( D => n220, CK => clk, Q => n6, QN 
                           => n51);
   need_to_fill_reg_0_inst : DLH_X1 port map( G => N436, D => N437, Q => 
                           need_to_fill_0_port);
   canrestoreNext_reg_1_inst : DLH_X1 port map( G => N442, D => N452, Q => 
                           canrestoreNext_1_port);
   canrestore_reg_1_inst : DFF_X1 port map( D => n222, CK => clk, Q => n_2092, 
                           QN => n53);
   spill_reg : DLH_X1 port map( G => N440, D => n235, Q => spill);
   fill_reg : DLH_X1 port map( G => N440, D => n234, Q => fill);
   dataACK_reg : DLH_X1 port map( G => N440, D => N441, Q => dataACK);
   cwp_reg_3_inst : DLH_X1 port map( G => N455, D => N459, Q => cwpOut_3_port);
   cwp_reg_0_inst : DLH_X1 port map( G => N455, D => N456, Q => cwpOut_0_port);
   cwp_reg_1_inst : DLH_X1 port map( G => N455, D => N457, Q => cwpOut_1_port);
   cansaveNext_reg_1_inst : DLH_X1 port map( G => N442, D => N444, Q => 
                           cansaveNext_1_port);
   cansave_reg_1_inst : DFF_X1 port map( D => n229, CK => clk, Q => n7, QN => 
                           n72);
   cansaveNext_reg_0_inst : DLH_X1 port map( G => N442, D => N443, Q => 
                           cansaveNext_0_port);
   cwp_reg_2_inst : DLH_X1 port map( G => N455, D => N458, Q => cwpOut_2_port);
   r243 : 
                           controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5_DW01_incdec_0 
                           port map( A(31) => actual_round_31_port, A(30) => 
                           actual_round_30_port, A(29) => actual_round_29_port,
                           A(28) => actual_round_28_port, A(27) => 
                           actual_round_27_port, A(26) => actual_round_26_port,
                           A(25) => actual_round_25_port, A(24) => 
                           actual_round_24_port, A(23) => actual_round_23_port,
                           A(22) => actual_round_22_port, A(21) => 
                           actual_round_21_port, A(20) => actual_round_20_port,
                           A(19) => actual_round_19_port, A(18) => 
                           actual_round_18_port, A(17) => actual_round_17_port,
                           A(16) => actual_round_16_port, A(15) => 
                           actual_round_15_port, A(14) => actual_round_14_port,
                           A(13) => actual_round_13_port, A(12) => 
                           actual_round_12_port, A(11) => actual_round_11_port,
                           A(10) => actual_round_10_port, A(9) => 
                           actual_round_9_port, A(8) => actual_round_8_port, 
                           A(7) => actual_round_7_port, A(6) => 
                           actual_round_6_port, A(5) => actual_round_5_port, 
                           A(4) => actual_round_4_port, A(3) => 
                           actual_round_3_port, A(2) => actual_round_2_port, 
                           A(1) => actual_round_1_port, A(0) => 
                           actual_round_0_port, INC_DEC => n12, SUM(31) => N497
                           , SUM(30) => N496, SUM(29) => N495, SUM(28) => N494,
                           SUM(27) => N493, SUM(26) => N492, SUM(25) => N491, 
                           SUM(24) => N490, SUM(23) => N489, SUM(22) => N488, 
                           SUM(21) => N487, SUM(20) => N486, SUM(19) => N485, 
                           SUM(18) => N484, SUM(17) => N483, SUM(16) => N482, 
                           SUM(15) => N481, SUM(14) => N480, SUM(13) => N479, 
                           SUM(12) => N478, SUM(11) => N477, SUM(10) => N476, 
                           SUM(9) => N475, SUM(8) => N474, SUM(7) => N473, 
                           SUM(6) => N472, SUM(5) => N471, SUM(4) => N470, 
                           SUM(3) => N469, SUM(2) => N468, SUM(1) => N467, 
                           SUM(0) => N466);
   U3 : OR3_X1 port map( A1 => swpOut_0_port, A2 => swpOut_1_port, A3 => n32, 
                           ZN => n3);
   U4 : INV_X1 port map( A => N465, ZN => n10);
   U5 : INV_X1 port map( A => n10, ZN => n11);
   U6 : INV_X4 port map( A => n3, ZN => n12);
   U7 : OR2_X1 port map( A1 => n13, A2 => n14, ZN => n230);
   U8 : MUX2_X1 port map( A => n1, B => cansaveNext_0_port, S => n15, Z => n14)
                           ;
   U9 : OR2_X1 port map( A1 => n13, A2 => n16, ZN => n229);
   U10 : MUX2_X1 port map( A => n7, B => cansaveNext_1_port, S => n15, Z => n16
                           );
   U11 : OAI21_X1 port map( B1 => n71, B2 => n15, A => n17, ZN => n228);
   U12 : NAND2_X1 port map( A1 => cansaveNext_2_port, A2 => n18, ZN => n17);
   U13 : OAI21_X1 port map( B1 => n70, B2 => n15, A => n19, ZN => n227);
   U14 : NAND2_X1 port map( A1 => cansaveNext_3_port, A2 => n18, ZN => n19);
   U15 : OR2_X1 port map( A1 => n13, A2 => n20, ZN => n226);
   U16 : MUX2_X1 port map( A => n2, B => nextState_0_port, S => n15, Z => n20);
   U17 : NOR2_X1 port map( A1 => n21, A2 => n18, ZN => n13);
   U18 : OAI21_X1 port map( B1 => n65, B2 => n15, A => n22, ZN => n225);
   U19 : NAND2_X1 port map( A1 => nextState_1_port, A2 => n18, ZN => n22);
   U20 : OAI21_X1 port map( B1 => n63, B2 => n15, A => n23, ZN => n224);
   U21 : NAND2_X1 port map( A1 => nextState_2_port, A2 => n18, ZN => n23);
   U22 : OAI21_X1 port map( B1 => n54, B2 => n15, A => n24, ZN => n223);
   U23 : NAND2_X1 port map( A1 => canrestoreNext_0_port, A2 => n18, ZN => n24);
   U24 : OAI21_X1 port map( B1 => n53, B2 => n15, A => n25, ZN => n222);
   U25 : NAND2_X1 port map( A1 => canrestoreNext_1_port, A2 => n18, ZN => n25);
   U26 : OAI21_X1 port map( B1 => n15, B2 => n4, A => n26, ZN => n221);
   U27 : NAND2_X1 port map( A1 => canrestoreNext_2_port, A2 => n18, ZN => n26);
   U28 : OAI21_X1 port map( B1 => n51, B2 => n15, A => n27, ZN => n220);
   U29 : NAND2_X1 port map( A1 => canrestoreNext_3_port, A2 => n18, ZN => n27);
   U30 : INV_X1 port map( A => n21, ZN => n15);
   U31 : NOR2_X1 port map( A1 => reset, A2 => n18, ZN => n21);
   U32 : NOR2_X1 port map( A1 => n28, A2 => reset, ZN => n18);
   U33 : INV_X1 port map( A => enable, ZN => n28);
   U34 : AOI21_X1 port map( B1 => n3, B2 => n29, A => n30, ZN => N465);
   U35 : NAND2_X1 port map( A1 => n235, A2 => n31, ZN => n29);
   U36 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => N464);
   U37 : XOR2_X1 port map( A => n35, B => n36, Z => n33);
   U38 : AOI22_X1 port map( A1 => n37, A2 => n235, B1 => swpOut_3_port, B2 => 
                           n234, ZN => n35);
   U39 : MUX2_X1 port map( A => n38, B => n39, S => n31, Z => n37);
   U40 : XNOR2_X1 port map( A => N467, B => n40, ZN => n39);
   U41 : XNOR2_X1 port map( A => actual_round_1_port, B => n40, ZN => n38);
   U42 : OAI221_X1 port map( B1 => n41, B2 => n42, C1 => n234, C2 => n41, A => 
                           n43, ZN => N463);
   U43 : NOR2_X1 port map( A1 => n44, A2 => n36, ZN => n43);
   U44 : AND3_X1 port map( A1 => n234, A2 => n41, A3 => n42, ZN => n36);
   U45 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => n42);
   U46 : AOI22_X1 port map( A1 => n234, A2 => swpOut_2_port, B1 => n47, B2 => 
                           n235, ZN => n41);
   U47 : INV_X1 port map( A => n40, ZN => n47);
   U48 : MUX2_X1 port map( A => actual_round_0_port, B => N466, S => n31, Z => 
                           n40);
   U49 : AND2_X1 port map( A1 => swpOut_1_port, A2 => swpOut_0_port, ZN => n31)
                           ;
   U50 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n34, ZN => N462);
   U51 : XOR2_X1 port map( A => n46, B => n45, Z => n49);
   U52 : AND2_X1 port map( A1 => swpOut_0_port, A2 => n234, ZN => n45);
   U53 : AND2_X1 port map( A1 => swpOut_1_port, A2 => n234, ZN => n46);
   U54 : AOI21_X1 port map( B1 => n235, B2 => n50, A => n234, ZN => n48);
   U55 : XOR2_X1 port map( A => swpOut_1_port, B => swpOut_0_port, Z => n50);
   U56 : OAI21_X1 port map( B1 => swpOut_0_port, B2 => n52, A => n34, ZN => 
                           N461);
   U57 : NAND2_X1 port map( A1 => n55, A2 => n34, ZN => N460);
   U58 : NOR2_X1 port map( A1 => n56, A2 => n57, ZN => N459);
   U59 : NOR2_X1 port map( A1 => n56, A2 => n58, ZN => N458);
   U60 : NOR2_X1 port map( A1 => n56, A2 => n59, ZN => N457);
   U61 : NOR2_X1 port map( A1 => n56, A2 => n60, ZN => N456);
   U62 : OR2_X1 port map( A1 => n61, A2 => n44, ZN => N455);
   U63 : OAI21_X1 port map( B1 => n62, B2 => n64, A => n67, ZN => N454);
   U64 : MUX2_X1 port map( A => n68, B => n69, S => n6, Z => n67);
   U65 : AOI21_X1 port map( B1 => n74, B2 => n4, A => n75, ZN => n69);
   U66 : INV_X1 port map( A => n76, ZN => n75);
   U67 : NAND3_X1 port map( A1 => n74, A2 => n174, A3 => n77, ZN => n68);
   U68 : XOR2_X1 port map( A => n78, B => n79, Z => n64);
   U69 : XNOR2_X1 port map( A => n51, B => n80, ZN => n79);
   U70 : AOI21_X1 port map( B1 => n81, B2 => n80, A => n82, ZN => n78);
   U71 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n4, ZN => n82);
   U72 : INV_X1 port map( A => n84, ZN => n81);
   U73 : OAI21_X1 port map( B1 => n62, B2 => n85, A => n86, ZN => N453);
   U74 : MUX2_X1 port map( A => n76, B => n87, S => n4, Z => n86);
   U75 : NAND2_X1 port map( A1 => n77, A2 => n74, ZN => n87);
   U76 : NAND2_X1 port map( A1 => n74, A2 => n88, ZN => n76);
   U77 : XNOR2_X1 port map( A => n84, B => n89, ZN => n85);
   U78 : XNOR2_X1 port map( A => n174, B => n80, ZN => n89);
   U79 : AOI21_X1 port map( B1 => n80, B2 => n90, A => n77, ZN => n84);
   U80 : OAI22_X1 port map( A1 => n91, A2 => n92, B1 => n62, B2 => n93, ZN => 
                           N452);
   U81 : XNOR2_X1 port map( A => n83, B => n92, ZN => n93);
   U82 : INV_X1 port map( A => n80, ZN => n83);
   U83 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n80);
   U84 : AND2_X1 port map( A1 => n97, A2 => n98, ZN => n62);
   U85 : NAND2_X1 port map( A1 => n90, A2 => n88, ZN => n92);
   U86 : INV_X1 port map( A => n77, ZN => n88);
   U87 : NOR2_X1 port map( A1 => n53, A2 => n54, ZN => n77);
   U88 : AOI21_X1 port map( B1 => n97, B2 => n99, A => n9, ZN => N451);
   U89 : OAI221_X1 port map( B1 => n100, B2 => n101, C1 => n102, C2 => n103, A 
                           => n104, ZN => N450);
   U90 : AOI222_X1 port map( A1 => n105, A2 => n30, B1 => n106, B2 => n107, C1 
                           => n108, C2 => n109, ZN => n104);
   U91 : OAI211_X1 port map( C1 => n110, C2 => n111, A => n112, B => n113, ZN 
                           => N449);
   U92 : NAND3_X1 port map( A1 => n114, A2 => n101, A3 => n115, ZN => n112);
   U93 : INV_X1 port map( A => n116, ZN => n101);
   U94 : INV_X1 port map( A => n108, ZN => n111);
   U95 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN 
                           => N448);
   U96 : AOI22_X1 port map( A1 => reset, A2 => n44, B1 => n234, B2 => n30, ZN 
                           => n120);
   U97 : OAI21_X1 port map( B1 => n121, B2 => n116, A => n114, ZN => n119);
   U98 : NAND3_X1 port map( A1 => n122, A2 => n123, A3 => n102, ZN => n117);
   U99 : NAND4_X1 port map( A1 => n56, A2 => call, A3 => n124, A4 => n65, ZN =>
                           N447);
   U100 : NOR2_X1 port map( A1 => n44, A2 => n115, ZN => n124);
   U101 : INV_X1 port map( A => n125, ZN => n115);
   U102 : INV_X1 port map( A => n34, ZN => n44);
   U103 : OAI22_X1 port map( A1 => n98, A2 => n57, B1 => n126, B2 => n127, ZN 
                           => N446);
   U104 : XOR2_X1 port map( A => n128, B => n129, Z => n127);
   U105 : XNOR2_X1 port map( A => n70, B => n130, ZN => n129);
   U106 : OAI21_X1 port map( B1 => n131, B2 => n130, A => n132, ZN => n128);
   U107 : OAI21_X1 port map( B1 => n133, B2 => n134, A => n71, ZN => n132);
   U108 : XOR2_X1 port map( A => n135, B => n136, Z => n57);
   U109 : XNOR2_X1 port map( A => n137, B => n138, ZN => n136);
   U110 : AOI22_X1 port map( A1 => cwpOut_3_port, A2 => n61, B1 => n139, B2 => 
                           n8, ZN => n137);
   U111 : AOI21_X1 port map( B1 => n140, B2 => n141, A => n142, ZN => n135);
   U112 : INV_X1 port map( A => n143, ZN => n142);
   U113 : OAI21_X1 port map( B1 => n141, B2 => n140, A => n138, ZN => n143);
   U114 : OAI22_X1 port map( A1 => n58, A2 => n98, B1 => n126, B2 => n144, ZN 
                           => N445);
   U115 : XNOR2_X1 port map( A => n133, B => n145, ZN => n144);
   U116 : XNOR2_X1 port map( A => n134, B => n71, ZN => n145);
   U117 : INV_X1 port map( A => n131, ZN => n133);
   U118 : OAI22_X1 port map( A1 => n73, A2 => n72, B1 => n146, B2 => n134, ZN 
                           => n131);
   U119 : XOR2_X1 port map( A => n147, B => n141, Z => n58);
   U120 : AOI21_X1 port map( B1 => n148, B2 => n149, A => n150, ZN => n141);
   U121 : AOI21_X1 port map( B1 => n138, B2 => n151, A => n60, ZN => n150);
   U122 : INV_X1 port map( A => n138, ZN => n149);
   U123 : XNOR2_X1 port map( A => n140, B => n138, ZN => n147);
   U124 : OAI21_X1 port map( B1 => n71, B2 => n98, A => n152, ZN => n140);
   U125 : NAND2_X1 port map( A1 => cwpOut_2_port, A2 => n61, ZN => n152);
   U126 : OAI221_X1 port map( B1 => n126, B2 => n153, C1 => n98, C2 => n59, A 
                           => n34, ZN => N444);
   U127 : XNOR2_X1 port map( A => n154, B => n148, ZN => n59);
   U128 : INV_X1 port map( A => n151, ZN => n148);
   U129 : OAI21_X1 port map( B1 => n72, B2 => n98, A => n155, ZN => n151);
   U130 : NAND2_X1 port map( A1 => cwpOut_1_port, A2 => n61, ZN => n155);
   U131 : XNOR2_X1 port map( A => n60, B => n138, ZN => n154);
   U132 : OAI21_X1 port map( B1 => n32, B2 => n30, A => n156, ZN => n138);
   U133 : AOI21_X1 port map( B1 => n146, B2 => n130, A => n157, ZN => n153);
   U134 : MUX2_X1 port map( A => n158, B => n159, S => n1, Z => n157);
   U135 : XNOR2_X1 port map( A => n134, B => n72, ZN => n159);
   U136 : INV_X1 port map( A => n130, ZN => n134);
   U137 : NOR2_X1 port map( A1 => n72, A2 => n130, ZN => n158);
   U138 : NAND2_X1 port map( A1 => n160, A2 => n161, ZN => n130);
   U139 : OAI221_X1 port map( B1 => n98, B2 => n60, C1 => n126, C2 => n1, A => 
                           n34, ZN => N443);
   U140 : AND2_X1 port map( A1 => n97, A2 => n91, ZN => n126);
   U141 : INV_X1 port map( A => n74, ZN => n91);
   U142 : AOI21_X1 port map( B1 => n162, B2 => n122, A => n99, ZN => n74);
   U143 : OAI21_X1 port map( B1 => n73, B2 => n98, A => n163, ZN => n60);
   U144 : NAND2_X1 port map( A1 => cwpOut_0_port, A2 => n61, ZN => n163);
   U145 : NAND3_X1 port map( A1 => n161, A2 => n55, A3 => n156, ZN => n61);
   U146 : NAND3_X1 port map( A1 => n164, A2 => n162, A3 => n114, ZN => n156);
   U147 : INV_X1 port map( A => N441, ZN => n55);
   U148 : INV_X1 port map( A => n139, ZN => n98);
   U149 : NAND3_X1 port map( A1 => n34, A2 => n160, A3 => n113, ZN => N442);
   U150 : NOR2_X1 port map( A1 => n165, A2 => n166, ZN => n113);
   U151 : AOI21_X1 port map( B1 => n94, B2 => n110, A => n95, ZN => n166);
   U152 : NAND2_X1 port map( A1 => n102, A2 => n167, ZN => n95);
   U153 : AND2_X1 port map( A1 => n168, A2 => n169, ZN => n102);
   U154 : NAND2_X1 port map( A1 => need_to_spill_0_port, A2 => n110, ZN => n169
                           );
   U155 : INV_X1 port map( A => n96, ZN => n165);
   U156 : AOI21_X1 port map( B1 => n114, B2 => n121, A => n139, ZN => n96);
   U157 : NOR2_X1 port map( A1 => n118, A2 => n106, ZN => n139);
   U158 : INV_X1 port map( A => n107, ZN => n118);
   U159 : NOR2_X1 port map( A1 => n99, A2 => n94, ZN => n107);
   U160 : INV_X1 port map( A => n122, ZN => n94);
   U161 : NOR2_X1 port map( A1 => n170, A2 => call, ZN => n122);
   U162 : NOR2_X1 port map( A1 => n170, A2 => n116, ZN => n121);
   U163 : MUX2_X1 port map( A => n106, B => need_to_fill_0_port, S => n171, Z 
                           => n116);
   U164 : NAND2_X1 port map( A1 => n108, A2 => n168, ZN => n160);
   U165 : NOR2_X1 port map( A1 => n125, A2 => n99, ZN => n108);
   U166 : NAND2_X1 port map( A1 => call, A2 => n170, ZN => n125);
   U167 : NOR2_X1 port map( A1 => n30, A2 => n52, ZN => N441);
   U168 : INV_X1 port map( A => MMUStrobe, ZN => n30);
   U169 : NAND3_X1 port map( A1 => n34, A2 => n99, A3 => n56, ZN => N440);
   U170 : AND2_X1 port map( A1 => n97, A2 => n52, ZN => n56);
   U171 : NOR2_X1 port map( A1 => n235, A2 => n234, ZN => n52);
   U172 : INV_X1 port map( A => n32, ZN => n234);
   U173 : INV_X1 port map( A => n172, ZN => n235);
   U174 : NOR2_X1 port map( A1 => n167, A2 => n114, ZN => n97);
   U175 : INV_X1 port map( A => n100, ZN => n114);
   U176 : INV_X1 port map( A => n103, ZN => n167);
   U177 : NAND3_X1 port map( A1 => n65, A2 => n2, A3 => n63, ZN => n34);
   U178 : NAND4_X1 port map( A1 => n161, A2 => n99, A3 => n173, A4 => n172, ZN 
                           => N438);
   U179 : NAND2_X1 port map( A1 => n66, A2 => n105, ZN => n172);
   U180 : INV_X1 port map( A => N439, ZN => n173);
   U181 : NOR2_X1 port map( A1 => n168, A2 => n103, ZN => N439);
   U182 : OR2_X1 port map( A1 => n103, A2 => n110, ZN => n161);
   U183 : NAND2_X1 port map( A1 => call, A2 => n168, ZN => n110);
   U184 : NAND2_X1 port map( A1 => n123, A2 => n5, ZN => n103);
   U185 : NOR2_X1 port map( A1 => n100, A2 => n162, ZN => N437);
   U186 : INV_X1 port map( A => n106, ZN => n162);
   U187 : OAI211_X1 port map( C1 => n171, C2 => n100, A => n99, B => n32, ZN =>
                           N436);
   U188 : NAND2_X1 port map( A1 => n105, A2 => n2, ZN => n32);
   U189 : NOR2_X1 port map( A1 => n5, A2 => n63, ZN => n105);
   U190 : NAND2_X1 port map( A1 => n123, A2 => n65, ZN => n99);
   U191 : AND2_X1 port map( A1 => n63, A2 => n66, ZN => n123);
   U192 : NAND3_X1 port map( A1 => n5, A2 => n2, A3 => n63, ZN => n100);
   U193 : NOR2_X1 port map( A1 => n164, A2 => n106, ZN => n171);
   U194 : NOR3_X1 port map( A1 => n90, A2 => n174, A3 => n6, ZN => n106);
   U195 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => n90);
   U196 : NOR2_X1 port map( A1 => n170, A2 => n109, ZN => n164);
   U197 : INV_X1 port map( A => n168, ZN => n109);
   U198 : NAND3_X1 port map( A1 => n70, A2 => n146, A3 => n71, ZN => n168);
   U199 : NOR2_X1 port map( A1 => n1, A2 => n7, ZN => n146);
   U200 : INV_X1 port map( A => ret, ZN => n170);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use 
   work.CONV_PACK_registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5.all;

entity registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5 is

   port( clk, reset, enable, rd1, rd2, wr1 : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  dataIn : in 
         std_logic_vector (31 downto 0);  dataOut1, dataOut2 : out 
         std_logic_vector (31 downto 0);  fill, spill : out std_logic;  call, 
         ret : in std_logic;  dataACK : out std_logic;  MMUStrobe : in 
         std_logic);

end registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5;

architecture SYN_struct of 
   registerFile_TLE_N8_M8_windowBlocks3_NData32_NAddr_Windowed5 is

   component physical_RF_NData32_NRegs72_NAddr7
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (6 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7
      port( clk, reset, enable, rd1, rd2, wr : in std_logic;  add_wr, add_rd1, 
            add_rd2 : in std_logic_vector (4 downto 0);  cwp : in 
            std_logic_vector (3 downto 0);  add_wr_out, add_rd1_out, 
            add_rd2_out : out std_logic_vector (6 downto 0));
   end component;
   
   component controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5
      port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
            std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, 
            spill : out std_logic;  MMUStrobe : in std_logic;  dataACK : out 
            std_logic);
   end component;
   
   signal cwp_s_3_port, cwp_s_2_port, cwp_s_1_port, cwp_s_0_port, 
      add_wr_out_s_6_port, add_wr_out_s_5_port, add_wr_out_s_4_port, 
      add_wr_out_s_3_port, add_wr_out_s_2_port, add_wr_out_s_1_port, 
      add_wr_out_s_0_port, add_rd1_out_s_6_port, add_rd1_out_s_5_port, 
      add_rd1_out_s_4_port, add_rd1_out_s_3_port, add_rd1_out_s_2_port, 
      add_rd1_out_s_1_port, add_rd1_out_s_0_port, add_rd2_out_s_6_port, 
      add_rd2_out_s_5_port, add_rd2_out_s_4_port, add_rd2_out_s_3_port, 
      add_rd2_out_s_2_port, add_rd2_out_s_1_port, add_rd2_out_s_0_port, n_2093,
      n_2094, n_2095, n_2096 : std_logic;

begin
   
   contrU : controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 port 
                           map( clk => clk, reset => reset, enable => enable, 
                           cwpOut(3) => cwp_s_3_port, cwpOut(2) => cwp_s_2_port
                           , cwpOut(1) => cwp_s_1_port, cwpOut(0) => 
                           cwp_s_0_port, swpOut(3) => n_2093, swpOut(2) => 
                           n_2094, swpOut(1) => n_2095, swpOut(0) => n_2096, 
                           call => call, ret => ret, fill => fill, spill => 
                           spill, MMUStrobe => MMUStrobe, dataACK => dataACK);
   translU : 
                           translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 
                           port map( clk => clk, reset => reset, enable => 
                           enable, rd1 => rd1, rd2 => rd2, wr => wr1, add_wr(4)
                           => add_wr(4), add_wr(3) => add_wr(3), add_wr(2) => 
                           add_wr(2), add_wr(1) => add_wr(1), add_wr(0) => 
                           add_wr(0), add_rd1(4) => add_rd1(4), add_rd1(3) => 
                           add_rd1(3), add_rd1(2) => add_rd1(2), add_rd1(1) => 
                           add_rd1(1), add_rd1(0) => add_rd1(0), add_rd2(4) => 
                           add_rd2(4), add_rd2(3) => add_rd2(3), add_rd2(2) => 
                           add_rd2(2), add_rd2(1) => add_rd2(1), add_rd2(0) => 
                           add_rd2(0), cwp(3) => cwp_s_3_port, cwp(2) => 
                           cwp_s_2_port, cwp(1) => cwp_s_1_port, cwp(0) => 
                           cwp_s_0_port, add_wr_out(6) => add_wr_out_s_6_port, 
                           add_wr_out(5) => add_wr_out_s_5_port, add_wr_out(4) 
                           => add_wr_out_s_4_port, add_wr_out(3) => 
                           add_wr_out_s_3_port, add_wr_out(2) => 
                           add_wr_out_s_2_port, add_wr_out(1) => 
                           add_wr_out_s_1_port, add_wr_out(0) => 
                           add_wr_out_s_0_port, add_rd1_out(6) => 
                           add_rd1_out_s_6_port, add_rd1_out(5) => 
                           add_rd1_out_s_5_port, add_rd1_out(4) => 
                           add_rd1_out_s_4_port, add_rd1_out(3) => 
                           add_rd1_out_s_3_port, add_rd1_out(2) => 
                           add_rd1_out_s_2_port, add_rd1_out(1) => 
                           add_rd1_out_s_1_port, add_rd1_out(0) => 
                           add_rd1_out_s_0_port, add_rd2_out(6) => 
                           add_rd2_out_s_6_port, add_rd2_out(5) => 
                           add_rd2_out_s_5_port, add_rd2_out(4) => 
                           add_rd2_out_s_4_port, add_rd2_out(3) => 
                           add_rd2_out_s_3_port, add_rd2_out(2) => 
                           add_rd2_out_s_2_port, add_rd2_out(1) => 
                           add_rd2_out_s_1_port, add_rd2_out(0) => 
                           add_rd2_out_s_0_port);
   physRF : physical_RF_NData32_NRegs72_NAddr7 port map( CLK => clk, RESET => 
                           reset, ENABLE => enable, RD1 => rd1, RD2 => rd2, WR 
                           => wr1, ADD_WR(6) => add_wr_out_s_6_port, ADD_WR(5) 
                           => add_wr_out_s_5_port, ADD_WR(4) => 
                           add_wr_out_s_4_port, ADD_WR(3) => 
                           add_wr_out_s_3_port, ADD_WR(2) => 
                           add_wr_out_s_2_port, ADD_WR(1) => 
                           add_wr_out_s_1_port, ADD_WR(0) => 
                           add_wr_out_s_0_port, ADD_RD1(6) => 
                           add_rd1_out_s_6_port, ADD_RD1(5) => 
                           add_rd1_out_s_5_port, ADD_RD1(4) => 
                           add_rd1_out_s_4_port, ADD_RD1(3) => 
                           add_rd1_out_s_3_port, ADD_RD1(2) => 
                           add_rd1_out_s_2_port, ADD_RD1(1) => 
                           add_rd1_out_s_1_port, ADD_RD1(0) => 
                           add_rd1_out_s_0_port, ADD_RD2(6) => 
                           add_rd2_out_s_6_port, ADD_RD2(5) => 
                           add_rd2_out_s_5_port, ADD_RD2(4) => 
                           add_rd2_out_s_4_port, ADD_RD2(3) => 
                           add_rd2_out_s_3_port, ADD_RD2(2) => 
                           add_rd2_out_s_2_port, ADD_RD2(1) => 
                           add_rd2_out_s_1_port, ADD_RD2(0) => 
                           add_rd2_out_s_0_port, DATAIN(31) => dataIn(31), 
                           DATAIN(30) => dataIn(30), DATAIN(29) => dataIn(29), 
                           DATAIN(28) => dataIn(28), DATAIN(27) => dataIn(27), 
                           DATAIN(26) => dataIn(26), DATAIN(25) => dataIn(25), 
                           DATAIN(24) => dataIn(24), DATAIN(23) => dataIn(23), 
                           DATAIN(22) => dataIn(22), DATAIN(21) => dataIn(21), 
                           DATAIN(20) => dataIn(20), DATAIN(19) => dataIn(19), 
                           DATAIN(18) => dataIn(18), DATAIN(17) => dataIn(17), 
                           DATAIN(16) => dataIn(16), DATAIN(15) => dataIn(15), 
                           DATAIN(14) => dataIn(14), DATAIN(13) => dataIn(13), 
                           DATAIN(12) => dataIn(12), DATAIN(11) => dataIn(11), 
                           DATAIN(10) => dataIn(10), DATAIN(9) => dataIn(9), 
                           DATAIN(8) => dataIn(8), DATAIN(7) => dataIn(7), 
                           DATAIN(6) => dataIn(6), DATAIN(5) => dataIn(5), 
                           DATAIN(4) => dataIn(4), DATAIN(3) => dataIn(3), 
                           DATAIN(2) => dataIn(2), DATAIN(1) => dataIn(1), 
                           DATAIN(0) => dataIn(0), OUT1(31) => dataOut1(31), 
                           OUT1(30) => dataOut1(30), OUT1(29) => dataOut1(29), 
                           OUT1(28) => dataOut1(28), OUT1(27) => dataOut1(27), 
                           OUT1(26) => dataOut1(26), OUT1(25) => dataOut1(25), 
                           OUT1(24) => dataOut1(24), OUT1(23) => dataOut1(23), 
                           OUT1(22) => dataOut1(22), OUT1(21) => dataOut1(21), 
                           OUT1(20) => dataOut1(20), OUT1(19) => dataOut1(19), 
                           OUT1(18) => dataOut1(18), OUT1(17) => dataOut1(17), 
                           OUT1(16) => dataOut1(16), OUT1(15) => dataOut1(15), 
                           OUT1(14) => dataOut1(14), OUT1(13) => dataOut1(13), 
                           OUT1(12) => dataOut1(12), OUT1(11) => dataOut1(11), 
                           OUT1(10) => dataOut1(10), OUT1(9) => dataOut1(9), 
                           OUT1(8) => dataOut1(8), OUT1(7) => dataOut1(7), 
                           OUT1(6) => dataOut1(6), OUT1(5) => dataOut1(5), 
                           OUT1(4) => dataOut1(4), OUT1(3) => dataOut1(3), 
                           OUT1(2) => dataOut1(2), OUT1(1) => dataOut1(1), 
                           OUT1(0) => dataOut1(0), OUT2(31) => dataOut2(31), 
                           OUT2(30) => dataOut2(30), OUT2(29) => dataOut2(29), 
                           OUT2(28) => dataOut2(28), OUT2(27) => dataOut2(27), 
                           OUT2(26) => dataOut2(26), OUT2(25) => dataOut2(25), 
                           OUT2(24) => dataOut2(24), OUT2(23) => dataOut2(23), 
                           OUT2(22) => dataOut2(22), OUT2(21) => dataOut2(21), 
                           OUT2(20) => dataOut2(20), OUT2(19) => dataOut2(19), 
                           OUT2(18) => dataOut2(18), OUT2(17) => dataOut2(17), 
                           OUT2(16) => dataOut2(16), OUT2(15) => dataOut2(15), 
                           OUT2(14) => dataOut2(14), OUT2(13) => dataOut2(13), 
                           OUT2(12) => dataOut2(12), OUT2(11) => dataOut2(11), 
                           OUT2(10) => dataOut2(10), OUT2(9) => dataOut2(9), 
                           OUT2(8) => dataOut2(8), OUT2(7) => dataOut2(7), 
                           OUT2(6) => dataOut2(6), OUT2(5) => dataOut2(5), 
                           OUT2(4) => dataOut2(4), OUT2(3) => dataOut2(3), 
                           OUT2(2) => dataOut2(2), OUT2(1) => dataOut2(1), 
                           OUT2(0) => dataOut2(0));

end SYN_struct;
