
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerFile_TLE is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerFile_TLE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity physical_RF_NData32_NRegs72_NAddr7 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR, RD_Mem, WR_Mem : in std_logic;  
         ADD_WR, ADD_RD1, ADD_RD2, ADD_SF : in std_logic_vector (6 downto 0);  
         DATAIN : in std_logic_vector (31 downto 0);  OUT1, OUT2, RFtoMEM_BUS :
         out std_logic_vector (31 downto 0));

end physical_RF_NData32_NRegs72_NAddr7;

architecture SYN_beh of physical_RF_NData32_NRegs72_NAddr7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9102, n9103, n9104, n9105, n9106, n9107, 
      n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
      n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, 
      n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, 
      n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, 
      n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, 
      n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
      n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, 
      n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
      n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, 
      n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, 
      n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, 
      n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, 
      n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, 
      n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, 
      n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, 
      n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, 
      n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, 
      n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, 
      n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, 
      n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, 
      n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, 
      n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, 
      n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, 
      n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, 
      n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, 
      n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, 
      n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, 
      n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, 
      n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, 
      n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
      n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, 
      n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, 
      n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, 
      n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, 
      n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, 
      n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, 
      n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, 
      n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, 
      n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, 
      n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, 
      n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, 
      n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, 
      n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, 
      n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, 
      n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, 
      n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, 
      n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, 
      n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, 
      n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, 
      n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, 
      n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, 
      n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, 
      n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, 
      n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, 
      n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, 
      n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, 
      n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, 
      n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, 
      n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, 
      n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, 
      n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, 
      n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, 
      n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, 
      n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, 
      n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, 
      n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
      n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, 
      n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, 
      n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, 
      n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, 
      n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, 
      n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, 
      n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, 
      n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
      n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, 
      n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, 
      n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, 
      n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
      n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, 
      n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, 
      n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, 
      n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
      n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, 
      n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, 
      n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, 
      n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, 
      n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, 
      n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, 
      n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
      n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, 
      n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, 
      n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
      n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, 
      n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, 
      n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
      n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, 
      n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, 
      n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, 
      n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
      n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, 
      n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, 
      n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, 
      n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, 
      n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, 
      n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, 
      n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, 
      n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, 
      n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, 
      n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, 
      n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, 
      n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, 
      n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, 
      n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, 
      n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, 
      n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
      n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, 
      n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, 
      n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, 
      n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, 
      n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, 
      n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, 
      n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, 
      n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, 
      n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, 
      n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
      n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, 
      n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, 
      n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, 
      n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, 
      n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, 
      n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, 
      n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, 
      n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, 
      n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, 
      n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, 
      n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, 
      n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, 
      n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, 
      n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, 
      n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, 
      n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, 
      n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, 
      n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, 
      n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, 
      n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, 
      n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, 
      n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, 
      n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, 
      n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, 
      n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, 
      n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, 
      n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, 
      n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, 
      n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, 
      n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, 
      n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, 
      n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, 
      n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, 
      n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, 
      n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, 
      n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, 
      n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, 
      n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, 
      n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, 
      n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, 
      n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, 
      n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, 
      n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, 
      n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, 
      n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, 
      n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, 
      n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, 
      n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, 
      n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, 
      n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, 
      n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, 
      n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
      n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, 
      n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, 
      n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, 
      n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, 
      n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
      n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, 
      n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
      n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, 
      n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, 
      n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, 
      n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, 
      n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, 
      n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
      n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, 
      n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, 
      n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, 
      n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, 
      n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, 
      n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, 
      n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, 
      n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, 
      n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, 
      n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, 
      n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, 
      n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, 
      n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, 
      n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, 
      n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, 
      n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, 
      n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, 
      n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, 
      n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, 
      n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, 
      n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, 
      n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, 
      n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, 
      n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, 
      n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, 
      n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, 
      n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, 
      n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, 
      n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, 
      n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, 
      n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, 
      n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, 
      n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, 
      n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, 
      n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, 
      n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, 
      n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, 
      n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, 
      n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, 
      n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, 
      n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, 
      n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, 
      n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, 
      n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, 
      n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, 
      n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, 
      n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, 
      n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, 
      n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
      n11501, n76, n82, n88, n94, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n899, n905, n911, n917, n923, n929, n935, n941, n947, n953, n959, 
      n965, n971, n977, n983, n989, n995, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, 
      n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
      n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
      n2275, n2276, n2277, n6726, n6727, n6728, n6731, n6734, n6737, n6740, 
      n6741, n6742, n6743, n6744, n6745, n6746, n6750, n6752, n6755, n6756, 
      n6758, n6761, n6762, n6764, n6765, n6766, n6767, n6768, n6770, n6774, 
      n6776, n6779, n6782, n6785, n6786, n6788, n6789, n6790, n6791, n6792, 
      n6794, n6798, n6800, n6803, n6804, n6806, n6809, n6810, n6812, n6813, 
      n6814, n6815, n6816, n6818, n6822, n6824, n6827, n6828, n6830, n6833, 
      n6834, n6836, n6837, n6838, n6839, n6840, n6842, n6846, n6848, n6851, 
      n6852, n6854, n6857, n6858, n6860, n6861, n6862, n6863, n6864, n6866, 
      n6870, n6872, n6875, n6876, n6878, n6881, n6882, n6884, n6885, n6886, 
      n6887, n6888, n6890, n6894, n6896, n6899, n6900, n6902, n6905, n6906, 
      n6908, n6909, n6910, n6911, n6912, n6914, n6918, n6920, n6923, n6924, 
      n6926, n6929, n6930, n6932, n6933, n6934, n6935, n6936, n6938, n6942, 
      n6944, n6947, n6948, n6950, n6953, n6954, n6956, n6957, n6958, n6959, 
      n6960, n6962, n6966, n6968, n6971, n6972, n6974, n6977, n6978, n6980, 
      n6981, n6982, n6983, n6984, n6986, n6990, n6992, n6995, n6996, n6998, 
      n7001, n7002, n7004, n7005, n7006, n7007, n7008, n7010, n7014, n7016, 
      n7019, n7020, n7022, n7025, n7028, n7029, n7030, n7031, n7034, n7038, 
      n7040, n7043, n7046, n7049, n7052, n7054, n7055, n7058, n7062, n7064, 
      n7067, n7070, n7073, n7076, n7078, n7079, n7082, n7086, n7088, n7091, 
      n7094, n7097, n7100, n7102, n7103, n7106, n7110, n7112, n7115, n7118, 
      n7121, n7124, n7126, n7127, n7130, n7134, n7136, n7139, n7142, n7145, 
      n7146, n7148, n7149, n7150, n7151, n7152, n7154, n7158, n7159, n7160, 
      n7163, n7166, n7169, n7172, n7173, n7174, n7175, n7176, n7177, n7178, 
      n7182, n7183, n7184, n7187, n7190, n7193, n7196, n7238, n7241, n7244, 
      n7245, n7246, n7247, n7248, n7249, n7250, n7254, n7255, n7256, n7259, 
      n7262, n7265, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7278, 
      n7279, n7280, n7283, n7286, n7289, n7292, n7293, n7294, n7295, n7296, 
      n7297, n7298, n7302, n7303, n7304, n7307, n7310, n7313, n7316, n7317, 
      n7318, n7319, n7320, n7321, n7322, n7326, n7327, n7328, n7331, n7334, 
      n7337, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7350, n7351, 
      n7352, n7355, n7358, n7361, n7364, n7365, n7366, n7367, n7368, n7369, 
      n7370, n7374, n7375, n7376, n7379, n7382, n7385, n7388, n7389, n7390, 
      n7391, n7392, n7393, n7394, n7398, n7399, n7400, n7403, n7406, n7409, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7422, n7423, n7424, 
      n7427, n7430, n7433, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7446, n7447, n7448, n7451, n7454, n7457, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7470, n7471, n7472, n7475, n7478, n7481, n7484, 
      n7485, n7486, n7487, n7488, n7489, n7490, n7496, n7498, n7502, n7504, 
      n7508, n7510, n7514, n7516, n7520, n7522, n7526, n7528, n7532, n7534, 
      n7538, n7540, n7544, n7546, n7550, n7552, n7556, n7558, n7562, n7564, 
      n7574, n7576, n7580, n7582, n7586, n7588, n7592, n7594, n7598, n7600, 
      n7604, n7606, n7610, n7612, n7616, n7618, n7622, n7624, n7628, n7630, 
      n7634, n7636, n7640, n7642, n7646, n7648, n7652, n7654, n7658, n7660, 
      n7664, n7666, n7670, n7672, n7676, n7678, n7682, n7684, n7686, n7688, 
      n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, 
      n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, 
      n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, 
      n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, 
      n7730, n7731, n7732, n7734, n7735, n7736, n7737, n7740, n7741, n7742, 
      n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
      n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
      n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, 
      n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, 
      n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7853, n7854, 
      n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, 
      n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, 
      n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, 
      n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, 
      n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, 
      n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, 
      n7915, n7916, n7917, n7918, n7919, n7921, n7922, n7923, n7924, n7925, 
      n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, 
      n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, 
      n7946, n7947, n7948, n7949, n7950, n7951, n7953, n7954, n7955, n7956, 
      n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, 
      n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, 
      n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7985, n7986, n7987, 
      n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, 
      n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, 
      n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8017, n8018, 
      n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, 
      n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, 
      n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8049, 
      n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, 
      n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, 
      n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, 
      n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, 
      n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, 
      n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, 
      n8111, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, 
      n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, 
      n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, 
      n8142, n8143, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, 
      n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, 
      n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, 
      n8173, n8174, n8175, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, 
      n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, 
      n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, 
      n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, 
      n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, 
      n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, 
      n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8353, n8354, n8385, 
      n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, 
      n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, 
      n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
      n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, 
      n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, 
      n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, 
      n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, 
      n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, 
      n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
      n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, 
      n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, 
      n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8576, n8577, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
      n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, 
      n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, 
      n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, 
      n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, 
      n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, 
      n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, 
      n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, 
      n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, 
      n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, 
      n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, 
      n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, 
      n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
      n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, 
      n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, 
      n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, 
      n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, 
      n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, 
      n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, 
      n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, 
      n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, 
      n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, 
      n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, 
      n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, 
      n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, 
      n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, 
      n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, 
      n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
      n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, 
      n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8898, n8902, 
      n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, 
      n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, 
      n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, 
      n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, 
      n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, 
      n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
      n8963, n8964, n8965, n727, n731, n734, n735, n736, n743, n752, n756, n761
      , n762, n763, n770, n774, n777, n784, n786, n791, n795, n798, n799, n800,
      n801, n802, n803, n805, n806, n807, n810, n811, n812, n814, n815, n816, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n6754, n6760,
      n6771, n6773, n6778, n6781, n6787, n6795, n6799, n6805, n6817, n6820, 
      n6826, n6832, n6843, n6845, n6853, n6859, n6868, n6871, n6880, n6889, 
      n6893, n6898, n6907, n6915, n6919, n6925, n6937, n6940, n6946, n6952, 
      n6963, n6965, n6973, n6979, n7013, n7018, n7026, n7032, n7036, n7039, 
      n7044, n7047, n7051, n7056, n7060, n7063, n7068, n7071, n7075, n7080, 
      n7084, n7087, n7092, n7095, n7099, n7104, n7107, n7108, n7113, n7114, 
      n7116, n7117, n7119, n7120, n7122, n7123, n7125, n7128, n7129, n7131, 
      n7132, n7133, n7135, n7137, n7138, n7140, n7141, n7143, n7153, n7155, 
      n7156, n7157, n7179, n7180, n7181, n7203, n7204, n7205, n7469, n7491, 
      n7492, n7493, n7494, n7495, n7497, n7499, n7500, n7501, n7503, n7505, 
      n7506, n7507, n7509, n7511, n7512, n7513, n7515, n7517, n7519, n7521, 
      n7523, n7524, n7525, n7527, n7529, n7530, n7531, n7533, n7535, n7584, 
      n7585, n7587, n7589, n7590, n7591, n7593, n7595, n7596, n7597, n7599, 
      n7601, n7602, n7603, n7605, n7607, n7608, n7609, n7611, n7613, n7614, 
      n7615, n7617, n7619, n7620, n7621, n7623, n7625, n7626, n7627, n7629, 
      n7631, n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n79, n80, 
      n85, n86, n91, n92, n97, n98, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n728, n729, n730, n732, 
      n733, n737, n738, n739, n740, n741, n742, n744, n745, n746, n747, n748, 
      n749, n750, n751, n755, n757, n758, n759, n760, n764, n765, n766, n767, 
      n768, n769, n771, n772, n773, n775, n776, n778, n779, n780, n781, n782, 
      n783, n785, n787, n788, n789, n790, n792, n793, n794, n796, n797, n804, 
      n808, n809, n813, n819, n898, n900, n904, n906, n910, n912, n916, n918, 
      n922, n924, n928, n930, n934, n936, n940, n942, n946, n948, n952, n954, 
      n958, n960, n964, n966, n970, n972, n976, n978, n982, n984, n988, n990, 
      n994, n996, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008
      , n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
      n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
      n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
      n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
      n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, 
      n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
      n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
      n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
      n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
      n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
      n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, 
      n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2524, n2525, n2526, n2527, n2528, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2558, n2559, n2563, n2565, 
      n2566, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
      n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, 
      n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, 
      n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, 
      n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, 
      n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
      n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2770, n2771, n2772, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
      n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
      n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
      n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2865, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
      n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, 
      n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, 
      n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
      n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, 
      n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, 
      n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
      n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, 
      n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, 
      n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, 
      n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, 
      n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, 
      n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, 
      n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, 
      n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, 
      n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, 
      n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
      n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, 
      n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, 
      n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, 
      n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6729, n6730, n6732, n6733, n6735, n6736, n6738, n6739, 
      n6747, n6748, n6749, n6751, n6753, n6757, n6759, n6763, n6769, n6772, 
      n6775, n6777, n6780, n6783, n6784, n6793, n6796, n6797, n6801, n6802, 
      n6807, n6808, n6811, n6819, n6821, n6823, n6825, n7325, n7329, n13220, 
      n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, 
      n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, 
      n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, 
      n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, 
      n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, 
      n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, 
      n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, 
      n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, 
      n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, 
      n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, 
      n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, 
      n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, 
      n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, 
      n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, 
      n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, 
      n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, 
      n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, 
      n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, 
      n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, 
      n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, 
      n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, 
      n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, 
      n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, 
      n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, 
      n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, 
      n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, 
      n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, 
      n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, 
      n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, 
      n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, 
      n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, 
      n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, 
      n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, 
      n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, 
      n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, 
      n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, 
      n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, 
      n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, 
      n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, 
      n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, 
      n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, 
      n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, 
      n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, 
      n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, 
      n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, 
      n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, 
      n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, 
      n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, 
      n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, 
      n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, 
      n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, 
      n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, 
      n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, 
      n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, 
      n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, 
      n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, 
      n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, 
      n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, 
      n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, 
      n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, 
      n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, 
      n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, 
      n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, 
      n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, 
      n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, 
      n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, 
      n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, 
      n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, 
      n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, 
      n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, 
      n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, 
      n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, 
      n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, 
      n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, 
      n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, 
      n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, 
      n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, 
      n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, 
      n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, 
      n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, 
      n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, 
      n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, 
      n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, 
      n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, 
      n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, 
      n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, 
      n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, 
      n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, 
      n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, 
      n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, 
      n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, 
      n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, 
      n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, 
      n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, 
      n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, 
      n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, 
      n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, 
      n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, 
      n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, 
      n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, 
      n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, 
      n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, 
      n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, 
      n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, 
      n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, 
      n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, 
      n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, 
      n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, 
      n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, 
      n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, 
      n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, 
      n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, 
      n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, 
      n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, 
      n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, 
      n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, 
      n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, 
      n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, 
      n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, 
      n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, 
      n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, 
      n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, 
      n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, 
      n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, 
      n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, 
      n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, 
      n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, 
      n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, 
      n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, 
      n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, 
      n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, 
      n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, 
      n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, 
      n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, 
      n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, 
      n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, 
      n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, 
      n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, 
      n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, 
      n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, 
      n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, 
      n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, 
      n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, 
      n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, 
      n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, 
      n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, 
      n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, 
      n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, 
      n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, 
      n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, 
      n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, 
      n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, 
      n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, 
      n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, 
      n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, 
      n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, 
      n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, 
      n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, 
      n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, 
      n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, 
      n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, 
      n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, 
      n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, 
      n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, 
      n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, 
      n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, 
      n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, 
      n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, 
      n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, 
      n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
      n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, 
      n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, 
      n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, 
      n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, 
      n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, 
      n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, 
      n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, 
      n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, 
      n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, 
      n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, 
      n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, 
      n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, 
      n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, 
      n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, 
      n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, 
      n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, 
      n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, 
      n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, 
      n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, 
      n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, 
      n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, 
      n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, 
      n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, 
      n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, 
      n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, 
      n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, 
      n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, 
      n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, 
      n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, 
      n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, 
      n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, 
      n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, 
      n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, 
      n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, 
      n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, 
      n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, 
      n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, 
      n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, 
      n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, 
      n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, 
      n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, 
      n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, 
      n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, 
      n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, 
      n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, 
      n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, 
      n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, 
      n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, 
      n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, 
      n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, 
      n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, 
      n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, 
      n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, 
      n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, 
      n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, 
      n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, 
      n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, 
      n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, 
      n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, 
      n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, 
      n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, 
      n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, 
      n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, 
      n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, 
      n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, 
      n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, 
      n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, 
      n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, 
      n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, 
      n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, 
      n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, 
      n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, 
      n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, 
      n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, 
      n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, 
      n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, 
      n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, 
      n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, 
      n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, 
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, 
      n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, 
      n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, 
      n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781 : 
      std_logic;

begin
   
   OUT1_tri_enable_reg_31_inst : DFF_X1 port map( D => n9006, CK => CLK, Q => 
                           n8902, QN => n2277);
   OUT1_tri_enable_reg_30_inst : DFF_X1 port map( D => n9007, CK => CLK, Q => 
                           n8903, QN => n2276);
   OUT1_tri_enable_reg_29_inst : DFF_X1 port map( D => n9008, CK => CLK, Q => 
                           n8904, QN => n2275);
   OUT1_tri_enable_reg_28_inst : DFF_X1 port map( D => n9009, CK => CLK, Q => 
                           n8905, QN => n2274);
   OUT1_tri_enable_reg_27_inst : DFF_X1 port map( D => n9010, CK => CLK, Q => 
                           n8906, QN => n2273);
   OUT1_tri_enable_reg_26_inst : DFF_X1 port map( D => n9011, CK => CLK, Q => 
                           n8907, QN => n2272);
   OUT1_tri_enable_reg_25_inst : DFF_X1 port map( D => n9012, CK => CLK, Q => 
                           n8908, QN => n2271);
   OUT1_tri_enable_reg_24_inst : DFF_X1 port map( D => n9013, CK => CLK, Q => 
                           n8909, QN => n2270);
   OUT1_tri_enable_reg_23_inst : DFF_X1 port map( D => n9014, CK => CLK, Q => 
                           n8910, QN => n2269);
   OUT1_tri_enable_reg_22_inst : DFF_X1 port map( D => n9015, CK => CLK, Q => 
                           n8911, QN => n2268);
   OUT1_tri_enable_reg_21_inst : DFF_X1 port map( D => n9016, CK => CLK, Q => 
                           n8912, QN => n2267);
   OUT1_tri_enable_reg_20_inst : DFF_X1 port map( D => n9017, CK => CLK, Q => 
                           n8913, QN => n2266);
   OUT1_tri_enable_reg_19_inst : DFF_X1 port map( D => n9018, CK => CLK, Q => 
                           n8914, QN => n2265);
   OUT1_tri_enable_reg_18_inst : DFF_X1 port map( D => n9019, CK => CLK, Q => 
                           n8915, QN => n2264);
   OUT1_tri_enable_reg_17_inst : DFF_X1 port map( D => n9020, CK => CLK, Q => 
                           n8916, QN => n2263);
   OUT1_tri_enable_reg_16_inst : DFF_X1 port map( D => n9021, CK => CLK, Q => 
                           n8917, QN => n2262);
   OUT1_tri_enable_reg_15_inst : DFF_X1 port map( D => n9022, CK => CLK, Q => 
                           n8918, QN => n2261);
   OUT1_tri_enable_reg_14_inst : DFF_X1 port map( D => n9023, CK => CLK, Q => 
                           n8919, QN => n2260);
   OUT1_tri_enable_reg_13_inst : DFF_X1 port map( D => n9024, CK => CLK, Q => 
                           n8920, QN => n2259);
   OUT1_tri_enable_reg_12_inst : DFF_X1 port map( D => n9025, CK => CLK, Q => 
                           n8921, QN => n2258);
   OUT1_tri_enable_reg_11_inst : DFF_X1 port map( D => n9026, CK => CLK, Q => 
                           n8922, QN => n2257);
   OUT1_tri_enable_reg_10_inst : DFF_X1 port map( D => n9027, CK => CLK, Q => 
                           n8923, QN => n2256);
   OUT1_tri_enable_reg_9_inst : DFF_X1 port map( D => n9028, CK => CLK, Q => 
                           n8924, QN => n2255);
   OUT1_tri_enable_reg_8_inst : DFF_X1 port map( D => n9029, CK => CLK, Q => 
                           n8925, QN => n2254);
   OUT1_tri_enable_reg_7_inst : DFF_X1 port map( D => n9030, CK => CLK, Q => 
                           n8926, QN => n2253);
   OUT1_tri_enable_reg_6_inst : DFF_X1 port map( D => n9031, CK => CLK, Q => 
                           n8927, QN => n2252);
   OUT1_tri_enable_reg_5_inst : DFF_X1 port map( D => n9032, CK => CLK, Q => 
                           n8928, QN => n2251);
   OUT1_tri_enable_reg_4_inst : DFF_X1 port map( D => n9033, CK => CLK, Q => 
                           n8929, QN => n2250);
   OUT1_tri_enable_reg_3_inst : DFF_X1 port map( D => n9034, CK => CLK, Q => 
                           n8930, QN => n2249);
   OUT1_tri_enable_reg_2_inst : DFF_X1 port map( D => n9035, CK => CLK, Q => 
                           n8931, QN => n2248);
   OUT1_tri_enable_reg_1_inst : DFF_X1 port map( D => n9036, CK => CLK, Q => 
                           n8932, QN => n2247);
   OUT1_tri_enable_reg_0_inst : DFF_X1 port map( D => n9037, CK => CLK, Q => 
                           n8933, QN => n2246);
   OUT2_tri_enable_reg_31_inst : DFF_X1 port map( D => n9038, CK => CLK, Q => 
                           n8934, QN => n2245);
   OUT2_tri_enable_reg_30_inst : DFF_X1 port map( D => n9039, CK => CLK, Q => 
                           n8935, QN => n2244);
   OUT2_tri_enable_reg_29_inst : DFF_X1 port map( D => n9040, CK => CLK, Q => 
                           n8936, QN => n2243);
   OUT2_tri_enable_reg_28_inst : DFF_X1 port map( D => n9041, CK => CLK, Q => 
                           n8937, QN => n2242);
   OUT2_tri_enable_reg_27_inst : DFF_X1 port map( D => n9042, CK => CLK, Q => 
                           n8938, QN => n2241);
   OUT2_tri_enable_reg_26_inst : DFF_X1 port map( D => n9043, CK => CLK, Q => 
                           n8939, QN => n2240);
   OUT2_tri_enable_reg_25_inst : DFF_X1 port map( D => n9044, CK => CLK, Q => 
                           n8940, QN => n2239);
   OUT2_tri_enable_reg_24_inst : DFF_X1 port map( D => n9045, CK => CLK, Q => 
                           n8941, QN => n2238);
   OUT2_tri_enable_reg_23_inst : DFF_X1 port map( D => n9046, CK => CLK, Q => 
                           n8942, QN => n2237);
   OUT2_tri_enable_reg_22_inst : DFF_X1 port map( D => n9047, CK => CLK, Q => 
                           n8943, QN => n2236);
   OUT2_tri_enable_reg_21_inst : DFF_X1 port map( D => n9048, CK => CLK, Q => 
                           n8944, QN => n2235);
   OUT2_tri_enable_reg_20_inst : DFF_X1 port map( D => n9049, CK => CLK, Q => 
                           n8945, QN => n2234);
   OUT2_tri_enable_reg_19_inst : DFF_X1 port map( D => n9050, CK => CLK, Q => 
                           n8946, QN => n2233);
   OUT2_tri_enable_reg_18_inst : DFF_X1 port map( D => n9051, CK => CLK, Q => 
                           n8947, QN => n2232);
   OUT2_tri_enable_reg_17_inst : DFF_X1 port map( D => n9052, CK => CLK, Q => 
                           n8948, QN => n2231);
   OUT2_tri_enable_reg_16_inst : DFF_X1 port map( D => n9053, CK => CLK, Q => 
                           n8949, QN => n2230);
   OUT2_tri_enable_reg_15_inst : DFF_X1 port map( D => n9054, CK => CLK, Q => 
                           n8950, QN => n2229);
   OUT2_tri_enable_reg_14_inst : DFF_X1 port map( D => n9055, CK => CLK, Q => 
                           n8951, QN => n2228);
   OUT2_tri_enable_reg_13_inst : DFF_X1 port map( D => n9056, CK => CLK, Q => 
                           n8952, QN => n2227);
   OUT2_tri_enable_reg_12_inst : DFF_X1 port map( D => n9057, CK => CLK, Q => 
                           n8953, QN => n2226);
   OUT2_tri_enable_reg_11_inst : DFF_X1 port map( D => n9058, CK => CLK, Q => 
                           n8954, QN => n2225);
   OUT2_tri_enable_reg_10_inst : DFF_X1 port map( D => n9059, CK => CLK, Q => 
                           n8955, QN => n2224);
   OUT2_tri_enable_reg_9_inst : DFF_X1 port map( D => n9060, CK => CLK, Q => 
                           n8956, QN => n2223);
   OUT2_tri_enable_reg_8_inst : DFF_X1 port map( D => n9061, CK => CLK, Q => 
                           n8957, QN => n2222);
   OUT2_tri_enable_reg_7_inst : DFF_X1 port map( D => n9062, CK => CLK, Q => 
                           n8958, QN => n2221);
   OUT2_tri_enable_reg_6_inst : DFF_X1 port map( D => n9063, CK => CLK, Q => 
                           n8959, QN => n2220);
   OUT2_tri_enable_reg_5_inst : DFF_X1 port map( D => n9064, CK => CLK, Q => 
                           n8960, QN => n2219);
   OUT2_tri_enable_reg_4_inst : DFF_X1 port map( D => n9065, CK => CLK, Q => 
                           n8961, QN => n2218);
   OUT2_tri_enable_reg_3_inst : DFF_X1 port map( D => n9066, CK => CLK, Q => 
                           n8962, QN => n2217);
   OUT2_tri_enable_reg_2_inst : DFF_X1 port map( D => n9067, CK => CLK, Q => 
                           n8963, QN => n2216);
   OUT2_tri_enable_reg_1_inst : DFF_X1 port map( D => n9068, CK => CLK, Q => 
                           n8964, QN => n2215);
   OUT2_tri_enable_reg_0_inst : DFF_X1 port map( D => n9069, CK => CLK, Q => 
                           n8965, QN => n2214);
   RFtoMEM_BUS_reg_31_inst : DFF_X1 port map( D => n9134, CK => CLK, Q => 
                           RFtoMEM_BUS(31), QN => n7631);
   RFtoMEM_BUS_reg_30_inst : DFF_X1 port map( D => n9168, CK => CLK, Q => 
                           RFtoMEM_BUS(30), QN => n7629);
   RFtoMEM_BUS_reg_29_inst : DFF_X1 port map( D => n9170, CK => CLK, Q => 
                           RFtoMEM_BUS(29), QN => n7627);
   RFtoMEM_BUS_reg_28_inst : DFF_X1 port map( D => n9172, CK => CLK, Q => 
                           RFtoMEM_BUS(28), QN => n7626);
   RFtoMEM_BUS_reg_27_inst : DFF_X1 port map( D => n9174, CK => CLK, Q => 
                           RFtoMEM_BUS(27), QN => n7625);
   RFtoMEM_BUS_reg_26_inst : DFF_X1 port map( D => n9176, CK => CLK, Q => 
                           RFtoMEM_BUS(26), QN => n7623);
   RFtoMEM_BUS_reg_25_inst : DFF_X1 port map( D => n9178, CK => CLK, Q => 
                           RFtoMEM_BUS(25), QN => n7621);
   RFtoMEM_BUS_reg_24_inst : DFF_X1 port map( D => n9180, CK => CLK, Q => 
                           RFtoMEM_BUS(24), QN => n7620);
   RFtoMEM_BUS_reg_23_inst : DFF_X1 port map( D => n9182, CK => CLK, Q => 
                           RFtoMEM_BUS(23), QN => n7619);
   RFtoMEM_BUS_reg_22_inst : DFF_X1 port map( D => n9184, CK => CLK, Q => 
                           RFtoMEM_BUS(22), QN => n7617);
   RFtoMEM_BUS_reg_21_inst : DFF_X1 port map( D => n9186, CK => CLK, Q => 
                           RFtoMEM_BUS(21), QN => n7615);
   RFtoMEM_BUS_reg_20_inst : DFF_X1 port map( D => n9188, CK => CLK, Q => 
                           RFtoMEM_BUS(20), QN => n7614);
   RFtoMEM_BUS_reg_19_inst : DFF_X1 port map( D => n9190, CK => CLK, Q => 
                           RFtoMEM_BUS(19), QN => n7613);
   RFtoMEM_BUS_reg_18_inst : DFF_X1 port map( D => n9192, CK => CLK, Q => 
                           RFtoMEM_BUS(18), QN => n7611);
   RFtoMEM_BUS_reg_17_inst : DFF_X1 port map( D => n9194, CK => CLK, Q => 
                           RFtoMEM_BUS(17), QN => n7609);
   RFtoMEM_BUS_reg_16_inst : DFF_X1 port map( D => n9196, CK => CLK, Q => 
                           RFtoMEM_BUS(16), QN => n7608);
   RFtoMEM_BUS_reg_15_inst : DFF_X1 port map( D => n9198, CK => CLK, Q => 
                           RFtoMEM_BUS(15), QN => n7607);
   RFtoMEM_BUS_reg_14_inst : DFF_X1 port map( D => n9200, CK => CLK, Q => 
                           RFtoMEM_BUS(14), QN => n7605);
   RFtoMEM_BUS_reg_13_inst : DFF_X1 port map( D => n9202, CK => CLK, Q => 
                           RFtoMEM_BUS(13), QN => n7603);
   RFtoMEM_BUS_reg_12_inst : DFF_X1 port map( D => n9204, CK => CLK, Q => 
                           RFtoMEM_BUS(12), QN => n7602);
   RFtoMEM_BUS_reg_11_inst : DFF_X1 port map( D => n9206, CK => CLK, Q => 
                           RFtoMEM_BUS(11), QN => n7601);
   RFtoMEM_BUS_reg_10_inst : DFF_X1 port map( D => n9208, CK => CLK, Q => 
                           RFtoMEM_BUS(10), QN => n7599);
   RFtoMEM_BUS_reg_9_inst : DFF_X1 port map( D => n9210, CK => CLK, Q => 
                           RFtoMEM_BUS(9), QN => n7597);
   RFtoMEM_BUS_reg_8_inst : DFF_X1 port map( D => n9212, CK => CLK, Q => 
                           RFtoMEM_BUS(8), QN => n7596);
   RFtoMEM_BUS_reg_7_inst : DFF_X1 port map( D => n9214, CK => CLK, Q => 
                           RFtoMEM_BUS(7), QN => n7595);
   RFtoMEM_BUS_reg_6_inst : DFF_X1 port map( D => n9216, CK => CLK, Q => 
                           RFtoMEM_BUS(6), QN => n7593);
   RFtoMEM_BUS_reg_5_inst : DFF_X1 port map( D => n9218, CK => CLK, Q => 
                           RFtoMEM_BUS(5), QN => n7591);
   RFtoMEM_BUS_reg_4_inst : DFF_X1 port map( D => n9220, CK => CLK, Q => 
                           RFtoMEM_BUS(4), QN => n7590);
   RFtoMEM_BUS_reg_3_inst : DFF_X1 port map( D => n9222, CK => CLK, Q => 
                           RFtoMEM_BUS(3), QN => n7589);
   RFtoMEM_BUS_reg_2_inst : DFF_X1 port map( D => n9224, CK => CLK, Q => 
                           RFtoMEM_BUS(2), QN => n7587);
   RFtoMEM_BUS_reg_1_inst : DFF_X1 port map( D => n9226, CK => CLK, Q => 
                           RFtoMEM_BUS(1), QN => n7585);
   RFtoMEM_BUS_reg_0_inst : DFF_X1 port map( D => n11501, CK => CLK, Q => 
                           RFtoMEM_BUS(0), QN => n7584);
   OUT1_reg_22_inst : DFF_X1 port map( D => n9144, CK => CLK, Q => n_1000, QN 
                           => n2172);
   OUT1_reg_21_inst : DFF_X1 port map( D => n9145, CK => CLK, Q => n_1001, QN 
                           => n2171);
   OUT1_reg_20_inst : DFF_X1 port map( D => n9146, CK => CLK, Q => n_1002, QN 
                           => n2170);
   U21 : TINV_X1 port map( I => n2181, EN => n8902, ZN => OUT1(31));
   U22 : TINV_X1 port map( I => n2180, EN => n8903, ZN => OUT1(30));
   U23 : TINV_X1 port map( I => n2179, EN => n8904, ZN => OUT1(29));
   U24 : TINV_X1 port map( I => n2178, EN => n8905, ZN => OUT1(28));
   U25 : TINV_X1 port map( I => n2177, EN => n8906, ZN => OUT1(27));
   U26 : TINV_X1 port map( I => n2176, EN => n8907, ZN => OUT1(26));
   U27 : TINV_X1 port map( I => n2175, EN => n8908, ZN => OUT1(25));
   U28 : TINV_X1 port map( I => n2174, EN => n8909, ZN => OUT1(24));
   U29 : TINV_X1 port map( I => n2173, EN => n8910, ZN => OUT1(23));
   U30 : TINV_X1 port map( I => n2172, EN => n8911, ZN => OUT1(22));
   U31 : TINV_X1 port map( I => n2171, EN => n8912, ZN => OUT1(21));
   U32 : TINV_X1 port map( I => n2170, EN => n8913, ZN => OUT1(20));
   U33 : TINV_X1 port map( I => n2169, EN => n8914, ZN => OUT1(19));
   U34 : TINV_X1 port map( I => n2168, EN => n8915, ZN => OUT1(18));
   U35 : TINV_X1 port map( I => n2167, EN => n8916, ZN => OUT1(17));
   U36 : TINV_X1 port map( I => n2166, EN => n8917, ZN => OUT1(16));
   U37 : TINV_X1 port map( I => n2165, EN => n8918, ZN => OUT1(15));
   U38 : TINV_X1 port map( I => n2164, EN => n8919, ZN => OUT1(14));
   U39 : TINV_X1 port map( I => n2163, EN => n8920, ZN => OUT1(13));
   U40 : TINV_X1 port map( I => n2162, EN => n8921, ZN => OUT1(12));
   U41 : TINV_X1 port map( I => n2161, EN => n8922, ZN => OUT1(11));
   U42 : TINV_X1 port map( I => n2160, EN => n8923, ZN => OUT1(10));
   U43 : TINV_X1 port map( I => n2159, EN => n8924, ZN => OUT1(9));
   U44 : TINV_X1 port map( I => n2158, EN => n8925, ZN => OUT1(8));
   U45 : TINV_X1 port map( I => n2157, EN => n8926, ZN => OUT1(7));
   U46 : TINV_X1 port map( I => n2156, EN => n8927, ZN => OUT1(6));
   U47 : TINV_X1 port map( I => n2155, EN => n8928, ZN => OUT1(5));
   U48 : TINV_X1 port map( I => n2154, EN => n8929, ZN => OUT1(4));
   U49 : TINV_X1 port map( I => n2153, EN => n8930, ZN => OUT1(3));
   U50 : TINV_X1 port map( I => n2152, EN => n8931, ZN => OUT1(2));
   U51 : TINV_X1 port map( I => n2151, EN => n8932, ZN => OUT1(1));
   U52 : TINV_X1 port map( I => n2150, EN => n8933, ZN => OUT1(0));
   U53 : TINV_X1 port map( I => n2213, EN => n8934, ZN => OUT2(31));
   U54 : TINV_X1 port map( I => n2212, EN => n8935, ZN => OUT2(30));
   U55 : TINV_X1 port map( I => n2211, EN => n8936, ZN => OUT2(29));
   U56 : TINV_X1 port map( I => n2210, EN => n8937, ZN => OUT2(28));
   U57 : TINV_X1 port map( I => n2209, EN => n8938, ZN => OUT2(27));
   U58 : TINV_X1 port map( I => n2208, EN => n8939, ZN => OUT2(26));
   U59 : TINV_X1 port map( I => n2207, EN => n8940, ZN => OUT2(25));
   U60 : TINV_X1 port map( I => n2206, EN => n8941, ZN => OUT2(24));
   U61 : TINV_X1 port map( I => n2205, EN => n8942, ZN => OUT2(23));
   U62 : TINV_X1 port map( I => n2204, EN => n8943, ZN => OUT2(22));
   U63 : TINV_X1 port map( I => n2203, EN => n8944, ZN => OUT2(21));
   U64 : TINV_X1 port map( I => n2202, EN => n8945, ZN => OUT2(20));
   U65 : TINV_X1 port map( I => n2201, EN => n8946, ZN => OUT2(19));
   U66 : TINV_X1 port map( I => n2200, EN => n8947, ZN => OUT2(18));
   U67 : TINV_X1 port map( I => n2199, EN => n8948, ZN => OUT2(17));
   U68 : TINV_X1 port map( I => n2198, EN => n8949, ZN => OUT2(16));
   U69 : TINV_X1 port map( I => n2197, EN => n8950, ZN => OUT2(15));
   U70 : TINV_X1 port map( I => n2196, EN => n8951, ZN => OUT2(14));
   U71 : TINV_X1 port map( I => n2195, EN => n8952, ZN => OUT2(13));
   U72 : TINV_X1 port map( I => n2194, EN => n8953, ZN => OUT2(12));
   U73 : TINV_X1 port map( I => n2193, EN => n8954, ZN => OUT2(11));
   U74 : TINV_X1 port map( I => n2192, EN => n8955, ZN => OUT2(10));
   U75 : TINV_X1 port map( I => n2191, EN => n8956, ZN => OUT2(9));
   U76 : TINV_X1 port map( I => n2190, EN => n8957, ZN => OUT2(8));
   U77 : TINV_X1 port map( I => n2189, EN => n8958, ZN => OUT2(7));
   U78 : TINV_X1 port map( I => n2188, EN => n8959, ZN => OUT2(6));
   U79 : TINV_X1 port map( I => n2187, EN => n8960, ZN => OUT2(5));
   U80 : TINV_X1 port map( I => n2186, EN => n8961, ZN => OUT2(4));
   U81 : TINV_X1 port map( I => n2185, EN => n8962, ZN => OUT2(3));
   U82 : TINV_X1 port map( I => n2184, EN => n8963, ZN => OUT2(2));
   U83 : TINV_X1 port map( I => n2183, EN => n8964, ZN => OUT2(1));
   U84 : TINV_X1 port map( I => n2182, EN => n8965, ZN => OUT2(0));
   U3271 : NOR4_X2 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(5), A4 => ADD_RD1(6), ZN => n5198);
   U4617 : NOR4_X2 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(5), A4 => ADD_RD2(6), ZN => n6519);
   U4711 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n6508);
   U8869 : NAND3_X1 port map( A1 => n2524, A2 => n14685, A3 => n2585, ZN => 
                           n2628);
   U8870 : NAND3_X1 port map( A1 => n2524, A2 => n14502, A3 => n2573, ZN => 
                           n2664);
   U8871 : NAND3_X1 port map( A1 => n2524, A2 => n14493, A3 => n2577, ZN => 
                           n2669);
   U8872 : NAND3_X1 port map( A1 => n2524, A2 => n14484, A3 => n2572, ZN => 
                           n2674);
   U8873 : NAND3_X1 port map( A1 => n2524, A2 => n14475, A3 => n2576, ZN => 
                           n2679);
   U8874 : NAND3_X1 port map( A1 => n2524, A2 => n14466, A3 => n2571, ZN => 
                           n2684);
   U8875 : NAND3_X1 port map( A1 => n2524, A2 => n14457, A3 => n2575, ZN => 
                           n2689);
   U8876 : NAND3_X1 port map( A1 => n2524, A2 => n14448, A3 => n2570, ZN => 
                           n2694);
   U8877 : NAND3_X1 port map( A1 => n2524, A2 => n14439, A3 => n2574, ZN => 
                           n2699);
   U8878 : NAND3_X1 port map( A1 => n2528, A2 => n14430, A3 => n2581, ZN => 
                           n2704);
   U8879 : NAND3_X1 port map( A1 => n2528, A2 => n14421, A3 => n2584, ZN => 
                           n2711);
   U8880 : NAND3_X1 port map( A1 => n2528, A2 => n14412, A3 => n2580, ZN => 
                           n2716);
   U8881 : NAND3_X1 port map( A1 => n2528, A2 => n14403, A3 => n2583, ZN => 
                           n2721);
   U8882 : NAND3_X1 port map( A1 => n2528, A2 => n14394, A3 => n2579, ZN => 
                           n2726);
   U8883 : NAND3_X1 port map( A1 => n2528, A2 => n14385, A3 => n2582, ZN => 
                           n2731);
   U8884 : NAND3_X1 port map( A1 => n2578, A2 => n14376, A3 => n2528, ZN => 
                           n2736);
   U8885 : NAND3_X1 port map( A1 => n2585, A2 => n14367, A3 => n2528, ZN => 
                           n2741);
   U8886 : NAND3_X1 port map( A1 => n2529, A2 => n14358, A3 => n13221, ZN => 
                           n2745);
   U8887 : NAND3_X1 port map( A1 => n2529, A2 => n14347, A3 => n14730, ZN => 
                           n2750);
   U8888 : NAND3_X1 port map( A1 => n2529, A2 => n14338, A3 => n14736, ZN => 
                           n2754);
   U8889 : NAND3_X1 port map( A1 => n2529, A2 => n14329, A3 => n14733, ZN => 
                           n2758);
   U8890 : NAND3_X1 port map( A1 => n2529, A2 => n14320, A3 => n14727, ZN => 
                           n2762);
   U8891 : NAND3_X1 port map( A1 => n2529, A2 => n14311, A3 => n13224, ZN => 
                           n2766);
   U8892 : NAND3_X1 port map( A1 => n2529, A2 => n14300, A3 => n13222, ZN => 
                           n2770);
   U8893 : NAND3_X1 port map( A1 => n2529, A2 => n14289, A3 => n13225, ZN => 
                           n2774);
   U8894 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD1(6), Z => n5236);
   U8895 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD1(5), Z => n5235);
   U8896 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD1(4), Z => n5234);
   U8897 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD1(3), Z => n5233);
   U8898 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD1(0), Z => n5237);
   U8899 : XOR2_X1 port map( A => n2537, B => ADD_RD1(1), Z => n5230);
   U8900 : XOR2_X1 port map( A => n2536, B => ADD_RD1(2), Z => n5229);
   U8901 : XOR2_X1 port map( A => ADD_WR(6), B => ADD_RD2(6), Z => n6557);
   U8902 : XOR2_X1 port map( A => ADD_WR(5), B => ADD_RD2(5), Z => n6556);
   U8903 : XOR2_X1 port map( A => ADD_WR(4), B => ADD_RD2(4), Z => n6555);
   U8904 : XOR2_X1 port map( A => ADD_WR(3), B => ADD_RD2(3), Z => n6554);
   U8905 : XOR2_X1 port map( A => ADD_WR(0), B => ADD_RD2(0), Z => n6558);
   U8906 : XOR2_X1 port map( A => n2537, B => ADD_RD2(1), Z => n6551);
   U8907 : XOR2_X1 port map( A => n2536, B => ADD_RD2(2), Z => n6550);
   U8908 : NAND3_X1 port map( A1 => n6572, A2 => n2589, A3 => ADD_SF(6), ZN => 
                           n2803);
   U8909 : NAND3_X1 port map( A1 => n6572, A2 => ADD_SF(0), A3 => ADD_SF(6), ZN
                           => n2802);
   U8910 : NAND3_X1 port map( A1 => n6573, A2 => ADD_SF(0), A3 => ADD_SF(6), ZN
                           => n2808);
   U8911 : NAND3_X1 port map( A1 => n6574, A2 => n2589, A3 => ADD_SF(6), ZN => 
                           n2807);
   U8912 : NAND3_X1 port map( A1 => n2573, A2 => n13633, A3 => n2527, ZN => 
                           n6605);
   U8913 : NAND3_X1 port map( A1 => n2577, A2 => n13624, A3 => n2527, ZN => 
                           n6609);
   U8914 : NAND3_X1 port map( A1 => n2572, A2 => n13615, A3 => n2527, ZN => 
                           n6612);
   U8915 : NAND3_X1 port map( A1 => n2576, A2 => n13606, A3 => n2527, ZN => 
                           n6615);
   U8916 : NAND3_X1 port map( A1 => n2571, A2 => n13597, A3 => n2527, ZN => 
                           n6618);
   U8917 : NAND3_X1 port map( A1 => n2575, A2 => n13588, A3 => n2527, ZN => 
                           n6621);
   U8918 : NAND3_X1 port map( A1 => n2570, A2 => n13579, A3 => n2527, ZN => 
                           n6624);
   U8919 : NAND3_X1 port map( A1 => n2574, A2 => n13570, A3 => n2527, ZN => 
                           n6627);
   U8920 : NAND3_X1 port map( A1 => n6601, A2 => n2529, A3 => ADD_SF(6), ZN => 
                           n6607);
   U8921 : NAND3_X1 port map( A1 => n2581, A2 => n13561, A3 => n2526, ZN => 
                           n6630);
   U8922 : NAND3_X1 port map( A1 => n2584, A2 => n13552, A3 => n2526, ZN => 
                           n6635);
   U8923 : NAND3_X1 port map( A1 => n2580, A2 => n13543, A3 => n2526, ZN => 
                           n6638);
   U8924 : NAND3_X1 port map( A1 => n2583, A2 => n13534, A3 => n2526, ZN => 
                           n6641);
   U8925 : NAND3_X1 port map( A1 => n2579, A2 => n13525, A3 => n2526, ZN => 
                           n6644);
   U8926 : NAND3_X1 port map( A1 => n2582, A2 => n13516, A3 => n2526, ZN => 
                           n6647);
   U8927 : NAND3_X1 port map( A1 => n2578, A2 => n13507, A3 => n2526, ZN => 
                           n6650);
   U8928 : NAND3_X1 port map( A1 => n2585, A2 => n13498, A3 => n2526, ZN => 
                           n6653);
   U8929 : NAND3_X1 port map( A1 => n2573, A2 => n13489, A3 => n2526, ZN => 
                           n6656);
   U8930 : NAND3_X1 port map( A1 => n2577, A2 => n13480, A3 => n2526, ZN => 
                           n6659);
   U8931 : NAND3_X1 port map( A1 => n2572, A2 => n13471, A3 => n2526, ZN => 
                           n6662);
   U8932 : NAND3_X1 port map( A1 => n2576, A2 => n13462, A3 => n2526, ZN => 
                           n6665);
   U8933 : NAND3_X1 port map( A1 => n2571, A2 => n13453, A3 => n2526, ZN => 
                           n6668);
   U8934 : NAND3_X1 port map( A1 => n2575, A2 => n13444, A3 => n2526, ZN => 
                           n6671);
   U8935 : NAND3_X1 port map( A1 => n2570, A2 => n13435, A3 => n2526, ZN => 
                           n6674);
   U8936 : NAND3_X1 port map( A1 => n2574, A2 => n13426, A3 => n2526, ZN => 
                           n6677);
   U8937 : NAND3_X1 port map( A1 => n2581, A2 => n13417, A3 => n2525, ZN => 
                           n6681);
   U8938 : NAND3_X1 port map( A1 => n2584, A2 => n13408, A3 => n2525, ZN => 
                           n6686);
   U8939 : NAND3_X1 port map( A1 => n2580, A2 => n13399, A3 => n2525, ZN => 
                           n6689);
   U8940 : NAND3_X1 port map( A1 => n2583, A2 => n13390, A3 => n2525, ZN => 
                           n6692);
   U8941 : NAND3_X1 port map( A1 => n2579, A2 => n13381, A3 => n2525, ZN => 
                           n6695);
   U8942 : NAND3_X1 port map( A1 => n2582, A2 => n13372, A3 => n2525, ZN => 
                           n6698);
   U8943 : NAND3_X1 port map( A1 => n2578, A2 => n13363, A3 => n2525, ZN => 
                           n6701);
   U8944 : NAND3_X1 port map( A1 => n2585, A2 => n13354, A3 => n2525, ZN => 
                           n6704);
   U8945 : NAND3_X1 port map( A1 => n2573, A2 => n13345, A3 => n2525, ZN => 
                           n6710);
   U8946 : NAND3_X1 port map( A1 => n2577, A2 => n13336, A3 => n2525, ZN => 
                           n6716);
   U8947 : NAND3_X1 port map( A1 => n2572, A2 => n13327, A3 => n2525, ZN => 
                           n6721);
   U8948 : NAND3_X1 port map( A1 => n2576, A2 => n13318, A3 => n2525, ZN => 
                           n6725);
   U8949 : NAND3_X1 port map( A1 => n2571, A2 => n13309, A3 => n2525, ZN => 
                           n6732);
   U8950 : NAND3_X1 port map( A1 => n2575, A2 => n13300, A3 => n2525, ZN => 
                           n6738);
   U8951 : NAND3_X1 port map( A1 => n2570, A2 => n13291, A3 => n2525, ZN => 
                           n6748);
   U8952 : NAND3_X1 port map( A1 => n2574, A2 => n13282, A3 => n2525, ZN => 
                           n6753);
   U8953 : NAND3_X1 port map( A1 => n2524, A2 => n13273, A3 => n2581, ZN => 
                           n6763);
   U8954 : NAND3_X1 port map( A1 => n2524, A2 => n13264, A3 => n2584, ZN => 
                           n6780);
   U8955 : NAND3_X1 port map( A1 => n2524, A2 => n13255, A3 => n2580, ZN => 
                           n6793);
   U8956 : NAND3_X1 port map( A1 => n2524, A2 => n13246, A3 => n2583, ZN => 
                           n6801);
   U8957 : NAND3_X1 port map( A1 => n2524, A2 => n13237, A3 => n2579, ZN => 
                           n6808);
   U8958 : NAND3_X1 port map( A1 => n2524, A2 => n13228, A3 => n2582, ZN => 
                           n6821);
   U8959 : NAND3_X1 port map( A1 => n2524, A2 => n14709, A3 => n2578, ZN => 
                           n2625);
   REGISTERS_reg_70_7_inst : DFF_X1 port map( D => n11461, CK => CLK, Q => n935
                           , QN => n1);
   REGISTERS_reg_70_6_inst : DFF_X1 port map( D => n11462, CK => CLK, Q => n929
                           , QN => n2);
   REGISTERS_reg_70_5_inst : DFF_X1 port map( D => n11463, CK => CLK, Q => n923
                           , QN => n3);
   REGISTERS_reg_70_4_inst : DFF_X1 port map( D => n11464, CK => CLK, Q => n917
                           , QN => n4);
   REGISTERS_reg_70_3_inst : DFF_X1 port map( D => n11465, CK => CLK, Q => n911
                           , QN => n5);
   REGISTERS_reg_70_2_inst : DFF_X1 port map( D => n11466, CK => CLK, Q => n905
                           , QN => n6);
   REGISTERS_reg_70_1_inst : DFF_X1 port map( D => n11467, CK => CLK, Q => n899
                           , QN => n7);
   REGISTERS_reg_68_7_inst : DFF_X1 port map( D => n11397, CK => CLK, Q => 
                           n8886, QN => n8);
   REGISTERS_reg_68_6_inst : DFF_X1 port map( D => n11398, CK => CLK, Q => 
                           n8887, QN => n10);
   REGISTERS_reg_68_5_inst : DFF_X1 port map( D => n11399, CK => CLK, Q => 
                           n8888, QN => n11);
   REGISTERS_reg_68_4_inst : DFF_X1 port map( D => n11400, CK => CLK, Q => 
                           n8889, QN => n12);
   REGISTERS_reg_68_3_inst : DFF_X1 port map( D => n11401, CK => CLK, Q => 
                           n8890, QN => n13);
   REGISTERS_reg_68_2_inst : DFF_X1 port map( D => n11402, CK => CLK, Q => 
                           n8891, QN => n14);
   REGISTERS_reg_68_1_inst : DFF_X1 port map( D => n11403, CK => CLK, Q => 
                           n8892, QN => n15);
   REGISTERS_reg_68_0_inst : DFF_X1 port map( D => n11404, CK => CLK, Q => 
                           n8893, QN => n16);
   REGISTERS_reg_67_7_inst : DFF_X1 port map( D => n11365, CK => CLK, Q => 
                           n8854, QN => n17);
   REGISTERS_reg_67_6_inst : DFF_X1 port map( D => n11366, CK => CLK, Q => 
                           n8855, QN => n18);
   REGISTERS_reg_67_5_inst : DFF_X1 port map( D => n11367, CK => CLK, Q => 
                           n8856, QN => n19);
   REGISTERS_reg_67_4_inst : DFF_X1 port map( D => n11368, CK => CLK, Q => 
                           n8857, QN => n20);
   REGISTERS_reg_67_3_inst : DFF_X1 port map( D => n11369, CK => CLK, Q => 
                           n8858, QN => n21);
   REGISTERS_reg_67_2_inst : DFF_X1 port map( D => n11370, CK => CLK, Q => 
                           n8859, QN => n22);
   REGISTERS_reg_67_1_inst : DFF_X1 port map( D => n11371, CK => CLK, Q => 
                           n8860, QN => n23);
   REGISTERS_reg_67_0_inst : DFF_X1 port map( D => n11372, CK => CLK, Q => 
                           n8861, QN => n24);
   REGISTERS_reg_66_7_inst : DFF_X1 port map( D => n11333, CK => CLK, Q => 
                           n7123, QN => n25);
   REGISTERS_reg_66_6_inst : DFF_X1 port map( D => n11334, CK => CLK, Q => 
                           n7122, QN => n26);
   REGISTERS_reg_66_5_inst : DFF_X1 port map( D => n11335, CK => CLK, Q => 
                           n7120, QN => n27);
   REGISTERS_reg_66_4_inst : DFF_X1 port map( D => n11336, CK => CLK, Q => 
                           n7119, QN => n28);
   REGISTERS_reg_66_3_inst : DFF_X1 port map( D => n11337, CK => CLK, Q => 
                           n7117, QN => n29);
   REGISTERS_reg_66_2_inst : DFF_X1 port map( D => n11338, CK => CLK, Q => 
                           n7116, QN => n30);
   REGISTERS_reg_66_1_inst : DFF_X1 port map( D => n11339, CK => CLK, Q => 
                           n7114, QN => n31);
   REGISTERS_reg_66_0_inst : DFF_X1 port map( D => n11340, CK => CLK, Q => 
                           n7113, QN => n32);
   REGISTERS_reg_65_7_inst : DFF_X1 port map( D => n11301, CK => CLK, Q => 
                           n_1003, QN => n33);
   REGISTERS_reg_65_6_inst : DFF_X1 port map( D => n11302, CK => CLK, Q => 
                           n_1004, QN => n34);
   REGISTERS_reg_65_5_inst : DFF_X1 port map( D => n11303, CK => CLK, Q => 
                           n_1005, QN => n35);
   REGISTERS_reg_65_4_inst : DFF_X1 port map( D => n11304, CK => CLK, Q => 
                           n_1006, QN => n36);
   REGISTERS_reg_65_3_inst : DFF_X1 port map( D => n11305, CK => CLK, Q => 
                           n_1007, QN => n37);
   REGISTERS_reg_65_2_inst : DFF_X1 port map( D => n11306, CK => CLK, Q => 
                           n_1008, QN => n38);
   REGISTERS_reg_65_1_inst : DFF_X1 port map( D => n11307, CK => CLK, Q => 
                           n_1009, QN => n39);
   REGISTERS_reg_65_0_inst : DFF_X1 port map( D => n11308, CK => CLK, Q => 
                           n_1010, QN => n40);
   REGISTERS_reg_64_7_inst : DFF_X1 port map( D => n11269, CK => CLK, Q => 
                           n8823, QN => n41);
   REGISTERS_reg_64_6_inst : DFF_X1 port map( D => n11270, CK => CLK, Q => 
                           n8824, QN => n42);
   REGISTERS_reg_64_5_inst : DFF_X1 port map( D => n11271, CK => CLK, Q => 
                           n8825, QN => n43);
   REGISTERS_reg_64_4_inst : DFF_X1 port map( D => n11272, CK => CLK, Q => 
                           n8826, QN => n44);
   REGISTERS_reg_64_3_inst : DFF_X1 port map( D => n11273, CK => CLK, Q => 
                           n8827, QN => n45);
   REGISTERS_reg_64_2_inst : DFF_X1 port map( D => n11274, CK => CLK, Q => 
                           n8828, QN => n46);
   REGISTERS_reg_64_1_inst : DFF_X1 port map( D => n11275, CK => CLK, Q => 
                           n8829, QN => n47);
   REGISTERS_reg_64_0_inst : DFF_X1 port map( D => n11276, CK => CLK, Q => 
                           n8894, QN => n48);
   REGISTERS_reg_63_7_inst : DFF_X1 port map( D => n11237, CK => CLK, Q => 
                           n8792, QN => n49);
   REGISTERS_reg_63_6_inst : DFF_X1 port map( D => n11238, CK => CLK, Q => 
                           n8793, QN => n50);
   REGISTERS_reg_63_5_inst : DFF_X1 port map( D => n11239, CK => CLK, Q => 
                           n8794, QN => n51);
   REGISTERS_reg_63_4_inst : DFF_X1 port map( D => n11240, CK => CLK, Q => 
                           n8795, QN => n52);
   REGISTERS_reg_63_3_inst : DFF_X1 port map( D => n11241, CK => CLK, Q => 
                           n8796, QN => n53);
   REGISTERS_reg_63_2_inst : DFF_X1 port map( D => n11242, CK => CLK, Q => 
                           n8797, QN => n54);
   REGISTERS_reg_63_1_inst : DFF_X1 port map( D => n11243, CK => CLK, Q => 
                           n8798, QN => n55);
   REGISTERS_reg_63_0_inst : DFF_X1 port map( D => n11244, CK => CLK, Q => 
                           n8895, QN => n56);
   REGISTERS_reg_62_7_inst : DFF_X1 port map( D => n11205, CK => CLK, Q => 
                           n_1011, QN => n1725);
   REGISTERS_reg_62_6_inst : DFF_X1 port map( D => n11206, CK => CLK, Q => 
                           n_1012, QN => n1726);
   REGISTERS_reg_62_5_inst : DFF_X1 port map( D => n11207, CK => CLK, Q => 
                           n_1013, QN => n1727);
   REGISTERS_reg_62_4_inst : DFF_X1 port map( D => n11208, CK => CLK, Q => 
                           n_1014, QN => n1728);
   REGISTERS_reg_62_3_inst : DFF_X1 port map( D => n11209, CK => CLK, Q => 
                           n_1015, QN => n1729);
   REGISTERS_reg_62_2_inst : DFF_X1 port map( D => n11210, CK => CLK, Q => 
                           n_1016, QN => n57);
   REGISTERS_reg_62_1_inst : DFF_X1 port map( D => n11211, CK => CLK, Q => 
                           n_1017, QN => n1730);
   REGISTERS_reg_62_0_inst : DFF_X1 port map( D => n11212, CK => CLK, Q => 
                           n_1018, QN => n1731);
   REGISTERS_reg_61_7_inst : DFF_X1 port map( D => n11173, CK => CLK, Q => 
                           n_1019, QN => n58);
   REGISTERS_reg_61_6_inst : DFF_X1 port map( D => n11174, CK => CLK, Q => 
                           n_1020, QN => n59);
   REGISTERS_reg_61_5_inst : DFF_X1 port map( D => n11175, CK => CLK, Q => 
                           n_1021, QN => n60);
   REGISTERS_reg_61_4_inst : DFF_X1 port map( D => n11176, CK => CLK, Q => 
                           n_1022, QN => n61);
   REGISTERS_reg_61_3_inst : DFF_X1 port map( D => n11177, CK => CLK, Q => 
                           n_1023, QN => n62);
   REGISTERS_reg_61_2_inst : DFF_X1 port map( D => n11178, CK => CLK, Q => 
                           n_1024, QN => n63);
   REGISTERS_reg_61_1_inst : DFF_X1 port map( D => n11179, CK => CLK, Q => 
                           n_1025, QN => n64);
   REGISTERS_reg_61_0_inst : DFF_X1 port map( D => n11180, CK => CLK, Q => 
                           n_1026, QN => n1732);
   REGISTERS_reg_59_7_inst : DFF_X1 port map( D => n11109, CK => CLK, Q => 
                           n8760, QN => n65);
   REGISTERS_reg_59_6_inst : DFF_X1 port map( D => n11110, CK => CLK, Q => 
                           n8761, QN => n66);
   REGISTERS_reg_59_5_inst : DFF_X1 port map( D => n11111, CK => CLK, Q => 
                           n8762, QN => n67);
   REGISTERS_reg_59_4_inst : DFF_X1 port map( D => n11112, CK => CLK, Q => 
                           n8763, QN => n68);
   REGISTERS_reg_59_3_inst : DFF_X1 port map( D => n11113, CK => CLK, Q => 
                           n8764, QN => n69);
   REGISTERS_reg_59_2_inst : DFF_X1 port map( D => n11114, CK => CLK, Q => 
                           n8765, QN => n70);
   REGISTERS_reg_59_1_inst : DFF_X1 port map( D => n11115, CK => CLK, Q => 
                           n8766, QN => n73);
   REGISTERS_reg_59_0_inst : DFF_X1 port map( D => n11116, CK => CLK, Q => 
                           n8767, QN => n74);
   REGISTERS_reg_58_7_inst : DFF_X1 port map( D => n11077, CK => CLK, Q => 
                           n8728, QN => n79);
   REGISTERS_reg_58_6_inst : DFF_X1 port map( D => n11078, CK => CLK, Q => 
                           n8729, QN => n80);
   REGISTERS_reg_58_5_inst : DFF_X1 port map( D => n11079, CK => CLK, Q => 
                           n8730, QN => n85);
   REGISTERS_reg_58_4_inst : DFF_X1 port map( D => n11080, CK => CLK, Q => 
                           n8731, QN => n86);
   REGISTERS_reg_58_3_inst : DFF_X1 port map( D => n11081, CK => CLK, Q => 
                           n8732, QN => n91);
   REGISTERS_reg_58_2_inst : DFF_X1 port map( D => n11082, CK => CLK, Q => 
                           n8733, QN => n92);
   REGISTERS_reg_58_1_inst : DFF_X1 port map( D => n11083, CK => CLK, Q => 
                           n8734, QN => n97);
   REGISTERS_reg_58_0_inst : DFF_X1 port map( D => n11084, CK => CLK, Q => 
                           n8735, QN => n98);
   REGISTERS_reg_57_7_inst : DFF_X1 port map( D => n11045, CK => CLK, Q => 
                           n8696, QN => n100);
   REGISTERS_reg_57_6_inst : DFF_X1 port map( D => n11046, CK => CLK, Q => 
                           n8697, QN => n101);
   REGISTERS_reg_57_5_inst : DFF_X1 port map( D => n11047, CK => CLK, Q => 
                           n8698, QN => n102);
   REGISTERS_reg_57_4_inst : DFF_X1 port map( D => n11048, CK => CLK, Q => 
                           n8699, QN => n103);
   REGISTERS_reg_57_3_inst : DFF_X1 port map( D => n11049, CK => CLK, Q => 
                           n8700, QN => n104);
   REGISTERS_reg_57_2_inst : DFF_X1 port map( D => n11050, CK => CLK, Q => 
                           n8701, QN => n105);
   REGISTERS_reg_57_1_inst : DFF_X1 port map( D => n11051, CK => CLK, Q => 
                           n8702, QN => n106);
   REGISTERS_reg_57_0_inst : DFF_X1 port map( D => n11052, CK => CLK, Q => 
                           n8703, QN => n107);
   REGISTERS_reg_56_7_inst : DFF_X1 port map( D => n11013, CK => CLK, Q => 
                           n8664, QN => n108);
   REGISTERS_reg_56_6_inst : DFF_X1 port map( D => n11014, CK => CLK, Q => 
                           n8665, QN => n109);
   REGISTERS_reg_56_5_inst : DFF_X1 port map( D => n11015, CK => CLK, Q => 
                           n8666, QN => n110);
   REGISTERS_reg_56_4_inst : DFF_X1 port map( D => n11016, CK => CLK, Q => 
                           n8667, QN => n111);
   REGISTERS_reg_56_3_inst : DFF_X1 port map( D => n11017, CK => CLK, Q => 
                           n8668, QN => n112);
   REGISTERS_reg_56_2_inst : DFF_X1 port map( D => n11018, CK => CLK, Q => 
                           n8669, QN => n113);
   REGISTERS_reg_56_1_inst : DFF_X1 port map( D => n11019, CK => CLK, Q => 
                           n8670, QN => n114);
   REGISTERS_reg_56_0_inst : DFF_X1 port map( D => n11020, CK => CLK, Q => 
                           n8671, QN => n115);
   REGISTERS_reg_55_7_inst : DFF_X1 port map( D => n10981, CK => CLK, Q => 
                           n7499, QN => n116);
   REGISTERS_reg_55_6_inst : DFF_X1 port map( D => n10982, CK => CLK, Q => 
                           n7497, QN => n117);
   REGISTERS_reg_55_5_inst : DFF_X1 port map( D => n10983, CK => CLK, Q => 
                           n7495, QN => n118);
   REGISTERS_reg_55_4_inst : DFF_X1 port map( D => n10984, CK => CLK, Q => 
                           n7494, QN => n119);
   REGISTERS_reg_55_3_inst : DFF_X1 port map( D => n10985, CK => CLK, Q => 
                           n7493, QN => n120);
   REGISTERS_reg_55_2_inst : DFF_X1 port map( D => n10986, CK => CLK, Q => 
                           n7492, QN => n121);
   REGISTERS_reg_55_1_inst : DFF_X1 port map( D => n10987, CK => CLK, Q => 
                           n7491, QN => n122);
   REGISTERS_reg_55_0_inst : DFF_X1 port map( D => n10988, CK => CLK, Q => 
                           n7469, QN => n123);
   REGISTERS_reg_54_7_inst : DFF_X1 port map( D => n10949, CK => CLK, Q => 
                           n_1027, QN => n124);
   REGISTERS_reg_54_6_inst : DFF_X1 port map( D => n10950, CK => CLK, Q => 
                           n_1028, QN => n125);
   REGISTERS_reg_54_5_inst : DFF_X1 port map( D => n10951, CK => CLK, Q => 
                           n_1029, QN => n126);
   REGISTERS_reg_54_4_inst : DFF_X1 port map( D => n10952, CK => CLK, Q => 
                           n_1030, QN => n127);
   REGISTERS_reg_54_3_inst : DFF_X1 port map( D => n10953, CK => CLK, Q => 
                           n_1031, QN => n128);
   REGISTERS_reg_54_2_inst : DFF_X1 port map( D => n10954, CK => CLK, Q => 
                           n_1032, QN => n129);
   REGISTERS_reg_54_1_inst : DFF_X1 port map( D => n10955, CK => CLK, Q => 
                           n_1033, QN => n130);
   REGISTERS_reg_54_0_inst : DFF_X1 port map( D => n10956, CK => CLK, Q => 
                           n_1034, QN => n131);
   REGISTERS_reg_53_2_inst : DFF_X1 port map( D => n10922, CK => CLK, Q => 
                           n_1035, QN => n132);
   REGISTERS_reg_53_0_inst : DFF_X1 port map( D => n10924, CK => CLK, Q => 
                           n_1036, QN => n1741);
   REGISTERS_reg_52_7_inst : DFF_X1 port map( D => n10885, CK => CLK, Q => 
                           n_1037, QN => n133);
   REGISTERS_reg_52_6_inst : DFF_X1 port map( D => n10886, CK => CLK, Q => 
                           n_1038, QN => n134);
   REGISTERS_reg_52_5_inst : DFF_X1 port map( D => n10887, CK => CLK, Q => 
                           n_1039, QN => n135);
   REGISTERS_reg_52_4_inst : DFF_X1 port map( D => n10888, CK => CLK, Q => 
                           n_1040, QN => n136);
   REGISTERS_reg_52_3_inst : DFF_X1 port map( D => n10889, CK => CLK, Q => 
                           n_1041, QN => n137);
   REGISTERS_reg_52_2_inst : DFF_X1 port map( D => n10890, CK => CLK, Q => 
                           n_1042, QN => n138);
   REGISTERS_reg_52_1_inst : DFF_X1 port map( D => n10891, CK => CLK, Q => 
                           n_1043, QN => n139);
   REGISTERS_reg_52_0_inst : DFF_X1 port map( D => n10892, CK => CLK, Q => 
                           n_1044, QN => n1742);
   REGISTERS_reg_50_7_inst : DFF_X1 port map( D => n10821, CK => CLK, Q => 
                           n8632, QN => n140);
   REGISTERS_reg_50_6_inst : DFF_X1 port map( D => n10822, CK => CLK, Q => 
                           n8633, QN => n141);
   REGISTERS_reg_50_5_inst : DFF_X1 port map( D => n10823, CK => CLK, Q => 
                           n8634, QN => n142);
   REGISTERS_reg_50_4_inst : DFF_X1 port map( D => n10824, CK => CLK, Q => 
                           n8635, QN => n143);
   REGISTERS_reg_50_3_inst : DFF_X1 port map( D => n10825, CK => CLK, Q => 
                           n8636, QN => n144);
   REGISTERS_reg_50_2_inst : DFF_X1 port map( D => n10826, CK => CLK, Q => 
                           n8637, QN => n145);
   REGISTERS_reg_50_1_inst : DFF_X1 port map( D => n10827, CK => CLK, Q => 
                           n8638, QN => n146);
   REGISTERS_reg_50_0_inst : DFF_X1 port map( D => n10828, CK => CLK, Q => 
                           n8639, QN => n147);
   REGISTERS_reg_49_7_inst : DFF_X1 port map( D => n10789, CK => CLK, Q => 
                           n8600, QN => n148);
   REGISTERS_reg_49_6_inst : DFF_X1 port map( D => n10790, CK => CLK, Q => 
                           n8601, QN => n149);
   REGISTERS_reg_49_5_inst : DFF_X1 port map( D => n10791, CK => CLK, Q => 
                           n8602, QN => n150);
   REGISTERS_reg_49_4_inst : DFF_X1 port map( D => n10792, CK => CLK, Q => 
                           n8603, QN => n151);
   REGISTERS_reg_49_3_inst : DFF_X1 port map( D => n10793, CK => CLK, Q => 
                           n8604, QN => n152);
   REGISTERS_reg_49_2_inst : DFF_X1 port map( D => n10794, CK => CLK, Q => 
                           n8605, QN => n153);
   REGISTERS_reg_49_1_inst : DFF_X1 port map( D => n10795, CK => CLK, Q => 
                           n8606, QN => n154);
   REGISTERS_reg_49_0_inst : DFF_X1 port map( D => n10796, CK => CLK, Q => 
                           n8607, QN => n155);
   REGISTERS_reg_48_7_inst : DFF_X1 port map( D => n10757, CK => CLK, Q => 
                           n_1045, QN => n156);
   REGISTERS_reg_48_6_inst : DFF_X1 port map( D => n10758, CK => CLK, Q => 
                           n_1046, QN => n157);
   REGISTERS_reg_48_5_inst : DFF_X1 port map( D => n10759, CK => CLK, Q => 
                           n_1047, QN => n158);
   REGISTERS_reg_48_4_inst : DFF_X1 port map( D => n10760, CK => CLK, Q => 
                           n_1048, QN => n159);
   REGISTERS_reg_48_3_inst : DFF_X1 port map( D => n10761, CK => CLK, Q => 
                           n_1049, QN => n160);
   REGISTERS_reg_48_2_inst : DFF_X1 port map( D => n10762, CK => CLK, Q => 
                           n_1050, QN => n161);
   REGISTERS_reg_48_1_inst : DFF_X1 port map( D => n10763, CK => CLK, Q => 
                           n_1051, QN => n162);
   REGISTERS_reg_48_0_inst : DFF_X1 port map( D => n10764, CK => CLK, Q => 
                           n_1052, QN => n163);
   REGISTERS_reg_47_7_inst : DFF_X1 port map( D => n10725, CK => CLK, Q => 
                           n_1053, QN => n164);
   REGISTERS_reg_47_6_inst : DFF_X1 port map( D => n10726, CK => CLK, Q => 
                           n_1054, QN => n165);
   REGISTERS_reg_47_5_inst : DFF_X1 port map( D => n10727, CK => CLK, Q => 
                           n_1055, QN => n166);
   REGISTERS_reg_47_4_inst : DFF_X1 port map( D => n10728, CK => CLK, Q => 
                           n_1056, QN => n167);
   REGISTERS_reg_47_3_inst : DFF_X1 port map( D => n10729, CK => CLK, Q => 
                           n_1057, QN => n168);
   REGISTERS_reg_47_2_inst : DFF_X1 port map( D => n10730, CK => CLK, Q => 
                           n_1058, QN => n169);
   REGISTERS_reg_47_1_inst : DFF_X1 port map( D => n10731, CK => CLK, Q => 
                           n_1059, QN => n170);
   REGISTERS_reg_47_0_inst : DFF_X1 port map( D => n10732, CK => CLK, Q => 
                           n_1060, QN => n171);
   REGISTERS_reg_46_7_inst : DFF_X1 port map( D => n10693, CK => CLK, Q => 
                           n8506, QN => n172);
   REGISTERS_reg_46_6_inst : DFF_X1 port map( D => n10694, CK => CLK, Q => 
                           n8507, QN => n173);
   REGISTERS_reg_46_5_inst : DFF_X1 port map( D => n10695, CK => CLK, Q => 
                           n8508, QN => n174);
   REGISTERS_reg_46_4_inst : DFF_X1 port map( D => n10696, CK => CLK, Q => 
                           n8509, QN => n175);
   REGISTERS_reg_46_3_inst : DFF_X1 port map( D => n10697, CK => CLK, Q => 
                           n8510, QN => n176);
   REGISTERS_reg_46_2_inst : DFF_X1 port map( D => n10698, CK => CLK, Q => 
                           n8511, QN => n177);
   REGISTERS_reg_46_1_inst : DFF_X1 port map( D => n10699, CK => CLK, Q => 
                           n8512, QN => n178);
   REGISTERS_reg_46_0_inst : DFF_X1 port map( D => n10700, CK => CLK, Q => 
                           n8513, QN => n179);
   REGISTERS_reg_45_7_inst : DFF_X1 port map( D => n10661, CK => CLK, Q => 
                           n8474, QN => n180);
   REGISTERS_reg_45_6_inst : DFF_X1 port map( D => n10662, CK => CLK, Q => 
                           n8475, QN => n181);
   REGISTERS_reg_45_5_inst : DFF_X1 port map( D => n10663, CK => CLK, Q => 
                           n8476, QN => n182);
   REGISTERS_reg_45_4_inst : DFF_X1 port map( D => n10664, CK => CLK, Q => 
                           n8477, QN => n183);
   REGISTERS_reg_45_3_inst : DFF_X1 port map( D => n10665, CK => CLK, Q => 
                           n8478, QN => n184);
   REGISTERS_reg_45_2_inst : DFF_X1 port map( D => n10666, CK => CLK, Q => 
                           n8479, QN => n185);
   REGISTERS_reg_45_1_inst : DFF_X1 port map( D => n10667, CK => CLK, Q => 
                           n8480, QN => n186);
   REGISTERS_reg_45_0_inst : DFF_X1 port map( D => n10668, CK => CLK, Q => 
                           n8481, QN => n187);
   REGISTERS_reg_44_7_inst : DFF_X1 port map( D => n10629, CK => CLK, Q => 
                           n_1061, QN => n1751);
   REGISTERS_reg_44_6_inst : DFF_X1 port map( D => n10630, CK => CLK, Q => 
                           n_1062, QN => n1752);
   REGISTERS_reg_44_5_inst : DFF_X1 port map( D => n10631, CK => CLK, Q => 
                           n_1063, QN => n1753);
   REGISTERS_reg_44_4_inst : DFF_X1 port map( D => n10632, CK => CLK, Q => 
                           n_1064, QN => n1754);
   REGISTERS_reg_44_3_inst : DFF_X1 port map( D => n10633, CK => CLK, Q => 
                           n_1065, QN => n1755);
   REGISTERS_reg_44_2_inst : DFF_X1 port map( D => n10634, CK => CLK, Q => 
                           n_1066, QN => n188);
   REGISTERS_reg_44_1_inst : DFF_X1 port map( D => n10635, CK => CLK, Q => 
                           n_1067, QN => n1756);
   REGISTERS_reg_44_0_inst : DFF_X1 port map( D => n10636, CK => CLK, Q => 
                           n_1068, QN => n1757);
   REGISTERS_reg_43_7_inst : DFF_X1 port map( D => n10597, CK => CLK, Q => 
                           n_1069, QN => n189);
   REGISTERS_reg_43_6_inst : DFF_X1 port map( D => n10598, CK => CLK, Q => 
                           n_1070, QN => n190);
   REGISTERS_reg_43_5_inst : DFF_X1 port map( D => n10599, CK => CLK, Q => 
                           n_1071, QN => n191);
   REGISTERS_reg_43_4_inst : DFF_X1 port map( D => n10600, CK => CLK, Q => 
                           n_1072, QN => n192);
   REGISTERS_reg_43_3_inst : DFF_X1 port map( D => n10601, CK => CLK, Q => 
                           n_1073, QN => n193);
   REGISTERS_reg_43_2_inst : DFF_X1 port map( D => n10602, CK => CLK, Q => 
                           n_1074, QN => n194);
   REGISTERS_reg_43_1_inst : DFF_X1 port map( D => n10603, CK => CLK, Q => 
                           n_1075, QN => n195);
   REGISTERS_reg_43_0_inst : DFF_X1 port map( D => n10604, CK => CLK, Q => 
                           n_1076, QN => n1758);
   REGISTERS_reg_41_7_inst : DFF_X1 port map( D => n10533, CK => CLK, Q => 
                           n8442, QN => n196);
   REGISTERS_reg_41_6_inst : DFF_X1 port map( D => n10534, CK => CLK, Q => 
                           n8443, QN => n197);
   REGISTERS_reg_41_5_inst : DFF_X1 port map( D => n10535, CK => CLK, Q => 
                           n8444, QN => n198);
   REGISTERS_reg_41_4_inst : DFF_X1 port map( D => n10536, CK => CLK, Q => 
                           n8445, QN => n199);
   REGISTERS_reg_41_3_inst : DFF_X1 port map( D => n10537, CK => CLK, Q => 
                           n8446, QN => n200);
   REGISTERS_reg_41_2_inst : DFF_X1 port map( D => n10538, CK => CLK, Q => 
                           n8447, QN => n201);
   REGISTERS_reg_41_1_inst : DFF_X1 port map( D => n10539, CK => CLK, Q => 
                           n8448, QN => n202);
   REGISTERS_reg_41_0_inst : DFF_X1 port map( D => n10540, CK => CLK, Q => 
                           n8449, QN => n203);
   REGISTERS_reg_40_7_inst : DFF_X1 port map( D => n10501, CK => CLK, Q => 
                           n8410, QN => n204);
   REGISTERS_reg_40_6_inst : DFF_X1 port map( D => n10502, CK => CLK, Q => 
                           n8411, QN => n205);
   REGISTERS_reg_40_5_inst : DFF_X1 port map( D => n10503, CK => CLK, Q => 
                           n8412, QN => n206);
   REGISTERS_reg_40_4_inst : DFF_X1 port map( D => n10504, CK => CLK, Q => 
                           n8413, QN => n207);
   REGISTERS_reg_40_3_inst : DFF_X1 port map( D => n10505, CK => CLK, Q => 
                           n8414, QN => n208);
   REGISTERS_reg_40_2_inst : DFF_X1 port map( D => n10506, CK => CLK, Q => 
                           n8415, QN => n209);
   REGISTERS_reg_40_1_inst : DFF_X1 port map( D => n10507, CK => CLK, Q => 
                           n8416, QN => n210);
   REGISTERS_reg_40_0_inst : DFF_X1 port map( D => n10508, CK => CLK, Q => 
                           n8417, QN => n211);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n10476, CK => CLK, Q => n830
                           , QN => n212);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n10405, CK => CLK, Q => 
                           n_1077, QN => n213);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n10406, CK => CLK, Q => 
                           n_1078, QN => n214);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n10407, CK => CLK, Q => 
                           n_1079, QN => n215);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n10408, CK => CLK, Q => 
                           n_1080, QN => n216);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n10409, CK => CLK, Q => 
                           n_1081, QN => n217);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n10410, CK => CLK, Q => 
                           n_1082, QN => n218);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n10411, CK => CLK, Q => 
                           n_1083, QN => n219);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n10412, CK => CLK, Q => 
                           n8385, QN => n220);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n10373, CK => CLK, Q => 
                           n_1084, QN => n221);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n10374, CK => CLK, Q => 
                           n_1085, QN => n222);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n10375, CK => CLK, Q => 
                           n_1086, QN => n223);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n10376, CK => CLK, Q => 
                           n_1087, QN => n224);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n10377, CK => CLK, Q => 
                           n_1088, QN => n225);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n10378, CK => CLK, Q => 
                           n_1089, QN => n226);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n10379, CK => CLK, Q => 
                           n_1090, QN => n227);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n10380, CK => CLK, Q => 
                           n8353, QN => n228);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n10348, CK => CLK, Q => 
                           n_1091, QN => n1782);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n10309, CK => CLK, Q => 
                           n_1092, QN => n229);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n10310, CK => CLK, Q => 
                           n_1093, QN => n230);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n10311, CK => CLK, Q => 
                           n_1094, QN => n231);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n10312, CK => CLK, Q => 
                           n_1095, QN => n232);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n10313, CK => CLK, Q => 
                           n_1096, QN => n233);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n10314, CK => CLK, Q => 
                           n_1097, QN => n234);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n10315, CK => CLK, Q => 
                           n_1098, QN => n235);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n10316, CK => CLK, Q => 
                           n_1099, QN => n1783);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n10245, CK => CLK, Q => 
                           n8314, QN => n236);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n10246, CK => CLK, Q => 
                           n8315, QN => n237);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n10247, CK => CLK, Q => 
                           n8316, QN => n238);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n10248, CK => CLK, Q => 
                           n8317, QN => n239);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n10249, CK => CLK, Q => 
                           n8318, QN => n240);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n10250, CK => CLK, Q => 
                           n8319, QN => n241);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n10251, CK => CLK, Q => 
                           n8320, QN => n242);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n10252, CK => CLK, Q => 
                           n8321, QN => n243);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n10213, CK => CLK, Q => 
                           n8282, QN => n244);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n10214, CK => CLK, Q => 
                           n8283, QN => n245);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n10215, CK => CLK, Q => 
                           n8284, QN => n246);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n10216, CK => CLK, Q => 
                           n8285, QN => n247);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n10217, CK => CLK, Q => 
                           n8286, QN => n248);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n10218, CK => CLK, Q => 
                           n8287, QN => n249);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n10219, CK => CLK, Q => 
                           n8288, QN => n250);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n10220, CK => CLK, Q => 
                           n8289, QN => n251);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n10188, CK => CLK, Q => n896
                           , QN => n252);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n10117, CK => CLK, Q => 
                           n_1100, QN => n253);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n10118, CK => CLK, Q => 
                           n_1101, QN => n254);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n10119, CK => CLK, Q => 
                           n_1102, QN => n255);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n10120, CK => CLK, Q => 
                           n_1103, QN => n256);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n10121, CK => CLK, Q => 
                           n_1104, QN => n257);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n10122, CK => CLK, Q => 
                           n_1105, QN => n258);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n10123, CK => CLK, Q => 
                           n_1106, QN => n259);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n10124, CK => CLK, Q => 
                           n_1107, QN => n260);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n10085, CK => CLK, Q => 
                           n_1108, QN => n261);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n10086, CK => CLK, Q => 
                           n_1109, QN => n262);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n10087, CK => CLK, Q => 
                           n_1110, QN => n263);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n10088, CK => CLK, Q => 
                           n_1111, QN => n264);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n10089, CK => CLK, Q => 
                           n_1112, QN => n265);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n10090, CK => CLK, Q => 
                           n_1113, QN => n266);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n10091, CK => CLK, Q => 
                           n_1114, QN => n267);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n10092, CK => CLK, Q => 
                           n_1115, QN => n268);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n9669, CK => CLK, Q => n8124
                           , QN => n269);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n9670, CK => CLK, Q => n8125
                           , QN => n270);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n9671, CK => CLK, Q => n8126
                           , QN => n271);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n9672, CK => CLK, Q => n8127
                           , QN => n272);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n9673, CK => CLK, Q => n8128
                           , QN => n273);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n9674, CK => CLK, Q => n8129
                           , QN => n274);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n9675, CK => CLK, Q => n8130
                           , QN => n275);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n9676, CK => CLK, Q => n8131
                           , QN => n276);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n9637, CK => CLK, Q => n8092
                           , QN => n277);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n9638, CK => CLK, Q => n8093
                           , QN => n278);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n9639, CK => CLK, Q => n8094
                           , QN => n279);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n9640, CK => CLK, Q => n8095
                           , QN => n280);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n9641, CK => CLK, Q => n8096
                           , QN => n281);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n9642, CK => CLK, Q => n8097
                           , QN => n282);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n9643, CK => CLK, Q => n8098
                           , QN => n283);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n9644, CK => CLK, Q => n8099
                           , QN => n284);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n9605, CK => CLK, Q => n846,
                           QN => n285);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n9606, CK => CLK, Q => n844,
                           QN => n286);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n9607, CK => CLK, Q => n842,
                           QN => n287);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n9608, CK => CLK, Q => n840,
                           QN => n288);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n9609, CK => CLK, Q => n838,
                           QN => n289);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n9610, CK => CLK, Q => n836,
                           QN => n290);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n9611, CK => CLK, Q => n834,
                           QN => n291);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n9612, CK => CLK, Q => n832,
                           QN => n292);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n9541, CK => CLK, Q => n8060
                           , QN => n293);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n9542, CK => CLK, Q => n8061
                           , QN => n294);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n9543, CK => CLK, Q => n8062
                           , QN => n295);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n9544, CK => CLK, Q => n8063
                           , QN => n296);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n9545, CK => CLK, Q => n8064
                           , QN => n297);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n9546, CK => CLK, Q => n8065
                           , QN => n298);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n9547, CK => CLK, Q => n8066
                           , QN => n299);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n9548, CK => CLK, Q => n8067
                           , QN => n300);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n9509, CK => CLK, Q => n8028,
                           QN => n301);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n9510, CK => CLK, Q => n8029,
                           QN => n302);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n9511, CK => CLK, Q => n8030,
                           QN => n303);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n9512, CK => CLK, Q => n8031,
                           QN => n304);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n9513, CK => CLK, Q => n8032,
                           QN => n305);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n9514, CK => CLK, Q => n8033,
                           QN => n306);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n9515, CK => CLK, Q => n8034,
                           QN => n307);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n9516, CK => CLK, Q => n8035,
                           QN => n308);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n9477, CK => CLK, Q => n_1116
                           , QN => n309);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n9478, CK => CLK, Q => n_1117
                           , QN => n310);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n9479, CK => CLK, Q => n_1118
                           , QN => n311);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n9480, CK => CLK, Q => n_1119
                           , QN => n312);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n9481, CK => CLK, Q => n_1120
                           , QN => n313);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n9482, CK => CLK, Q => n_1121
                           , QN => n314);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n9483, CK => CLK, Q => n_1122
                           , QN => n315);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n9484, CK => CLK, Q => n_1123
                           , QN => n316);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n9445, CK => CLK, Q => n_1124
                           , QN => n317);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n9446, CK => CLK, Q => n_1125
                           , QN => n318);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n9447, CK => CLK, Q => n_1126
                           , QN => n319);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n9448, CK => CLK, Q => n_1127
                           , QN => n320);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n9449, CK => CLK, Q => n_1128
                           , QN => n321);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n9450, CK => CLK, Q => n_1129
                           , QN => n322);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n9451, CK => CLK, Q => n_1130
                           , QN => n323);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n9452, CK => CLK, Q => n_1131
                           , QN => n324);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n9413, CK => CLK, Q => n6826,
                           QN => n325);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n9414, CK => CLK, Q => n6817,
                           QN => n326);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n9415, CK => CLK, Q => n6799,
                           QN => n327);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n9416, CK => CLK, Q => n6787,
                           QN => n328);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n9417, CK => CLK, Q => n6778,
                           QN => n329);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n9418, CK => CLK, Q => n6771,
                           QN => n330);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n9419, CK => CLK, Q => n6754,
                           QN => n331);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n9420, CK => CLK, Q => n7108,
                           QN => n332);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n9381, CK => CLK, Q => n7996,
                           QN => n333);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n9382, CK => CLK, Q => n7997,
                           QN => n334);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n9383, CK => CLK, Q => n7998,
                           QN => n335);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n9384, CK => CLK, Q => n7999,
                           QN => n336);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n9385, CK => CLK, Q => n8000,
                           QN => n337);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n9386, CK => CLK, Q => n8001,
                           QN => n338);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n9387, CK => CLK, Q => n8002,
                           QN => n339);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n9388, CK => CLK, Q => n8003,
                           QN => n340);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n9349, CK => CLK, Q => n7964,
                           QN => n341);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n9350, CK => CLK, Q => n7965,
                           QN => n342);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n9351, CK => CLK, Q => n7966,
                           QN => n343);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n9352, CK => CLK, Q => n7967,
                           QN => n344);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n9353, CK => CLK, Q => n7968,
                           QN => n345);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n9354, CK => CLK, Q => n7969,
                           QN => n346);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n9355, CK => CLK, Q => n7970,
                           QN => n347);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n9356, CK => CLK, Q => n7971,
                           QN => n348);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n9317, CK => CLK, Q => n847, 
                           QN => n349);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n9318, CK => CLK, Q => n845, 
                           QN => n350);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n9319, CK => CLK, Q => n843, 
                           QN => n351);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n9320, CK => CLK, Q => n841, 
                           QN => n352);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n9321, CK => CLK, Q => n839, 
                           QN => n353);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n9322, CK => CLK, Q => n837, 
                           QN => n354);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n9323, CK => CLK, Q => n835, 
                           QN => n355);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n9324, CK => CLK, Q => n833, 
                           QN => n356);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n9253, CK => CLK, Q => n7932,
                           QN => n357);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n9254, CK => CLK, Q => n7933,
                           QN => n358);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n9255, CK => CLK, Q => n7934,
                           QN => n359);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n9256, CK => CLK, Q => n7935,
                           QN => n360);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n9257, CK => CLK, Q => n7936,
                           QN => n361);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n9258, CK => CLK, Q => n7937,
                           QN => n362);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n9259, CK => CLK, Q => n7938,
                           QN => n363);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n9260, CK => CLK, Q => n7939,
                           QN => n364);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n9215, CK => CLK, Q => n7888,
                           QN => n365);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n9217, CK => CLK, Q => n7891,
                           QN => n366);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n9219, CK => CLK, Q => n7894,
                           QN => n367);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n9221, CK => CLK, Q => n7897,
                           QN => n368);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n9223, CK => CLK, Q => n7900,
                           QN => n369);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n9225, CK => CLK, Q => n7903,
                           QN => n370);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n9227, CK => CLK, Q => n7906,
                           QN => n371);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n9228, CK => CLK, Q => n7907,
                           QN => n372);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n9957, CK => CLK, Q => n8188
                           , QN => n373);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n9958, CK => CLK, Q => n8189
                           , QN => n374);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n9959, CK => CLK, Q => n8190
                           , QN => n375);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n9960, CK => CLK, Q => n8191
                           , QN => n376);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n9961, CK => CLK, Q => n8192
                           , QN => n377);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n9962, CK => CLK, Q => n8193
                           , QN => n378);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n9963, CK => CLK, Q => n8194
                           , QN => n379);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n9964, CK => CLK, Q => n8195
                           , QN => n380);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n9925, CK => CLK, Q => n8156
                           , QN => n381);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n9926, CK => CLK, Q => n8157
                           , QN => n382);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n9927, CK => CLK, Q => n8158
                           , QN => n383);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n9928, CK => CLK, Q => n8159
                           , QN => n384);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n9929, CK => CLK, Q => n8160
                           , QN => n385);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n9930, CK => CLK, Q => n8161
                           , QN => n386);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n9931, CK => CLK, Q => n8162
                           , QN => n387);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n9932, CK => CLK, Q => n8163
                           , QN => n388);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n9829, CK => CLK, Q => n6832
                           , QN => n389);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n9830, CK => CLK, Q => n6820
                           , QN => n390);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n9831, CK => CLK, Q => n6805
                           , QN => n391);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n9832, CK => CLK, Q => n6795
                           , QN => n392);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n9833, CK => CLK, Q => n6781
                           , QN => n393);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n9834, CK => CLK, Q => n6773
                           , QN => n394);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n9835, CK => CLK, Q => n6760
                           , QN => n395);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n9836, CK => CLK, Q => n7107
                           , QN => n396);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n9797, CK => CLK, Q => 
                           n_1132, QN => n397);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n9798, CK => CLK, Q => 
                           n_1133, QN => n398);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n9799, CK => CLK, Q => 
                           n_1134, QN => n399);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n9800, CK => CLK, Q => 
                           n_1135, QN => n400);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n9801, CK => CLK, Q => 
                           n_1136, QN => n401);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n9802, CK => CLK, Q => 
                           n_1137, QN => n402);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n9803, CK => CLK, Q => 
                           n_1138, QN => n403);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n9804, CK => CLK, Q => 
                           n_1139, QN => n404);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n9733, CK => CLK, Q => 
                           n_1140, QN => n405);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n9734, CK => CLK, Q => 
                           n_1141, QN => n406);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n9735, CK => CLK, Q => 
                           n_1142, QN => n407);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n9736, CK => CLK, Q => 
                           n_1143, QN => n408);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n9737, CK => CLK, Q => 
                           n_1144, QN => n409);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n9738, CK => CLK, Q => 
                           n_1145, QN => n410);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n9739, CK => CLK, Q => 
                           n_1146, QN => n411);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n9645, CK => CLK, Q => 
                           n8100, QN => n412);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n9646, CK => CLK, Q => 
                           n8101, QN => n413);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n9647, CK => CLK, Q => 
                           n8102, QN => n414);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n9649, CK => CLK, Q => 
                           n8104, QN => n416);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n9650, CK => CLK, Q => 
                           n8105, QN => n417);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n9651, CK => CLK, Q => 
                           n8106, QN => n418);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n9652, CK => CLK, Q => 
                           n8107, QN => n419);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n9653, CK => CLK, Q => 
                           n8108, QN => n420);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n9654, CK => CLK, Q => 
                           n8109, QN => n421);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n9655, CK => CLK, Q => 
                           n8110, QN => n422);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n9656, CK => CLK, Q => 
                           n8111, QN => n423);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n9658, CK => CLK, Q => 
                           n8113, QN => n425);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n9659, CK => CLK, Q => 
                           n8114, QN => n426);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n9660, CK => CLK, Q => 
                           n8115, QN => n427);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n9661, CK => CLK, Q => 
                           n8116, QN => n428);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n9662, CK => CLK, Q => 
                           n8117, QN => n429);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n9663, CK => CLK, Q => 
                           n8118, QN => n430);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n9664, CK => CLK, Q => 
                           n8119, QN => n431);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n9665, CK => CLK, Q => 
                           n8120, QN => n432);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n9666, CK => CLK, Q => 
                           n8121, QN => n433);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n9667, CK => CLK, Q => n8122
                           , QN => n434);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n9668, CK => CLK, Q => n8123
                           , QN => n435);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n9613, CK => CLK, Q => 
                           n8068, QN => n436);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n9614, CK => CLK, Q => 
                           n8069, QN => n437);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n9615, CK => CLK, Q => 
                           n8070, QN => n438);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n9616, CK => CLK, Q => 
                           n8071, QN => n439);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n9617, CK => CLK, Q => 
                           n8072, QN => n440);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n9618, CK => CLK, Q => 
                           n8073, QN => n441);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n9619, CK => CLK, Q => 
                           n8074, QN => n442);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n9620, CK => CLK, Q => 
                           n8075, QN => n443);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n9621, CK => CLK, Q => 
                           n8076, QN => n444);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n9622, CK => CLK, Q => 
                           n8077, QN => n445);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n9623, CK => CLK, Q => 
                           n8078, QN => n446);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n9624, CK => CLK, Q => 
                           n8079, QN => n447);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n9626, CK => CLK, Q => 
                           n8081, QN => n449);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n9627, CK => CLK, Q => 
                           n8082, QN => n450);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n9628, CK => CLK, Q => 
                           n8083, QN => n451);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n9629, CK => CLK, Q => 
                           n8084, QN => n452);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n9630, CK => CLK, Q => 
                           n8085, QN => n453);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n9631, CK => CLK, Q => 
                           n8086, QN => n454);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n9632, CK => CLK, Q => 
                           n8087, QN => n455);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n9633, CK => CLK, Q => 
                           n8088, QN => n456);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n9634, CK => CLK, Q => 
                           n8089, QN => n457);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n9635, CK => CLK, Q => n8090
                           , QN => n458);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n9636, CK => CLK, Q => n8091
                           , QN => n459);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n9581, CK => CLK, Q => n894
                           , QN => n460);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n9582, CK => CLK, Q => n892
                           , QN => n461);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n9583, CK => CLK, Q => n890
                           , QN => n462);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n9584, CK => CLK, Q => n888
                           , QN => n463);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n9585, CK => CLK, Q => n886
                           , QN => n464);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n9586, CK => CLK, Q => n884
                           , QN => n465);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n9587, CK => CLK, Q => n882
                           , QN => n466);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n9588, CK => CLK, Q => n880
                           , QN => n467);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n9589, CK => CLK, Q => n878
                           , QN => n468);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n9590, CK => CLK, Q => n876
                           , QN => n469);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n9591, CK => CLK, Q => n874
                           , QN => n470);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n9592, CK => CLK, Q => n872
                           , QN => n471);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n9593, CK => CLK, Q => n870
                           , QN => n472);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n9594, CK => CLK, Q => n868
                           , QN => n473);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n9595, CK => CLK, Q => n866
                           , QN => n474);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n9596, CK => CLK, Q => n864
                           , QN => n475);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n9597, CK => CLK, Q => n862
                           , QN => n476);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n9598, CK => CLK, Q => n860
                           , QN => n477);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n9599, CK => CLK, Q => n858
                           , QN => n478);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n9600, CK => CLK, Q => n856
                           , QN => n479);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n9601, CK => CLK, Q => n854
                           , QN => n480);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n9602, CK => CLK, Q => n852
                           , QN => n481);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n9603, CK => CLK, Q => n850,
                           QN => n482);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n9604, CK => CLK, Q => n848,
                           QN => n483);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n9561, CK => CLK, Q => n812
                           , QN => n1868);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n9517, CK => CLK, Q => 
                           n8036, QN => n484);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n9518, CK => CLK, Q => 
                           n8037, QN => n485);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n9519, CK => CLK, Q => 
                           n8038, QN => n486);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n9520, CK => CLK, Q => 
                           n8039, QN => n487);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n9521, CK => CLK, Q => 
                           n8040, QN => n488);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n9522, CK => CLK, Q => 
                           n8041, QN => n489);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n9523, CK => CLK, Q => 
                           n8042, QN => n490);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n9524, CK => CLK, Q => 
                           n8043, QN => n491);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n9525, CK => CLK, Q => 
                           n8044, QN => n492);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n9526, CK => CLK, Q => 
                           n8045, QN => n493);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n9527, CK => CLK, Q => 
                           n8046, QN => n494);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n9528, CK => CLK, Q => 
                           n8047, QN => n495);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n9530, CK => CLK, Q => 
                           n8049, QN => n497);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n9531, CK => CLK, Q => 
                           n8050, QN => n498);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n9532, CK => CLK, Q => 
                           n8051, QN => n499);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n9533, CK => CLK, Q => 
                           n8052, QN => n500);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n9534, CK => CLK, Q => 
                           n8053, QN => n501);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n9535, CK => CLK, Q => 
                           n8054, QN => n502);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n9536, CK => CLK, Q => 
                           n8055, QN => n503);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n9537, CK => CLK, Q => 
                           n8056, QN => n504);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n9538, CK => CLK, Q => 
                           n8057, QN => n505);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n9539, CK => CLK, Q => n8058
                           , QN => n506);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n9540, CK => CLK, Q => n8059
                           , QN => n507);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n9421, CK => CLK, Q => 
                           n_1147, QN => n508);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n9422, CK => CLK, Q => 
                           n_1148, QN => n509);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n9423, CK => CLK, Q => 
                           n_1149, QN => n510);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n9424, CK => CLK, Q => 
                           n_1150, QN => n511);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n9425, CK => CLK, Q => 
                           n_1151, QN => n512);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n9426, CK => CLK, Q => 
                           n_1152, QN => n513);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n9427, CK => CLK, Q => 
                           n_1153, QN => n514);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n9428, CK => CLK, Q => 
                           n_1154, QN => n515);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n9429, CK => CLK, Q => 
                           n_1155, QN => n516);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n9430, CK => CLK, Q => 
                           n_1156, QN => n517);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n9431, CK => CLK, Q => 
                           n_1157, QN => n518);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n9432, CK => CLK, Q => 
                           n_1158, QN => n519);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n9433, CK => CLK, Q => n7329
                           , QN => n520);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n9434, CK => CLK, Q => 
                           n_1159, QN => n521);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n9435, CK => CLK, Q => 
                           n_1160, QN => n522);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n9436, CK => CLK, Q => 
                           n_1161, QN => n523);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n9437, CK => CLK, Q => 
                           n_1162, QN => n524);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n9438, CK => CLK, Q => 
                           n_1163, QN => n525);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n9439, CK => CLK, Q => 
                           n_1164, QN => n526);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n9440, CK => CLK, Q => 
                           n_1165, QN => n527);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n9441, CK => CLK, Q => 
                           n_1166, QN => n528);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n9442, CK => CLK, Q => 
                           n_1167, QN => n529);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n9443, CK => CLK, Q => n_1168
                           , QN => n530);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n9444, CK => CLK, Q => n_1169
                           , QN => n531);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n9389, CK => CLK, Q => n7099
                           , QN => n966);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n9390, CK => CLK, Q => n7092
                           , QN => n970);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n9391, CK => CLK, Q => n7084
                           , QN => n972);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n9392, CK => CLK, Q => n7075
                           , QN => n976);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n9393, CK => CLK, Q => n7068
                           , QN => n978);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n9394, CK => CLK, Q => n7060
                           , QN => n982);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n9395, CK => CLK, Q => n7051
                           , QN => n984);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n9396, CK => CLK, Q => n7044
                           , QN => n988);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n9397, CK => CLK, Q => n7036
                           , QN => n990);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n9398, CK => CLK, Q => n7026
                           , QN => n994);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n9399, CK => CLK, Q => n7013
                           , QN => n996);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n9402, CK => CLK, Q => n6973
                           , QN => n1002);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n9403, CK => CLK, Q => n6963
                           , QN => n1003);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n9404, CK => CLK, Q => n6946
                           , QN => n1004);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n9405, CK => CLK, Q => n6937
                           , QN => n1005);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n9406, CK => CLK, Q => n6919
                           , QN => n1006);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n9407, CK => CLK, Q => n6907
                           , QN => n1007);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n9408, CK => CLK, Q => n6893
                           , QN => n1008);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n9409, CK => CLK, Q => n6880
                           , QN => n1009);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n9410, CK => CLK, Q => n6868
                           , QN => n1010);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n9411, CK => CLK, Q => n6853,
                           QN => n1011);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n9412, CK => CLK, Q => n6843,
                           QN => n1012);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n9357, CK => CLK, Q => n7972
                           , QN => n1013);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n9358, CK => CLK, Q => n7973
                           , QN => n1014);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n9359, CK => CLK, Q => n7974
                           , QN => n1015);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n9360, CK => CLK, Q => n7975
                           , QN => n1016);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n9361, CK => CLK, Q => n7976
                           , QN => n1017);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n9362, CK => CLK, Q => n7977
                           , QN => n1018);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n9363, CK => CLK, Q => n7978
                           , QN => n1019);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n9364, CK => CLK, Q => n7979
                           , QN => n1020);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n9365, CK => CLK, Q => n7980
                           , QN => n1021);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n9366, CK => CLK, Q => n7981
                           , QN => n1022);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n9367, CK => CLK, Q => n7982
                           , QN => n1023);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n9368, CK => CLK, Q => n7983
                           , QN => n1024);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n9370, CK => CLK, Q => n7985
                           , QN => n1026);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n9371, CK => CLK, Q => n7986
                           , QN => n1027);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n9372, CK => CLK, Q => n7987
                           , QN => n1028);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n9373, CK => CLK, Q => n7988
                           , QN => n1029);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n9374, CK => CLK, Q => n7989
                           , QN => n1030);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n9375, CK => CLK, Q => n7990
                           , QN => n1031);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n9376, CK => CLK, Q => n7991
                           , QN => n1032);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n9377, CK => CLK, Q => n7992
                           , QN => n1033);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n9378, CK => CLK, Q => n7993
                           , QN => n1034);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n9379, CK => CLK, Q => n7994,
                           QN => n1035);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n9380, CK => CLK, Q => n7995,
                           QN => n1036);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n9325, CK => CLK, Q => n7940
                           , QN => n532);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n9326, CK => CLK, Q => n7941
                           , QN => n533);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n9327, CK => CLK, Q => n7942
                           , QN => n534);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n9328, CK => CLK, Q => n7943
                           , QN => n535);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n9329, CK => CLK, Q => n7944
                           , QN => n536);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n9330, CK => CLK, Q => n7945
                           , QN => n537);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n9331, CK => CLK, Q => n7946
                           , QN => n538);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n9332, CK => CLK, Q => n7947
                           , QN => n539);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n9333, CK => CLK, Q => n7948
                           , QN => n540);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n9334, CK => CLK, Q => n7949
                           , QN => n541);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n9335, CK => CLK, Q => n7950
                           , QN => n542);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n9336, CK => CLK, Q => n7951
                           , QN => n543);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n9338, CK => CLK, Q => n7953
                           , QN => n545);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n9339, CK => CLK, Q => n7954
                           , QN => n546);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n9340, CK => CLK, Q => n7955
                           , QN => n547);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n9341, CK => CLK, Q => n7956
                           , QN => n548);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n9342, CK => CLK, Q => n7957
                           , QN => n549);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n9343, CK => CLK, Q => n7958
                           , QN => n550);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n9344, CK => CLK, Q => n7959
                           , QN => n551);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n9345, CK => CLK, Q => n7960
                           , QN => n552);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n9346, CK => CLK, Q => n7961
                           , QN => n553);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n9347, CK => CLK, Q => n7962,
                           QN => n554);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n9348, CK => CLK, Q => n7963,
                           QN => n555);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n9273, CK => CLK, Q => n803,
                           QN => n1892);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n9229, CK => CLK, Q => n7908
                           , QN => n580);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n9230, CK => CLK, Q => n7909
                           , QN => n581);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n9231, CK => CLK, Q => n7910
                           , QN => n582);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n9232, CK => CLK, Q => n7911
                           , QN => n583);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n9233, CK => CLK, Q => n7912
                           , QN => n584);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n9234, CK => CLK, Q => n7913
                           , QN => n585);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n9235, CK => CLK, Q => n7914
                           , QN => n586);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n9236, CK => CLK, Q => n7915
                           , QN => n587);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n9237, CK => CLK, Q => n7916
                           , QN => n588);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n9238, CK => CLK, Q => n7917
                           , QN => n589);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n9239, CK => CLK, Q => n7918
                           , QN => n590);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n9240, CK => CLK, Q => n7919
                           , QN => n591);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n9242, CK => CLK, Q => n7921
                           , QN => n593);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n9243, CK => CLK, Q => n7922
                           , QN => n594);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n9244, CK => CLK, Q => n7923
                           , QN => n595);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n9245, CK => CLK, Q => n7924
                           , QN => n596);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n9246, CK => CLK, Q => n7925
                           , QN => n597);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n9247, CK => CLK, Q => n7926
                           , QN => n598);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n9248, CK => CLK, Q => n7927
                           , QN => n599);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n9249, CK => CLK, Q => n7928
                           , QN => n600);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n9250, CK => CLK, Q => n7929
                           , QN => n601);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n9251, CK => CLK, Q => n7930,
                           QN => n602);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n9252, CK => CLK, Q => n7931,
                           QN => n603);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n9167, CK => CLK, Q => n7816
                           , QN => n604);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n9169, CK => CLK, Q => n7819
                           , QN => n605);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n9171, CK => CLK, Q => n7822
                           , QN => n606);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n9173, CK => CLK, Q => n7825
                           , QN => n607);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n9175, CK => CLK, Q => n7828
                           , QN => n608);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n9177, CK => CLK, Q => n7831
                           , QN => n609);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n9179, CK => CLK, Q => n7834
                           , QN => n610);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n9181, CK => CLK, Q => n7837
                           , QN => n611);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n9183, CK => CLK, Q => n7840
                           , QN => n612);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n9185, CK => CLK, Q => n7843
                           , QN => n613);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n9187, CK => CLK, Q => n7846
                           , QN => n614);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n9189, CK => CLK, Q => n7849
                           , QN => n615);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n9193, CK => CLK, Q => n7855
                           , QN => n617);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n9195, CK => CLK, Q => n7858
                           , QN => n618);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n9197, CK => CLK, Q => n7861
                           , QN => n619);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n9199, CK => CLK, Q => n7864
                           , QN => n620);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n9201, CK => CLK, Q => n7867
                           , QN => n621);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n9203, CK => CLK, Q => n7870
                           , QN => n622);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n9205, CK => CLK, Q => n7873
                           , QN => n623);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n9207, CK => CLK, Q => n7876
                           , QN => n624);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n9209, CK => CLK, Q => n7879
                           , QN => n625);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n9211, CK => CLK, Q => n7882,
                           QN => n626);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n9213, CK => CLK, Q => n7885,
                           QN => n627);
   REGISTERS_reg_70_21_inst : DFF_X1 port map( D => n11447, CK => CLK, Q => 
                           n735, QN => n1914);
   REGISTERS_reg_70_20_inst : DFF_X1 port map( D => n11448, CK => CLK, Q => 
                           n799, QN => n1915);
   REGISTERS_reg_70_17_inst : DFF_X1 port map( D => n11451, CK => CLK, Q => 
                           n995, QN => n628);
   REGISTERS_reg_70_16_inst : DFF_X1 port map( D => n11452, CK => CLK, Q => 
                           n989, QN => n629);
   REGISTERS_reg_70_15_inst : DFF_X1 port map( D => n11453, CK => CLK, Q => 
                           n983, QN => n630);
   REGISTERS_reg_70_14_inst : DFF_X1 port map( D => n11454, CK => CLK, Q => 
                           n977, QN => n631);
   REGISTERS_reg_70_13_inst : DFF_X1 port map( D => n11455, CK => CLK, Q => 
                           n971, QN => n632);
   REGISTERS_reg_70_12_inst : DFF_X1 port map( D => n11456, CK => CLK, Q => 
                           n965, QN => n633);
   REGISTERS_reg_70_11_inst : DFF_X1 port map( D => n11457, CK => CLK, Q => 
                           n959, QN => n634);
   REGISTERS_reg_70_10_inst : DFF_X1 port map( D => n11458, CK => CLK, Q => 
                           n953, QN => n635);
   REGISTERS_reg_70_9_inst : DFF_X1 port map( D => n11459, CK => CLK, Q => n947
                           , QN => n636);
   REGISTERS_reg_70_8_inst : DFF_X1 port map( D => n11460, CK => CLK, Q => n941
                           , QN => n637);
   REGISTERS_reg_69_21_inst : DFF_X1 port map( D => n11415, CK => CLK, Q => 
                           n734, QN => n1928);
   REGISTERS_reg_69_20_inst : DFF_X1 port map( D => n11416, CK => CLK, Q => 
                           n798, QN => n1929);
   REGISTERS_reg_68_31_inst : DFF_X1 port map( D => n11373, CK => CLK, Q => 
                           n8862, QN => n638);
   REGISTERS_reg_68_30_inst : DFF_X1 port map( D => n11374, CK => CLK, Q => 
                           n8863, QN => n639);
   REGISTERS_reg_68_29_inst : DFF_X1 port map( D => n11375, CK => CLK, Q => 
                           n8864, QN => n640);
   REGISTERS_reg_68_28_inst : DFF_X1 port map( D => n11376, CK => CLK, Q => 
                           n8865, QN => n641);
   REGISTERS_reg_68_27_inst : DFF_X1 port map( D => n11377, CK => CLK, Q => 
                           n8866, QN => n642);
   REGISTERS_reg_68_26_inst : DFF_X1 port map( D => n11378, CK => CLK, Q => 
                           n8867, QN => n643);
   REGISTERS_reg_68_25_inst : DFF_X1 port map( D => n11379, CK => CLK, Q => 
                           n8868, QN => n644);
   REGISTERS_reg_68_24_inst : DFF_X1 port map( D => n11380, CK => CLK, Q => 
                           n8869, QN => n645);
   REGISTERS_reg_68_23_inst : DFF_X1 port map( D => n11381, CK => CLK, Q => 
                           n8870, QN => n646);
   REGISTERS_reg_68_22_inst : DFF_X1 port map( D => n11382, CK => CLK, Q => 
                           n8871, QN => n647);
   REGISTERS_reg_68_21_inst : DFF_X1 port map( D => n11383, CK => CLK, Q => 
                           n8872, QN => n648);
   REGISTERS_reg_68_20_inst : DFF_X1 port map( D => n11384, CK => CLK, Q => 
                           n8873, QN => n649);
   REGISTERS_reg_68_19_inst : DFF_X1 port map( D => n11385, CK => CLK, Q => 
                           n8874, QN => n650);
   REGISTERS_reg_68_18_inst : DFF_X1 port map( D => n11386, CK => CLK, Q => 
                           n8875, QN => n651);
   REGISTERS_reg_68_17_inst : DFF_X1 port map( D => n11387, CK => CLK, Q => 
                           n8876, QN => n652);
   REGISTERS_reg_68_16_inst : DFF_X1 port map( D => n11388, CK => CLK, Q => 
                           n8877, QN => n653);
   REGISTERS_reg_68_15_inst : DFF_X1 port map( D => n11389, CK => CLK, Q => 
                           n8878, QN => n654);
   REGISTERS_reg_68_14_inst : DFF_X1 port map( D => n11390, CK => CLK, Q => 
                           n8879, QN => n655);
   REGISTERS_reg_68_13_inst : DFF_X1 port map( D => n11391, CK => CLK, Q => 
                           n8880, QN => n656);
   REGISTERS_reg_68_12_inst : DFF_X1 port map( D => n11392, CK => CLK, Q => 
                           n8881, QN => n657);
   REGISTERS_reg_68_11_inst : DFF_X1 port map( D => n11393, CK => CLK, Q => 
                           n8882, QN => n658);
   REGISTERS_reg_68_10_inst : DFF_X1 port map( D => n11394, CK => CLK, Q => 
                           n8883, QN => n659);
   REGISTERS_reg_68_9_inst : DFF_X1 port map( D => n11395, CK => CLK, Q => 
                           n8884, QN => n660);
   REGISTERS_reg_68_8_inst : DFF_X1 port map( D => n11396, CK => CLK, Q => 
                           n8885, QN => n661);
   REGISTERS_reg_67_31_inst : DFF_X1 port map( D => n11341, CK => CLK, Q => 
                           n8830, QN => n662);
   REGISTERS_reg_67_30_inst : DFF_X1 port map( D => n11342, CK => CLK, Q => 
                           n8831, QN => n663);
   REGISTERS_reg_67_29_inst : DFF_X1 port map( D => n11343, CK => CLK, Q => 
                           n8832, QN => n664);
   REGISTERS_reg_67_28_inst : DFF_X1 port map( D => n11344, CK => CLK, Q => 
                           n8833, QN => n665);
   REGISTERS_reg_67_27_inst : DFF_X1 port map( D => n11345, CK => CLK, Q => 
                           n8834, QN => n666);
   REGISTERS_reg_67_26_inst : DFF_X1 port map( D => n11346, CK => CLK, Q => 
                           n8835, QN => n667);
   REGISTERS_reg_67_25_inst : DFF_X1 port map( D => n11347, CK => CLK, Q => 
                           n8836, QN => n668);
   REGISTERS_reg_67_24_inst : DFF_X1 port map( D => n11348, CK => CLK, Q => 
                           n8837, QN => n669);
   REGISTERS_reg_67_23_inst : DFF_X1 port map( D => n11349, CK => CLK, Q => 
                           n8838, QN => n670);
   REGISTERS_reg_67_22_inst : DFF_X1 port map( D => n11350, CK => CLK, Q => 
                           n8839, QN => n671);
   REGISTERS_reg_67_21_inst : DFF_X1 port map( D => n11351, CK => CLK, Q => 
                           n8840, QN => n672);
   REGISTERS_reg_67_20_inst : DFF_X1 port map( D => n11352, CK => CLK, Q => 
                           n8841, QN => n673);
   REGISTERS_reg_67_19_inst : DFF_X1 port map( D => n11353, CK => CLK, Q => 
                           n8842, QN => n674);
   REGISTERS_reg_67_18_inst : DFF_X1 port map( D => n11354, CK => CLK, Q => 
                           n8843, QN => n675);
   REGISTERS_reg_67_17_inst : DFF_X1 port map( D => n11355, CK => CLK, Q => 
                           n8844, QN => n676);
   REGISTERS_reg_67_16_inst : DFF_X1 port map( D => n11356, CK => CLK, Q => 
                           n8845, QN => n677);
   REGISTERS_reg_67_15_inst : DFF_X1 port map( D => n11357, CK => CLK, Q => 
                           n8846, QN => n678);
   REGISTERS_reg_67_14_inst : DFF_X1 port map( D => n11358, CK => CLK, Q => 
                           n8847, QN => n679);
   REGISTERS_reg_67_13_inst : DFF_X1 port map( D => n11359, CK => CLK, Q => 
                           n8848, QN => n680);
   REGISTERS_reg_67_12_inst : DFF_X1 port map( D => n11360, CK => CLK, Q => 
                           n8849, QN => n681);
   REGISTERS_reg_67_11_inst : DFF_X1 port map( D => n11361, CK => CLK, Q => 
                           n8850, QN => n682);
   REGISTERS_reg_67_10_inst : DFF_X1 port map( D => n11362, CK => CLK, Q => 
                           n8851, QN => n683);
   REGISTERS_reg_67_9_inst : DFF_X1 port map( D => n11363, CK => CLK, Q => 
                           n8852, QN => n684);
   REGISTERS_reg_67_8_inst : DFF_X1 port map( D => n11364, CK => CLK, Q => 
                           n8853, QN => n685);
   REGISTERS_reg_66_31_inst : DFF_X1 port map( D => n11309, CK => CLK, Q => 
                           n7205, QN => n686);
   REGISTERS_reg_66_30_inst : DFF_X1 port map( D => n11310, CK => CLK, Q => 
                           n7204, QN => n687);
   REGISTERS_reg_66_29_inst : DFF_X1 port map( D => n11311, CK => CLK, Q => 
                           n7203, QN => n688);
   REGISTERS_reg_66_28_inst : DFF_X1 port map( D => n11312, CK => CLK, Q => 
                           n7181, QN => n689);
   REGISTERS_reg_66_27_inst : DFF_X1 port map( D => n11313, CK => CLK, Q => 
                           n7180, QN => n690);
   REGISTERS_reg_66_26_inst : DFF_X1 port map( D => n11314, CK => CLK, Q => 
                           n7179, QN => n691);
   REGISTERS_reg_66_25_inst : DFF_X1 port map( D => n11315, CK => CLK, Q => 
                           n7157, QN => n692);
   REGISTERS_reg_66_24_inst : DFF_X1 port map( D => n11316, CK => CLK, Q => 
                           n7156, QN => n693);
   REGISTERS_reg_66_23_inst : DFF_X1 port map( D => n11317, CK => CLK, Q => 
                           n7155, QN => n694);
   REGISTERS_reg_66_22_inst : DFF_X1 port map( D => n11318, CK => CLK, Q => 
                           n7153, QN => n695);
   REGISTERS_reg_66_19_inst : DFF_X1 port map( D => n11321, CK => CLK, Q => 
                           n7143, QN => n698);
   REGISTERS_reg_66_18_inst : DFF_X1 port map( D => n11322, CK => CLK, Q => 
                           n7141, QN => n699);
   REGISTERS_reg_66_17_inst : DFF_X1 port map( D => n11323, CK => CLK, Q => 
                           n7140, QN => n700);
   REGISTERS_reg_66_16_inst : DFF_X1 port map( D => n11324, CK => CLK, Q => 
                           n7138, QN => n701);
   REGISTERS_reg_66_15_inst : DFF_X1 port map( D => n11325, CK => CLK, Q => 
                           n7137, QN => n702);
   REGISTERS_reg_66_14_inst : DFF_X1 port map( D => n11326, CK => CLK, Q => 
                           n7135, QN => n703);
   REGISTERS_reg_66_13_inst : DFF_X1 port map( D => n11327, CK => CLK, Q => 
                           n7133, QN => n704);
   REGISTERS_reg_66_12_inst : DFF_X1 port map( D => n11328, CK => CLK, Q => 
                           n7132, QN => n705);
   REGISTERS_reg_66_11_inst : DFF_X1 port map( D => n11329, CK => CLK, Q => 
                           n7131, QN => n706);
   REGISTERS_reg_66_10_inst : DFF_X1 port map( D => n11330, CK => CLK, Q => 
                           n7129, QN => n707);
   REGISTERS_reg_66_9_inst : DFF_X1 port map( D => n11331, CK => CLK, Q => 
                           n7128, QN => n708);
   REGISTERS_reg_66_8_inst : DFF_X1 port map( D => n11332, CK => CLK, Q => 
                           n7125, QN => n709);
   REGISTERS_reg_65_31_inst : DFF_X1 port map( D => n11277, CK => CLK, Q => 
                           n_1170, QN => n710);
   REGISTERS_reg_65_30_inst : DFF_X1 port map( D => n11278, CK => CLK, Q => 
                           n_1171, QN => n711);
   REGISTERS_reg_65_29_inst : DFF_X1 port map( D => n11279, CK => CLK, Q => 
                           n_1172, QN => n712);
   REGISTERS_reg_65_28_inst : DFF_X1 port map( D => n11280, CK => CLK, Q => 
                           n_1173, QN => n713);
   REGISTERS_reg_65_27_inst : DFF_X1 port map( D => n11281, CK => CLK, Q => 
                           n_1174, QN => n714);
   REGISTERS_reg_65_26_inst : DFF_X1 port map( D => n11282, CK => CLK, Q => 
                           n_1175, QN => n715);
   REGISTERS_reg_65_25_inst : DFF_X1 port map( D => n11283, CK => CLK, Q => 
                           n_1176, QN => n716);
   REGISTERS_reg_65_24_inst : DFF_X1 port map( D => n11284, CK => CLK, Q => 
                           n_1177, QN => n717);
   REGISTERS_reg_65_23_inst : DFF_X1 port map( D => n11285, CK => CLK, Q => 
                           n_1178, QN => n718);
   REGISTERS_reg_65_22_inst : DFF_X1 port map( D => n11286, CK => CLK, Q => 
                           n_1179, QN => n719);
   REGISTERS_reg_65_21_inst : DFF_X1 port map( D => n11287, CK => CLK, Q => 
                           n_1180, QN => n720);
   REGISTERS_reg_65_20_inst : DFF_X1 port map( D => n11288, CK => CLK, Q => 
                           n_1181, QN => n721);
   REGISTERS_reg_65_19_inst : DFF_X1 port map( D => n11289, CK => CLK, Q => 
                           n_1182, QN => n722);
   REGISTERS_reg_65_18_inst : DFF_X1 port map( D => n11290, CK => CLK, Q => 
                           n_1183, QN => n723);
   REGISTERS_reg_65_17_inst : DFF_X1 port map( D => n11291, CK => CLK, Q => 
                           n_1184, QN => n724);
   REGISTERS_reg_65_16_inst : DFF_X1 port map( D => n11292, CK => CLK, Q => 
                           n_1185, QN => n725);
   REGISTERS_reg_65_15_inst : DFF_X1 port map( D => n11293, CK => CLK, Q => 
                           n_1186, QN => n726);
   REGISTERS_reg_65_14_inst : DFF_X1 port map( D => n11294, CK => CLK, Q => 
                           n_1187, QN => n728);
   REGISTERS_reg_65_13_inst : DFF_X1 port map( D => n11295, CK => CLK, Q => 
                           n_1188, QN => n729);
   REGISTERS_reg_65_12_inst : DFF_X1 port map( D => n11296, CK => CLK, Q => 
                           n_1189, QN => n730);
   REGISTERS_reg_65_11_inst : DFF_X1 port map( D => n11297, CK => CLK, Q => 
                           n_1190, QN => n732);
   REGISTERS_reg_65_10_inst : DFF_X1 port map( D => n11298, CK => CLK, Q => 
                           n_1191, QN => n733);
   REGISTERS_reg_65_9_inst : DFF_X1 port map( D => n11299, CK => CLK, Q => 
                           n_1192, QN => n737);
   REGISTERS_reg_65_8_inst : DFF_X1 port map( D => n11300, CK => CLK, Q => 
                           n_1193, QN => n738);
   REGISTERS_reg_64_31_inst : DFF_X1 port map( D => n11245, CK => CLK, Q => 
                           n8799, QN => n739);
   REGISTERS_reg_64_30_inst : DFF_X1 port map( D => n11246, CK => CLK, Q => 
                           n8800, QN => n740);
   REGISTERS_reg_64_29_inst : DFF_X1 port map( D => n11247, CK => CLK, Q => 
                           n8801, QN => n741);
   REGISTERS_reg_64_28_inst : DFF_X1 port map( D => n11248, CK => CLK, Q => 
                           n8802, QN => n742);
   REGISTERS_reg_64_27_inst : DFF_X1 port map( D => n11249, CK => CLK, Q => 
                           n8803, QN => n744);
   REGISTERS_reg_64_26_inst : DFF_X1 port map( D => n11250, CK => CLK, Q => 
                           n8804, QN => n745);
   REGISTERS_reg_64_25_inst : DFF_X1 port map( D => n11251, CK => CLK, Q => 
                           n8805, QN => n746);
   REGISTERS_reg_64_24_inst : DFF_X1 port map( D => n11252, CK => CLK, Q => 
                           n8806, QN => n747);
   REGISTERS_reg_64_23_inst : DFF_X1 port map( D => n11253, CK => CLK, Q => 
                           n8807, QN => n748);
   REGISTERS_reg_64_22_inst : DFF_X1 port map( D => n11254, CK => CLK, Q => 
                           n8808, QN => n749);
   REGISTERS_reg_64_21_inst : DFF_X1 port map( D => n11255, CK => CLK, Q => 
                           n8809, QN => n750);
   REGISTERS_reg_64_20_inst : DFF_X1 port map( D => n11256, CK => CLK, Q => 
                           n8810, QN => n751);
   REGISTERS_reg_64_19_inst : DFF_X1 port map( D => n11257, CK => CLK, Q => 
                           n8811, QN => n755);
   REGISTERS_reg_64_18_inst : DFF_X1 port map( D => n11258, CK => CLK, Q => 
                           n8812, QN => n757);
   REGISTERS_reg_64_17_inst : DFF_X1 port map( D => n11259, CK => CLK, Q => 
                           n8813, QN => n758);
   REGISTERS_reg_64_16_inst : DFF_X1 port map( D => n11260, CK => CLK, Q => 
                           n8814, QN => n759);
   REGISTERS_reg_64_15_inst : DFF_X1 port map( D => n11261, CK => CLK, Q => 
                           n8815, QN => n760);
   REGISTERS_reg_64_14_inst : DFF_X1 port map( D => n11262, CK => CLK, Q => 
                           n8816, QN => n764);
   REGISTERS_reg_64_13_inst : DFF_X1 port map( D => n11263, CK => CLK, Q => 
                           n8817, QN => n765);
   REGISTERS_reg_64_12_inst : DFF_X1 port map( D => n11264, CK => CLK, Q => 
                           n8818, QN => n766);
   REGISTERS_reg_64_11_inst : DFF_X1 port map( D => n11265, CK => CLK, Q => 
                           n8819, QN => n767);
   REGISTERS_reg_64_10_inst : DFF_X1 port map( D => n11266, CK => CLK, Q => 
                           n8820, QN => n768);
   REGISTERS_reg_64_9_inst : DFF_X1 port map( D => n11267, CK => CLK, Q => 
                           n8821, QN => n769);
   REGISTERS_reg_64_8_inst : DFF_X1 port map( D => n11268, CK => CLK, Q => 
                           n8822, QN => n771);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n9485, CK => CLK, Q => n8004
                           , QN => n772);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n9486, CK => CLK, Q => n8005
                           , QN => n773);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n9487, CK => CLK, Q => n8006
                           , QN => n775);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n9488, CK => CLK, Q => n8007
                           , QN => n776);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n9489, CK => CLK, Q => n8008
                           , QN => n778);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n9490, CK => CLK, Q => n8009
                           , QN => n779);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n9491, CK => CLK, Q => n8010
                           , QN => n780);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n9492, CK => CLK, Q => n8011
                           , QN => n781);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n9493, CK => CLK, Q => n8012
                           , QN => n782);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n9494, CK => CLK, Q => n8013
                           , QN => n783);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n9495, CK => CLK, Q => n8014
                           , QN => n785);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n9496, CK => CLK, Q => n8015
                           , QN => n787);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n9498, CK => CLK, Q => n8017
                           , QN => n789);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n9499, CK => CLK, Q => n8018
                           , QN => n790);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n9500, CK => CLK, Q => n8019
                           , QN => n792);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n9501, CK => CLK, Q => n8020
                           , QN => n793);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n9502, CK => CLK, Q => n8021
                           , QN => n794);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n9503, CK => CLK, Q => n8022
                           , QN => n796);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n9504, CK => CLK, Q => n8023
                           , QN => n797);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n9505, CK => CLK, Q => n8024
                           , QN => n804);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n9506, CK => CLK, Q => n8025
                           , QN => n808);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n9507, CK => CLK, Q => n8026,
                           QN => n809);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n9508, CK => CLK, Q => n8027,
                           QN => n813);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n9453, CK => CLK, Q => 
                           n_1194, QN => n819);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n9454, CK => CLK, Q => 
                           n_1195, QN => n898);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n9455, CK => CLK, Q => 
                           n_1196, QN => n900);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n9456, CK => CLK, Q => 
                           n_1197, QN => n904);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n9457, CK => CLK, Q => 
                           n_1198, QN => n906);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n9458, CK => CLK, Q => 
                           n_1199, QN => n910);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n9459, CK => CLK, Q => 
                           n_1200, QN => n912);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n9460, CK => CLK, Q => 
                           n_1201, QN => n916);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n9461, CK => CLK, Q => 
                           n_1202, QN => n918);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n9462, CK => CLK, Q => 
                           n_1203, QN => n922);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n9463, CK => CLK, Q => 
                           n_1204, QN => n924);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n9464, CK => CLK, Q => 
                           n_1205, QN => n928);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n9465, CK => CLK, Q => n7325
                           , QN => n930);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n9466, CK => CLK, Q => 
                           n_1206, QN => n934);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n9467, CK => CLK, Q => 
                           n_1207, QN => n936);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n9468, CK => CLK, Q => 
                           n_1208, QN => n940);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n9469, CK => CLK, Q => 
                           n_1209, QN => n942);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n9470, CK => CLK, Q => 
                           n_1210, QN => n946);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n9471, CK => CLK, Q => 
                           n_1211, QN => n948);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n9472, CK => CLK, Q => 
                           n_1212, QN => n952);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n9473, CK => CLK, Q => 
                           n_1213, QN => n954);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n9474, CK => CLK, Q => 
                           n_1214, QN => n958);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n9475, CK => CLK, Q => n_1215
                           , QN => n960);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n9476, CK => CLK, Q => n_1216
                           , QN => n964);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n9293, CK => CLK, Q => n895,
                           QN => n556);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n9294, CK => CLK, Q => n893,
                           QN => n557);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n9295, CK => CLK, Q => n891,
                           QN => n558);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n9296, CK => CLK, Q => n889,
                           QN => n559);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n9297, CK => CLK, Q => n887,
                           QN => n560);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n9298, CK => CLK, Q => n885,
                           QN => n561);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n9299, CK => CLK, Q => n883,
                           QN => n562);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n9300, CK => CLK, Q => n881,
                           QN => n563);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n9301, CK => CLK, Q => n879,
                           QN => n564);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n9302, CK => CLK, Q => n877,
                           QN => n565);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n9303, CK => CLK, Q => n875,
                           QN => n566);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n9304, CK => CLK, Q => n873,
                           QN => n567);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n9305, CK => CLK, Q => n871,
                           QN => n568);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n9306, CK => CLK, Q => n869,
                           QN => n569);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n9307, CK => CLK, Q => n867,
                           QN => n570);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n9308, CK => CLK, Q => n865,
                           QN => n571);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n9309, CK => CLK, Q => n863,
                           QN => n572);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n9310, CK => CLK, Q => n861,
                           QN => n573);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n9311, CK => CLK, Q => n859,
                           QN => n574);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n9312, CK => CLK, Q => n857,
                           QN => n575);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n9313, CK => CLK, Q => n855,
                           QN => n576);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n9314, CK => CLK, Q => n853,
                           QN => n577);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n9315, CK => CLK, Q => n851, 
                           QN => n578);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n9316, CK => CLK, Q => n849, 
                           QN => n579);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n10189, CK => CLK, Q => 
                           n8258, QN => n1037);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n10190, CK => CLK, Q => 
                           n8259, QN => n1038);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n10191, CK => CLK, Q => 
                           n8260, QN => n1039);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n10192, CK => CLK, Q => 
                           n8261, QN => n1040);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n10193, CK => CLK, Q => 
                           n8262, QN => n1041);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n10194, CK => CLK, Q => 
                           n8263, QN => n1042);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n10195, CK => CLK, Q => 
                           n8264, QN => n1043);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n10196, CK => CLK, Q => 
                           n8265, QN => n1044);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n10197, CK => CLK, Q => 
                           n8266, QN => n1045);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n10198, CK => CLK, Q => 
                           n8267, QN => n1046);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n10199, CK => CLK, Q => 
                           n8268, QN => n1047);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n10200, CK => CLK, Q => 
                           n8269, QN => n1048);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n10201, CK => CLK, Q => 
                           n8270, QN => n1049);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n10202, CK => CLK, Q => 
                           n8271, QN => n1050);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n10203, CK => CLK, Q => 
                           n8272, QN => n1051);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n10204, CK => CLK, Q => 
                           n8273, QN => n1052);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n10205, CK => CLK, Q => 
                           n8274, QN => n1053);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n10206, CK => CLK, Q => 
                           n8275, QN => n1054);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n10207, CK => CLK, Q => 
                           n8276, QN => n1055);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n10208, CK => CLK, Q => 
                           n8277, QN => n1056);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n10209, CK => CLK, Q => 
                           n8278, QN => n1057);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n10210, CK => CLK, Q => 
                           n8279, QN => n1058);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n10211, CK => CLK, Q => 
                           n8280, QN => n1059);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n10212, CK => CLK, Q => 
                           n8281, QN => n1060);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n10157, CK => CLK, Q => 
                           n897, QN => n1061);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n10093, CK => CLK, Q => 
                           n_1217, QN => n1062);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n10094, CK => CLK, Q => 
                           n_1218, QN => n1063);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n10095, CK => CLK, Q => 
                           n_1219, QN => n1064);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n10096, CK => CLK, Q => 
                           n_1220, QN => n1065);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n10097, CK => CLK, Q => 
                           n_1221, QN => n1066);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n10098, CK => CLK, Q => 
                           n_1222, QN => n1067);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n10099, CK => CLK, Q => 
                           n_1223, QN => n1068);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n10100, CK => CLK, Q => 
                           n_1224, QN => n1069);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n10101, CK => CLK, Q => 
                           n_1225, QN => n1070);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n10102, CK => CLK, Q => 
                           n_1226, QN => n1071);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n10103, CK => CLK, Q => 
                           n_1227, QN => n1072);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n10104, CK => CLK, Q => 
                           n_1228, QN => n1073);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n10106, CK => CLK, Q => 
                           n_1229, QN => n1074);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n10107, CK => CLK, Q => 
                           n_1230, QN => n1075);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n10108, CK => CLK, Q => 
                           n_1231, QN => n1076);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n10109, CK => CLK, Q => 
                           n_1232, QN => n1077);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n10110, CK => CLK, Q => 
                           n_1233, QN => n1078);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n10111, CK => CLK, Q => 
                           n_1234, QN => n1079);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n10112, CK => CLK, Q => 
                           n_1235, QN => n1080);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n10113, CK => CLK, Q => 
                           n_1236, QN => n1081);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n10114, CK => CLK, Q => 
                           n_1237, QN => n1082);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n10115, CK => CLK, Q => 
                           n_1238, QN => n1083);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n10116, CK => CLK, Q => 
                           n_1239, QN => n1084);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n10061, CK => CLK, Q => 
                           n_1240, QN => n1607);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n10064, CK => CLK, Q => 
                           n_1241, QN => n1707);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n10065, CK => CLK, Q => 
                           n_1242, QN => n1087);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n10066, CK => CLK, Q => 
                           n_1243, QN => n1088);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n10067, CK => CLK, Q => 
                           n_1244, QN => n1089);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n10068, CK => CLK, Q => 
                           n_1245, QN => n1090);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n10069, CK => CLK, Q => 
                           n_1246, QN => n1091);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n10070, CK => CLK, Q => 
                           n_1247, QN => n1092);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n10071, CK => CLK, Q => 
                           n_1248, QN => n1093);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n10072, CK => CLK, Q => 
                           n_1249, QN => n1094);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n10074, CK => CLK, Q => 
                           n_1250, QN => n1095);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n10075, CK => CLK, Q => 
                           n_1251, QN => n1096);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n10076, CK => CLK, Q => 
                           n_1252, QN => n1097);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n10077, CK => CLK, Q => 
                           n_1253, QN => n1098);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n10078, CK => CLK, Q => 
                           n_1254, QN => n1099);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n10079, CK => CLK, Q => 
                           n_1255, QN => n1100);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n10080, CK => CLK, Q => 
                           n_1256, QN => n1101);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n10081, CK => CLK, Q => 
                           n_1257, QN => n1102);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n10082, CK => CLK, Q => 
                           n_1258, QN => n1103);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n10083, CK => CLK, Q => 
                           n_1259, QN => n1104);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n10084, CK => CLK, Q => 
                           n_1260, QN => n1105);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n9976, CK => CLK, Q => n761
                           , QN => n1997);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n9977, CK => CLK, Q => n825
                           , QN => n1998);
   REGISTERS_reg_63_31_inst : DFF_X1 port map( D => n11213, CK => CLK, Q => 
                           n8768, QN => n1106);
   REGISTERS_reg_63_30_inst : DFF_X1 port map( D => n11214, CK => CLK, Q => 
                           n8769, QN => n1107);
   REGISTERS_reg_63_29_inst : DFF_X1 port map( D => n11215, CK => CLK, Q => 
                           n8770, QN => n1108);
   REGISTERS_reg_63_28_inst : DFF_X1 port map( D => n11216, CK => CLK, Q => 
                           n8771, QN => n1109);
   REGISTERS_reg_63_27_inst : DFF_X1 port map( D => n11217, CK => CLK, Q => 
                           n8772, QN => n1110);
   REGISTERS_reg_63_26_inst : DFF_X1 port map( D => n11218, CK => CLK, Q => 
                           n8773, QN => n1111);
   REGISTERS_reg_63_25_inst : DFF_X1 port map( D => n11219, CK => CLK, Q => 
                           n8774, QN => n1112);
   REGISTERS_reg_63_24_inst : DFF_X1 port map( D => n11220, CK => CLK, Q => 
                           n8775, QN => n1113);
   REGISTERS_reg_63_23_inst : DFF_X1 port map( D => n11221, CK => CLK, Q => 
                           n8776, QN => n1114);
   REGISTERS_reg_63_22_inst : DFF_X1 port map( D => n11222, CK => CLK, Q => 
                           n8777, QN => n1115);
   REGISTERS_reg_63_21_inst : DFF_X1 port map( D => n11223, CK => CLK, Q => 
                           n8778, QN => n1116);
   REGISTERS_reg_63_20_inst : DFF_X1 port map( D => n11224, CK => CLK, Q => 
                           n8779, QN => n1117);
   REGISTERS_reg_63_19_inst : DFF_X1 port map( D => n11225, CK => CLK, Q => 
                           n8780, QN => n1118);
   REGISTERS_reg_63_18_inst : DFF_X1 port map( D => n11226, CK => CLK, Q => 
                           n8781, QN => n1119);
   REGISTERS_reg_63_17_inst : DFF_X1 port map( D => n11227, CK => CLK, Q => 
                           n8782, QN => n1120);
   REGISTERS_reg_63_16_inst : DFF_X1 port map( D => n11228, CK => CLK, Q => 
                           n8783, QN => n1121);
   REGISTERS_reg_63_15_inst : DFF_X1 port map( D => n11229, CK => CLK, Q => 
                           n8784, QN => n1122);
   REGISTERS_reg_63_14_inst : DFF_X1 port map( D => n11230, CK => CLK, Q => 
                           n8785, QN => n1123);
   REGISTERS_reg_63_13_inst : DFF_X1 port map( D => n11231, CK => CLK, Q => 
                           n8786, QN => n1124);
   REGISTERS_reg_63_12_inst : DFF_X1 port map( D => n11232, CK => CLK, Q => 
                           n8787, QN => n1125);
   REGISTERS_reg_63_11_inst : DFF_X1 port map( D => n11233, CK => CLK, Q => 
                           n8788, QN => n1126);
   REGISTERS_reg_63_10_inst : DFF_X1 port map( D => n11234, CK => CLK, Q => 
                           n8789, QN => n1127);
   REGISTERS_reg_63_9_inst : DFF_X1 port map( D => n11235, CK => CLK, Q => 
                           n8790, QN => n1128);
   REGISTERS_reg_63_8_inst : DFF_X1 port map( D => n11236, CK => CLK, Q => 
                           n8791, QN => n1129);
   REGISTERS_reg_62_31_inst : DFF_X1 port map( D => n11181, CK => CLK, Q => 
                           n_1261, QN => n2010);
   REGISTERS_reg_62_30_inst : DFF_X1 port map( D => n11182, CK => CLK, Q => 
                           n_1262, QN => n2011);
   REGISTERS_reg_62_29_inst : DFF_X1 port map( D => n11183, CK => CLK, Q => 
                           n_1263, QN => n2012);
   REGISTERS_reg_62_28_inst : DFF_X1 port map( D => n11184, CK => CLK, Q => 
                           n_1264, QN => n2013);
   REGISTERS_reg_62_27_inst : DFF_X1 port map( D => n11185, CK => CLK, Q => 
                           n_1265, QN => n2014);
   REGISTERS_reg_62_26_inst : DFF_X1 port map( D => n11186, CK => CLK, Q => 
                           n_1266, QN => n2015);
   REGISTERS_reg_62_25_inst : DFF_X1 port map( D => n11187, CK => CLK, Q => 
                           n_1267, QN => n2016);
   REGISTERS_reg_62_24_inst : DFF_X1 port map( D => n11188, CK => CLK, Q => 
                           n_1268, QN => n2017);
   REGISTERS_reg_62_23_inst : DFF_X1 port map( D => n11189, CK => CLK, Q => 
                           n_1269, QN => n2018);
   REGISTERS_reg_62_22_inst : DFF_X1 port map( D => n11190, CK => CLK, Q => 
                           n_1270, QN => n2019);
   REGISTERS_reg_62_21_inst : DFF_X1 port map( D => n11191, CK => CLK, Q => 
                           n_1271, QN => n2020);
   REGISTERS_reg_62_20_inst : DFF_X1 port map( D => n11192, CK => CLK, Q => 
                           n_1272, QN => n2021);
   REGISTERS_reg_62_19_inst : DFF_X1 port map( D => n11193, CK => CLK, Q => 
                           n_1273, QN => n2022);
   REGISTERS_reg_62_18_inst : DFF_X1 port map( D => n11194, CK => CLK, Q => 
                           n_1274, QN => n2023);
   REGISTERS_reg_62_17_inst : DFF_X1 port map( D => n11195, CK => CLK, Q => 
                           n_1275, QN => n1130);
   REGISTERS_reg_62_16_inst : DFF_X1 port map( D => n11196, CK => CLK, Q => 
                           n_1276, QN => n1131);
   REGISTERS_reg_62_15_inst : DFF_X1 port map( D => n11197, CK => CLK, Q => 
                           n_1277, QN => n1132);
   REGISTERS_reg_62_14_inst : DFF_X1 port map( D => n11198, CK => CLK, Q => 
                           n_1278, QN => n1133);
   REGISTERS_reg_62_13_inst : DFF_X1 port map( D => n11199, CK => CLK, Q => 
                           n_1279, QN => n1134);
   REGISTERS_reg_62_12_inst : DFF_X1 port map( D => n11200, CK => CLK, Q => 
                           n_1280, QN => n2024);
   REGISTERS_reg_62_11_inst : DFF_X1 port map( D => n11201, CK => CLK, Q => 
                           n_1281, QN => n2025);
   REGISTERS_reg_62_10_inst : DFF_X1 port map( D => n11202, CK => CLK, Q => 
                           n_1282, QN => n2026);
   REGISTERS_reg_62_9_inst : DFF_X1 port map( D => n11203, CK => CLK, Q => 
                           n_1283, QN => n2027);
   REGISTERS_reg_62_8_inst : DFF_X1 port map( D => n11204, CK => CLK, Q => 
                           n_1284, QN => n2028);
   REGISTERS_reg_61_31_inst : DFF_X1 port map( D => n11149, CK => CLK, Q => 
                           n_1285, QN => n2029);
   REGISTERS_reg_61_30_inst : DFF_X1 port map( D => n11150, CK => CLK, Q => 
                           n_1286, QN => n2030);
   REGISTERS_reg_61_29_inst : DFF_X1 port map( D => n11151, CK => CLK, Q => 
                           n_1287, QN => n2031);
   REGISTERS_reg_61_28_inst : DFF_X1 port map( D => n11152, CK => CLK, Q => 
                           n_1288, QN => n2032);
   REGISTERS_reg_61_27_inst : DFF_X1 port map( D => n11153, CK => CLK, Q => 
                           n_1289, QN => n2033);
   REGISTERS_reg_61_26_inst : DFF_X1 port map( D => n11154, CK => CLK, Q => 
                           n_1290, QN => n2034);
   REGISTERS_reg_61_25_inst : DFF_X1 port map( D => n11155, CK => CLK, Q => 
                           n_1291, QN => n2035);
   REGISTERS_reg_61_24_inst : DFF_X1 port map( D => n11156, CK => CLK, Q => 
                           n_1292, QN => n2036);
   REGISTERS_reg_61_23_inst : DFF_X1 port map( D => n11157, CK => CLK, Q => 
                           n_1293, QN => n2037);
   REGISTERS_reg_61_22_inst : DFF_X1 port map( D => n11158, CK => CLK, Q => 
                           n_1294, QN => n2038);
   REGISTERS_reg_61_21_inst : DFF_X1 port map( D => n11159, CK => CLK, Q => 
                           n_1295, QN => n2039);
   REGISTERS_reg_61_20_inst : DFF_X1 port map( D => n11160, CK => CLK, Q => 
                           n_1296, QN => n2040);
   REGISTERS_reg_61_19_inst : DFF_X1 port map( D => n11161, CK => CLK, Q => 
                           n_1297, QN => n2041);
   REGISTERS_reg_61_18_inst : DFF_X1 port map( D => n11162, CK => CLK, Q => 
                           n_1298, QN => n2042);
   REGISTERS_reg_61_17_inst : DFF_X1 port map( D => n11163, CK => CLK, Q => 
                           n_1299, QN => n1135);
   REGISTERS_reg_61_16_inst : DFF_X1 port map( D => n11164, CK => CLK, Q => 
                           n_1300, QN => n1136);
   REGISTERS_reg_61_15_inst : DFF_X1 port map( D => n11165, CK => CLK, Q => 
                           n_1301, QN => n1137);
   REGISTERS_reg_61_14_inst : DFF_X1 port map( D => n11166, CK => CLK, Q => 
                           n_1302, QN => n1138);
   REGISTERS_reg_61_13_inst : DFF_X1 port map( D => n11167, CK => CLK, Q => 
                           n_1303, QN => n1139);
   REGISTERS_reg_61_12_inst : DFF_X1 port map( D => n11168, CK => CLK, Q => 
                           n_1304, QN => n1140);
   REGISTERS_reg_61_11_inst : DFF_X1 port map( D => n11169, CK => CLK, Q => 
                           n_1305, QN => n1141);
   REGISTERS_reg_61_10_inst : DFF_X1 port map( D => n11170, CK => CLK, Q => 
                           n_1306, QN => n1142);
   REGISTERS_reg_61_9_inst : DFF_X1 port map( D => n11171, CK => CLK, Q => 
                           n_1307, QN => n1143);
   REGISTERS_reg_61_8_inst : DFF_X1 port map( D => n11172, CK => CLK, Q => 
                           n_1308, QN => n1144);
   REGISTERS_reg_60_21_inst : DFF_X1 port map( D => n11127, CK => CLK, Q => 
                           n727, QN => n2053);
   REGISTERS_reg_60_20_inst : DFF_X1 port map( D => n11128, CK => CLK, Q => 
                           n791, QN => n2054);
   REGISTERS_reg_59_31_inst : DFF_X1 port map( D => n11085, CK => CLK, Q => 
                           n8736, QN => n1145);
   REGISTERS_reg_59_30_inst : DFF_X1 port map( D => n11086, CK => CLK, Q => 
                           n8737, QN => n1146);
   REGISTERS_reg_59_29_inst : DFF_X1 port map( D => n11087, CK => CLK, Q => 
                           n8738, QN => n1147);
   REGISTERS_reg_59_28_inst : DFF_X1 port map( D => n11088, CK => CLK, Q => 
                           n8739, QN => n1148);
   REGISTERS_reg_59_27_inst : DFF_X1 port map( D => n11089, CK => CLK, Q => 
                           n8740, QN => n1149);
   REGISTERS_reg_59_26_inst : DFF_X1 port map( D => n11090, CK => CLK, Q => 
                           n8741, QN => n1150);
   REGISTERS_reg_59_25_inst : DFF_X1 port map( D => n11091, CK => CLK, Q => 
                           n8742, QN => n1151);
   REGISTERS_reg_59_24_inst : DFF_X1 port map( D => n11092, CK => CLK, Q => 
                           n8743, QN => n1152);
   REGISTERS_reg_59_23_inst : DFF_X1 port map( D => n11093, CK => CLK, Q => 
                           n8744, QN => n1153);
   REGISTERS_reg_59_22_inst : DFF_X1 port map( D => n11094, CK => CLK, Q => 
                           n8745, QN => n1154);
   REGISTERS_reg_59_21_inst : DFF_X1 port map( D => n11095, CK => CLK, Q => 
                           n8746, QN => n1155);
   REGISTERS_reg_59_20_inst : DFF_X1 port map( D => n11096, CK => CLK, Q => 
                           n8747, QN => n1156);
   REGISTERS_reg_59_19_inst : DFF_X1 port map( D => n11097, CK => CLK, Q => 
                           n8748, QN => n1157);
   REGISTERS_reg_59_18_inst : DFF_X1 port map( D => n11098, CK => CLK, Q => 
                           n8749, QN => n1158);
   REGISTERS_reg_59_17_inst : DFF_X1 port map( D => n11099, CK => CLK, Q => 
                           n8750, QN => n1159);
   REGISTERS_reg_59_16_inst : DFF_X1 port map( D => n11100, CK => CLK, Q => 
                           n8751, QN => n1160);
   REGISTERS_reg_59_15_inst : DFF_X1 port map( D => n11101, CK => CLK, Q => 
                           n8752, QN => n1161);
   REGISTERS_reg_59_14_inst : DFF_X1 port map( D => n11102, CK => CLK, Q => 
                           n8753, QN => n1162);
   REGISTERS_reg_59_13_inst : DFF_X1 port map( D => n11103, CK => CLK, Q => 
                           n8754, QN => n1163);
   REGISTERS_reg_59_12_inst : DFF_X1 port map( D => n11104, CK => CLK, Q => 
                           n8755, QN => n1164);
   REGISTERS_reg_59_11_inst : DFF_X1 port map( D => n11105, CK => CLK, Q => 
                           n8756, QN => n1165);
   REGISTERS_reg_59_10_inst : DFF_X1 port map( D => n11106, CK => CLK, Q => 
                           n8757, QN => n1166);
   REGISTERS_reg_59_9_inst : DFF_X1 port map( D => n11107, CK => CLK, Q => 
                           n8758, QN => n1167);
   REGISTERS_reg_59_8_inst : DFF_X1 port map( D => n11108, CK => CLK, Q => 
                           n8759, QN => n1168);
   REGISTERS_reg_58_31_inst : DFF_X1 port map( D => n11053, CK => CLK, Q => 
                           n8704, QN => n1169);
   REGISTERS_reg_58_30_inst : DFF_X1 port map( D => n11054, CK => CLK, Q => 
                           n8705, QN => n1170);
   REGISTERS_reg_58_29_inst : DFF_X1 port map( D => n11055, CK => CLK, Q => 
                           n8706, QN => n1171);
   REGISTERS_reg_58_28_inst : DFF_X1 port map( D => n11056, CK => CLK, Q => 
                           n8707, QN => n1172);
   REGISTERS_reg_58_27_inst : DFF_X1 port map( D => n11057, CK => CLK, Q => 
                           n8708, QN => n1173);
   REGISTERS_reg_58_26_inst : DFF_X1 port map( D => n11058, CK => CLK, Q => 
                           n8709, QN => n1174);
   REGISTERS_reg_58_25_inst : DFF_X1 port map( D => n11059, CK => CLK, Q => 
                           n8710, QN => n1175);
   REGISTERS_reg_58_24_inst : DFF_X1 port map( D => n11060, CK => CLK, Q => 
                           n8711, QN => n1176);
   REGISTERS_reg_58_23_inst : DFF_X1 port map( D => n11061, CK => CLK, Q => 
                           n8712, QN => n1177);
   REGISTERS_reg_58_22_inst : DFF_X1 port map( D => n11062, CK => CLK, Q => 
                           n8713, QN => n1178);
   REGISTERS_reg_58_21_inst : DFF_X1 port map( D => n11063, CK => CLK, Q => 
                           n8714, QN => n1179);
   REGISTERS_reg_58_20_inst : DFF_X1 port map( D => n11064, CK => CLK, Q => 
                           n8715, QN => n1180);
   REGISTERS_reg_58_19_inst : DFF_X1 port map( D => n11065, CK => CLK, Q => 
                           n8716, QN => n1181);
   REGISTERS_reg_58_18_inst : DFF_X1 port map( D => n11066, CK => CLK, Q => 
                           n8717, QN => n1182);
   REGISTERS_reg_58_17_inst : DFF_X1 port map( D => n11067, CK => CLK, Q => 
                           n8718, QN => n1183);
   REGISTERS_reg_58_16_inst : DFF_X1 port map( D => n11068, CK => CLK, Q => 
                           n8719, QN => n1184);
   REGISTERS_reg_58_15_inst : DFF_X1 port map( D => n11069, CK => CLK, Q => 
                           n8720, QN => n1185);
   REGISTERS_reg_58_14_inst : DFF_X1 port map( D => n11070, CK => CLK, Q => 
                           n8721, QN => n1186);
   REGISTERS_reg_58_13_inst : DFF_X1 port map( D => n11071, CK => CLK, Q => 
                           n8722, QN => n1187);
   REGISTERS_reg_58_12_inst : DFF_X1 port map( D => n11072, CK => CLK, Q => 
                           n8723, QN => n1188);
   REGISTERS_reg_58_11_inst : DFF_X1 port map( D => n11073, CK => CLK, Q => 
                           n8724, QN => n1189);
   REGISTERS_reg_58_10_inst : DFF_X1 port map( D => n11074, CK => CLK, Q => 
                           n8725, QN => n1190);
   REGISTERS_reg_58_9_inst : DFF_X1 port map( D => n11075, CK => CLK, Q => 
                           n8726, QN => n1191);
   REGISTERS_reg_58_8_inst : DFF_X1 port map( D => n11076, CK => CLK, Q => 
                           n8727, QN => n1192);
   REGISTERS_reg_57_31_inst : DFF_X1 port map( D => n11021, CK => CLK, Q => 
                           n8672, QN => n1193);
   REGISTERS_reg_57_30_inst : DFF_X1 port map( D => n11022, CK => CLK, Q => 
                           n8673, QN => n1194);
   REGISTERS_reg_57_29_inst : DFF_X1 port map( D => n11023, CK => CLK, Q => 
                           n8674, QN => n1195);
   REGISTERS_reg_57_28_inst : DFF_X1 port map( D => n11024, CK => CLK, Q => 
                           n8675, QN => n1196);
   REGISTERS_reg_57_27_inst : DFF_X1 port map( D => n11025, CK => CLK, Q => 
                           n8676, QN => n1197);
   REGISTERS_reg_57_26_inst : DFF_X1 port map( D => n11026, CK => CLK, Q => 
                           n8677, QN => n1198);
   REGISTERS_reg_57_25_inst : DFF_X1 port map( D => n11027, CK => CLK, Q => 
                           n8678, QN => n1199);
   REGISTERS_reg_57_24_inst : DFF_X1 port map( D => n11028, CK => CLK, Q => 
                           n8679, QN => n1200);
   REGISTERS_reg_57_23_inst : DFF_X1 port map( D => n11029, CK => CLK, Q => 
                           n8680, QN => n1201);
   REGISTERS_reg_57_22_inst : DFF_X1 port map( D => n11030, CK => CLK, Q => 
                           n8681, QN => n1202);
   REGISTERS_reg_57_21_inst : DFF_X1 port map( D => n11031, CK => CLK, Q => 
                           n8682, QN => n1203);
   REGISTERS_reg_57_20_inst : DFF_X1 port map( D => n11032, CK => CLK, Q => 
                           n8683, QN => n1204);
   REGISTERS_reg_57_19_inst : DFF_X1 port map( D => n11033, CK => CLK, Q => 
                           n8684, QN => n1205);
   REGISTERS_reg_57_18_inst : DFF_X1 port map( D => n11034, CK => CLK, Q => 
                           n8685, QN => n1206);
   REGISTERS_reg_57_17_inst : DFF_X1 port map( D => n11035, CK => CLK, Q => 
                           n8686, QN => n1207);
   REGISTERS_reg_57_16_inst : DFF_X1 port map( D => n11036, CK => CLK, Q => 
                           n8687, QN => n1208);
   REGISTERS_reg_57_15_inst : DFF_X1 port map( D => n11037, CK => CLK, Q => 
                           n8688, QN => n1209);
   REGISTERS_reg_57_14_inst : DFF_X1 port map( D => n11038, CK => CLK, Q => 
                           n8689, QN => n1210);
   REGISTERS_reg_57_13_inst : DFF_X1 port map( D => n11039, CK => CLK, Q => 
                           n8690, QN => n1211);
   REGISTERS_reg_57_12_inst : DFF_X1 port map( D => n11040, CK => CLK, Q => 
                           n8691, QN => n1212);
   REGISTERS_reg_57_11_inst : DFF_X1 port map( D => n11041, CK => CLK, Q => 
                           n8692, QN => n1213);
   REGISTERS_reg_57_10_inst : DFF_X1 port map( D => n11042, CK => CLK, Q => 
                           n8693, QN => n1214);
   REGISTERS_reg_57_9_inst : DFF_X1 port map( D => n11043, CK => CLK, Q => 
                           n8694, QN => n1215);
   REGISTERS_reg_57_8_inst : DFF_X1 port map( D => n11044, CK => CLK, Q => 
                           n8695, QN => n1216);
   REGISTERS_reg_56_31_inst : DFF_X1 port map( D => n10989, CK => CLK, Q => 
                           n8640, QN => n1217);
   REGISTERS_reg_56_30_inst : DFF_X1 port map( D => n10990, CK => CLK, Q => 
                           n8641, QN => n1218);
   REGISTERS_reg_56_29_inst : DFF_X1 port map( D => n10991, CK => CLK, Q => 
                           n8642, QN => n1219);
   REGISTERS_reg_56_28_inst : DFF_X1 port map( D => n10992, CK => CLK, Q => 
                           n8643, QN => n1220);
   REGISTERS_reg_56_27_inst : DFF_X1 port map( D => n10993, CK => CLK, Q => 
                           n8644, QN => n1221);
   REGISTERS_reg_56_26_inst : DFF_X1 port map( D => n10994, CK => CLK, Q => 
                           n8645, QN => n1222);
   REGISTERS_reg_56_25_inst : DFF_X1 port map( D => n10995, CK => CLK, Q => 
                           n8646, QN => n1223);
   REGISTERS_reg_56_24_inst : DFF_X1 port map( D => n10996, CK => CLK, Q => 
                           n8647, QN => n1224);
   REGISTERS_reg_56_23_inst : DFF_X1 port map( D => n10997, CK => CLK, Q => 
                           n8648, QN => n1225);
   REGISTERS_reg_56_22_inst : DFF_X1 port map( D => n10998, CK => CLK, Q => 
                           n8649, QN => n1226);
   REGISTERS_reg_56_21_inst : DFF_X1 port map( D => n10999, CK => CLK, Q => 
                           n8650, QN => n1227);
   REGISTERS_reg_56_20_inst : DFF_X1 port map( D => n11000, CK => CLK, Q => 
                           n8651, QN => n1228);
   REGISTERS_reg_56_19_inst : DFF_X1 port map( D => n11001, CK => CLK, Q => 
                           n8652, QN => n1229);
   REGISTERS_reg_56_18_inst : DFF_X1 port map( D => n11002, CK => CLK, Q => 
                           n8653, QN => n1230);
   REGISTERS_reg_56_17_inst : DFF_X1 port map( D => n11003, CK => CLK, Q => 
                           n8654, QN => n1231);
   REGISTERS_reg_56_16_inst : DFF_X1 port map( D => n11004, CK => CLK, Q => 
                           n8655, QN => n1232);
   REGISTERS_reg_56_15_inst : DFF_X1 port map( D => n11005, CK => CLK, Q => 
                           n8656, QN => n1233);
   REGISTERS_reg_56_14_inst : DFF_X1 port map( D => n11006, CK => CLK, Q => 
                           n8657, QN => n1234);
   REGISTERS_reg_56_13_inst : DFF_X1 port map( D => n11007, CK => CLK, Q => 
                           n8658, QN => n1235);
   REGISTERS_reg_56_12_inst : DFF_X1 port map( D => n11008, CK => CLK, Q => 
                           n8659, QN => n1236);
   REGISTERS_reg_56_11_inst : DFF_X1 port map( D => n11009, CK => CLK, Q => 
                           n8660, QN => n1237);
   REGISTERS_reg_56_10_inst : DFF_X1 port map( D => n11010, CK => CLK, Q => 
                           n8661, QN => n1238);
   REGISTERS_reg_56_9_inst : DFF_X1 port map( D => n11011, CK => CLK, Q => 
                           n8662, QN => n1239);
   REGISTERS_reg_56_8_inst : DFF_X1 port map( D => n11012, CK => CLK, Q => 
                           n8663, QN => n1240);
   REGISTERS_reg_55_31_inst : DFF_X1 port map( D => n10957, CK => CLK, Q => 
                           n7535, QN => n1241);
   REGISTERS_reg_55_30_inst : DFF_X1 port map( D => n10958, CK => CLK, Q => 
                           n7533, QN => n1242);
   REGISTERS_reg_55_29_inst : DFF_X1 port map( D => n10959, CK => CLK, Q => 
                           n7531, QN => n1243);
   REGISTERS_reg_55_28_inst : DFF_X1 port map( D => n10960, CK => CLK, Q => 
                           n7530, QN => n1244);
   REGISTERS_reg_55_27_inst : DFF_X1 port map( D => n10961, CK => CLK, Q => 
                           n7529, QN => n1245);
   REGISTERS_reg_55_26_inst : DFF_X1 port map( D => n10962, CK => CLK, Q => 
                           n7527, QN => n1246);
   REGISTERS_reg_55_25_inst : DFF_X1 port map( D => n10963, CK => CLK, Q => 
                           n7525, QN => n1247);
   REGISTERS_reg_55_24_inst : DFF_X1 port map( D => n10964, CK => CLK, Q => 
                           n7524, QN => n1248);
   REGISTERS_reg_55_23_inst : DFF_X1 port map( D => n10965, CK => CLK, Q => 
                           n7523, QN => n1249);
   REGISTERS_reg_55_22_inst : DFF_X1 port map( D => n10966, CK => CLK, Q => 
                           n7521, QN => n1250);
   REGISTERS_reg_55_21_inst : DFF_X1 port map( D => n10967, CK => CLK, Q => 
                           n7519, QN => n1251);
   REGISTERS_reg_55_19_inst : DFF_X1 port map( D => n10969, CK => CLK, Q => 
                           n7517, QN => n1253);
   REGISTERS_reg_55_18_inst : DFF_X1 port map( D => n10970, CK => CLK, Q => 
                           n7515, QN => n1254);
   REGISTERS_reg_55_17_inst : DFF_X1 port map( D => n10971, CK => CLK, Q => 
                           n7513, QN => n1255);
   REGISTERS_reg_55_16_inst : DFF_X1 port map( D => n10972, CK => CLK, Q => 
                           n7512, QN => n1256);
   REGISTERS_reg_55_15_inst : DFF_X1 port map( D => n10973, CK => CLK, Q => 
                           n7511, QN => n1257);
   REGISTERS_reg_55_14_inst : DFF_X1 port map( D => n10974, CK => CLK, Q => 
                           n7509, QN => n1258);
   REGISTERS_reg_55_13_inst : DFF_X1 port map( D => n10975, CK => CLK, Q => 
                           n7507, QN => n1259);
   REGISTERS_reg_55_12_inst : DFF_X1 port map( D => n10976, CK => CLK, Q => 
                           n7506, QN => n1260);
   REGISTERS_reg_55_11_inst : DFF_X1 port map( D => n10977, CK => CLK, Q => 
                           n7505, QN => n1261);
   REGISTERS_reg_55_10_inst : DFF_X1 port map( D => n10978, CK => CLK, Q => 
                           n7503, QN => n1262);
   REGISTERS_reg_55_9_inst : DFF_X1 port map( D => n10979, CK => CLK, Q => 
                           n7501, QN => n1263);
   REGISTERS_reg_55_8_inst : DFF_X1 port map( D => n10980, CK => CLK, Q => 
                           n7500, QN => n1264);
   REGISTERS_reg_54_31_inst : DFF_X1 port map( D => n10925, CK => CLK, Q => 
                           n_1309, QN => n1265);
   REGISTERS_reg_54_30_inst : DFF_X1 port map( D => n10926, CK => CLK, Q => 
                           n_1310, QN => n1266);
   REGISTERS_reg_54_29_inst : DFF_X1 port map( D => n10927, CK => CLK, Q => 
                           n_1311, QN => n1267);
   REGISTERS_reg_54_28_inst : DFF_X1 port map( D => n10928, CK => CLK, Q => 
                           n_1312, QN => n1268);
   REGISTERS_reg_54_27_inst : DFF_X1 port map( D => n10929, CK => CLK, Q => 
                           n_1313, QN => n1269);
   REGISTERS_reg_54_26_inst : DFF_X1 port map( D => n10930, CK => CLK, Q => 
                           n_1314, QN => n1270);
   REGISTERS_reg_54_25_inst : DFF_X1 port map( D => n10931, CK => CLK, Q => 
                           n_1315, QN => n1271);
   REGISTERS_reg_54_24_inst : DFF_X1 port map( D => n10932, CK => CLK, Q => 
                           n_1316, QN => n1272);
   REGISTERS_reg_54_23_inst : DFF_X1 port map( D => n10933, CK => CLK, Q => 
                           n_1317, QN => n1273);
   REGISTERS_reg_54_22_inst : DFF_X1 port map( D => n10934, CK => CLK, Q => 
                           n_1318, QN => n1274);
   REGISTERS_reg_54_21_inst : DFF_X1 port map( D => n10935, CK => CLK, Q => 
                           n_1319, QN => n1275);
   REGISTERS_reg_54_20_inst : DFF_X1 port map( D => n10936, CK => CLK, Q => 
                           n_1320, QN => n1276);
   REGISTERS_reg_54_19_inst : DFF_X1 port map( D => n10937, CK => CLK, Q => 
                           n_1321, QN => n1277);
   REGISTERS_reg_54_18_inst : DFF_X1 port map( D => n10938, CK => CLK, Q => 
                           n_1322, QN => n1278);
   REGISTERS_reg_54_17_inst : DFF_X1 port map( D => n10939, CK => CLK, Q => 
                           n_1323, QN => n1279);
   REGISTERS_reg_54_16_inst : DFF_X1 port map( D => n10940, CK => CLK, Q => 
                           n_1324, QN => n1280);
   REGISTERS_reg_54_15_inst : DFF_X1 port map( D => n10941, CK => CLK, Q => 
                           n_1325, QN => n1281);
   REGISTERS_reg_54_14_inst : DFF_X1 port map( D => n10942, CK => CLK, Q => 
                           n_1326, QN => n1282);
   REGISTERS_reg_54_13_inst : DFF_X1 port map( D => n10943, CK => CLK, Q => 
                           n_1327, QN => n1283);
   REGISTERS_reg_54_12_inst : DFF_X1 port map( D => n10944, CK => CLK, Q => 
                           n_1328, QN => n1284);
   REGISTERS_reg_54_11_inst : DFF_X1 port map( D => n10945, CK => CLK, Q => 
                           n_1329, QN => n1285);
   REGISTERS_reg_54_10_inst : DFF_X1 port map( D => n10946, CK => CLK, Q => 
                           n_1330, QN => n1286);
   REGISTERS_reg_54_9_inst : DFF_X1 port map( D => n10947, CK => CLK, Q => 
                           n_1331, QN => n1287);
   REGISTERS_reg_54_8_inst : DFF_X1 port map( D => n10948, CK => CLK, Q => 
                           n_1332, QN => n1288);
   REGISTERS_reg_53_31_inst : DFF_X1 port map( D => n10893, CK => CLK, Q => 
                           n_1333, QN => n2067);
   REGISTERS_reg_53_30_inst : DFF_X1 port map( D => n10894, CK => CLK, Q => 
                           n_1334, QN => n2068);
   REGISTERS_reg_53_29_inst : DFF_X1 port map( D => n10895, CK => CLK, Q => 
                           n_1335, QN => n2069);
   REGISTERS_reg_53_28_inst : DFF_X1 port map( D => n10896, CK => CLK, Q => 
                           n_1336, QN => n2070);
   REGISTERS_reg_53_27_inst : DFF_X1 port map( D => n10897, CK => CLK, Q => 
                           n_1337, QN => n2071);
   REGISTERS_reg_53_26_inst : DFF_X1 port map( D => n10898, CK => CLK, Q => 
                           n_1338, QN => n2072);
   REGISTERS_reg_53_25_inst : DFF_X1 port map( D => n10899, CK => CLK, Q => 
                           n_1339, QN => n2073);
   REGISTERS_reg_53_24_inst : DFF_X1 port map( D => n10900, CK => CLK, Q => 
                           n_1340, QN => n2074);
   REGISTERS_reg_53_23_inst : DFF_X1 port map( D => n10901, CK => CLK, Q => 
                           n_1341, QN => n2075);
   REGISTERS_reg_53_22_inst : DFF_X1 port map( D => n10902, CK => CLK, Q => 
                           n_1342, QN => n2076);
   REGISTERS_reg_53_21_inst : DFF_X1 port map( D => n10903, CK => CLK, Q => 
                           n_1343, QN => n2077);
   REGISTERS_reg_53_20_inst : DFF_X1 port map( D => n10904, CK => CLK, Q => 
                           n_1344, QN => n2078);
   REGISTERS_reg_53_19_inst : DFF_X1 port map( D => n10905, CK => CLK, Q => 
                           n_1345, QN => n2079);
   REGISTERS_reg_53_18_inst : DFF_X1 port map( D => n10906, CK => CLK, Q => 
                           n_1346, QN => n2080);
   REGISTERS_reg_53_17_inst : DFF_X1 port map( D => n10907, CK => CLK, Q => 
                           n_1347, QN => n1289);
   REGISTERS_reg_53_16_inst : DFF_X1 port map( D => n10908, CK => CLK, Q => 
                           n_1348, QN => n1290);
   REGISTERS_reg_53_15_inst : DFF_X1 port map( D => n10909, CK => CLK, Q => 
                           n_1349, QN => n1291);
   REGISTERS_reg_53_14_inst : DFF_X1 port map( D => n10910, CK => CLK, Q => 
                           n_1350, QN => n1292);
   REGISTERS_reg_53_13_inst : DFF_X1 port map( D => n10911, CK => CLK, Q => 
                           n_1351, QN => n1293);
   REGISTERS_reg_52_31_inst : DFF_X1 port map( D => n10861, CK => CLK, Q => 
                           n_1352, QN => n2081);
   REGISTERS_reg_52_30_inst : DFF_X1 port map( D => n10862, CK => CLK, Q => 
                           n_1353, QN => n2082);
   REGISTERS_reg_52_29_inst : DFF_X1 port map( D => n10863, CK => CLK, Q => 
                           n_1354, QN => n2083);
   REGISTERS_reg_52_28_inst : DFF_X1 port map( D => n10864, CK => CLK, Q => 
                           n_1355, QN => n2084);
   REGISTERS_reg_52_27_inst : DFF_X1 port map( D => n10865, CK => CLK, Q => 
                           n_1356, QN => n2085);
   REGISTERS_reg_52_26_inst : DFF_X1 port map( D => n10866, CK => CLK, Q => 
                           n_1357, QN => n2086);
   REGISTERS_reg_52_25_inst : DFF_X1 port map( D => n10867, CK => CLK, Q => 
                           n_1358, QN => n2087);
   REGISTERS_reg_52_24_inst : DFF_X1 port map( D => n10868, CK => CLK, Q => 
                           n_1359, QN => n2088);
   REGISTERS_reg_52_23_inst : DFF_X1 port map( D => n10869, CK => CLK, Q => 
                           n_1360, QN => n2089);
   REGISTERS_reg_52_22_inst : DFF_X1 port map( D => n10870, CK => CLK, Q => 
                           n_1361, QN => n2090);
   REGISTERS_reg_52_21_inst : DFF_X1 port map( D => n10871, CK => CLK, Q => 
                           n_1362, QN => n2091);
   REGISTERS_reg_52_20_inst : DFF_X1 port map( D => n10872, CK => CLK, Q => 
                           n_1363, QN => n2092);
   REGISTERS_reg_52_19_inst : DFF_X1 port map( D => n10873, CK => CLK, Q => 
                           n_1364, QN => n2093);
   REGISTERS_reg_52_18_inst : DFF_X1 port map( D => n10874, CK => CLK, Q => 
                           n_1365, QN => n2094);
   REGISTERS_reg_52_17_inst : DFF_X1 port map( D => n10875, CK => CLK, Q => 
                           n_1366, QN => n1294);
   REGISTERS_reg_52_16_inst : DFF_X1 port map( D => n10876, CK => CLK, Q => 
                           n_1367, QN => n1295);
   REGISTERS_reg_52_15_inst : DFF_X1 port map( D => n10877, CK => CLK, Q => 
                           n_1368, QN => n1296);
   REGISTERS_reg_52_14_inst : DFF_X1 port map( D => n10878, CK => CLK, Q => 
                           n_1369, QN => n1297);
   REGISTERS_reg_52_13_inst : DFF_X1 port map( D => n10879, CK => CLK, Q => 
                           n_1370, QN => n1298);
   REGISTERS_reg_52_12_inst : DFF_X1 port map( D => n10880, CK => CLK, Q => 
                           n_1371, QN => n1299);
   REGISTERS_reg_52_11_inst : DFF_X1 port map( D => n10881, CK => CLK, Q => 
                           n_1372, QN => n1300);
   REGISTERS_reg_52_10_inst : DFF_X1 port map( D => n10882, CK => CLK, Q => 
                           n_1373, QN => n1301);
   REGISTERS_reg_52_9_inst : DFF_X1 port map( D => n10883, CK => CLK, Q => 
                           n_1374, QN => n1302);
   REGISTERS_reg_52_8_inst : DFF_X1 port map( D => n10884, CK => CLK, Q => 
                           n_1375, QN => n1303);
   REGISTERS_reg_51_20_inst : DFF_X1 port map( D => n10840, CK => CLK, Q => 
                           n784, QN => n2106);
   REGISTERS_reg_50_31_inst : DFF_X1 port map( D => n10797, CK => CLK, Q => 
                           n8608, QN => n1304);
   REGISTERS_reg_50_30_inst : DFF_X1 port map( D => n10798, CK => CLK, Q => 
                           n8609, QN => n1305);
   REGISTERS_reg_50_29_inst : DFF_X1 port map( D => n10799, CK => CLK, Q => 
                           n8610, QN => n1306);
   REGISTERS_reg_50_28_inst : DFF_X1 port map( D => n10800, CK => CLK, Q => 
                           n8611, QN => n1307);
   REGISTERS_reg_50_27_inst : DFF_X1 port map( D => n10801, CK => CLK, Q => 
                           n8612, QN => n1308);
   REGISTERS_reg_50_26_inst : DFF_X1 port map( D => n10802, CK => CLK, Q => 
                           n8613, QN => n1309);
   REGISTERS_reg_50_25_inst : DFF_X1 port map( D => n10803, CK => CLK, Q => 
                           n8614, QN => n1310);
   REGISTERS_reg_50_24_inst : DFF_X1 port map( D => n10804, CK => CLK, Q => 
                           n8615, QN => n1311);
   REGISTERS_reg_50_23_inst : DFF_X1 port map( D => n10805, CK => CLK, Q => 
                           n8616, QN => n1312);
   REGISTERS_reg_50_22_inst : DFF_X1 port map( D => n10806, CK => CLK, Q => 
                           n8617, QN => n1313);
   REGISTERS_reg_50_21_inst : DFF_X1 port map( D => n10807, CK => CLK, Q => 
                           n8618, QN => n1314);
   REGISTERS_reg_50_20_inst : DFF_X1 port map( D => n10808, CK => CLK, Q => 
                           n8619, QN => n1315);
   REGISTERS_reg_50_19_inst : DFF_X1 port map( D => n10809, CK => CLK, Q => 
                           n8620, QN => n1316);
   REGISTERS_reg_50_18_inst : DFF_X1 port map( D => n10810, CK => CLK, Q => 
                           n8621, QN => n1317);
   REGISTERS_reg_50_17_inst : DFF_X1 port map( D => n10811, CK => CLK, Q => 
                           n8622, QN => n1318);
   REGISTERS_reg_50_16_inst : DFF_X1 port map( D => n10812, CK => CLK, Q => 
                           n8623, QN => n1319);
   REGISTERS_reg_50_15_inst : DFF_X1 port map( D => n10813, CK => CLK, Q => 
                           n8624, QN => n1320);
   REGISTERS_reg_50_14_inst : DFF_X1 port map( D => n10814, CK => CLK, Q => 
                           n8625, QN => n1321);
   REGISTERS_reg_50_13_inst : DFF_X1 port map( D => n10815, CK => CLK, Q => 
                           n8626, QN => n1322);
   REGISTERS_reg_50_12_inst : DFF_X1 port map( D => n10816, CK => CLK, Q => 
                           n8627, QN => n1323);
   REGISTERS_reg_50_11_inst : DFF_X1 port map( D => n10817, CK => CLK, Q => 
                           n8628, QN => n1324);
   REGISTERS_reg_50_10_inst : DFF_X1 port map( D => n10818, CK => CLK, Q => 
                           n8629, QN => n1325);
   REGISTERS_reg_50_9_inst : DFF_X1 port map( D => n10819, CK => CLK, Q => 
                           n8630, QN => n1326);
   REGISTERS_reg_50_8_inst : DFF_X1 port map( D => n10820, CK => CLK, Q => 
                           n8631, QN => n1327);
   REGISTERS_reg_49_31_inst : DFF_X1 port map( D => n10765, CK => CLK, Q => 
                           n8576, QN => n1328);
   REGISTERS_reg_49_30_inst : DFF_X1 port map( D => n10766, CK => CLK, Q => 
                           n8577, QN => n1329);
   REGISTERS_reg_49_29_inst : DFF_X1 port map( D => n10767, CK => CLK, Q => 
                           n8578, QN => n1330);
   REGISTERS_reg_49_28_inst : DFF_X1 port map( D => n10768, CK => CLK, Q => 
                           n8579, QN => n1331);
   REGISTERS_reg_49_27_inst : DFF_X1 port map( D => n10769, CK => CLK, Q => 
                           n8580, QN => n1332);
   REGISTERS_reg_49_26_inst : DFF_X1 port map( D => n10770, CK => CLK, Q => 
                           n8581, QN => n1333);
   REGISTERS_reg_49_25_inst : DFF_X1 port map( D => n10771, CK => CLK, Q => 
                           n8582, QN => n1334);
   REGISTERS_reg_49_24_inst : DFF_X1 port map( D => n10772, CK => CLK, Q => 
                           n8583, QN => n1335);
   REGISTERS_reg_49_23_inst : DFF_X1 port map( D => n10773, CK => CLK, Q => 
                           n8584, QN => n1336);
   REGISTERS_reg_49_22_inst : DFF_X1 port map( D => n10774, CK => CLK, Q => 
                           n8585, QN => n1337);
   REGISTERS_reg_49_21_inst : DFF_X1 port map( D => n10775, CK => CLK, Q => 
                           n8586, QN => n1338);
   REGISTERS_reg_49_20_inst : DFF_X1 port map( D => n10776, CK => CLK, Q => 
                           n8587, QN => n1339);
   REGISTERS_reg_49_19_inst : DFF_X1 port map( D => n10777, CK => CLK, Q => 
                           n8588, QN => n1340);
   REGISTERS_reg_49_18_inst : DFF_X1 port map( D => n10778, CK => CLK, Q => 
                           n8589, QN => n1341);
   REGISTERS_reg_49_17_inst : DFF_X1 port map( D => n10779, CK => CLK, Q => 
                           n8590, QN => n1342);
   REGISTERS_reg_49_16_inst : DFF_X1 port map( D => n10780, CK => CLK, Q => 
                           n8591, QN => n1343);
   REGISTERS_reg_49_15_inst : DFF_X1 port map( D => n10781, CK => CLK, Q => 
                           n8592, QN => n1344);
   REGISTERS_reg_49_14_inst : DFF_X1 port map( D => n10782, CK => CLK, Q => 
                           n8593, QN => n1345);
   REGISTERS_reg_49_13_inst : DFF_X1 port map( D => n10783, CK => CLK, Q => 
                           n8594, QN => n1346);
   REGISTERS_reg_49_12_inst : DFF_X1 port map( D => n10784, CK => CLK, Q => 
                           n8595, QN => n1347);
   REGISTERS_reg_49_11_inst : DFF_X1 port map( D => n10785, CK => CLK, Q => 
                           n8596, QN => n1348);
   REGISTERS_reg_49_10_inst : DFF_X1 port map( D => n10786, CK => CLK, Q => 
                           n8597, QN => n1349);
   REGISTERS_reg_49_9_inst : DFF_X1 port map( D => n10787, CK => CLK, Q => 
                           n8598, QN => n1350);
   REGISTERS_reg_49_8_inst : DFF_X1 port map( D => n10788, CK => CLK, Q => 
                           n8599, QN => n1351);
   REGISTERS_reg_48_31_inst : DFF_X1 port map( D => n10733, CK => CLK, Q => 
                           n_1376, QN => n1352);
   REGISTERS_reg_48_30_inst : DFF_X1 port map( D => n10734, CK => CLK, Q => 
                           n_1377, QN => n1353);
   REGISTERS_reg_48_29_inst : DFF_X1 port map( D => n10735, CK => CLK, Q => 
                           n_1378, QN => n1354);
   REGISTERS_reg_48_28_inst : DFF_X1 port map( D => n10736, CK => CLK, Q => 
                           n_1379, QN => n1355);
   REGISTERS_reg_48_27_inst : DFF_X1 port map( D => n10737, CK => CLK, Q => 
                           n_1380, QN => n1356);
   REGISTERS_reg_48_26_inst : DFF_X1 port map( D => n10738, CK => CLK, Q => 
                           n_1381, QN => n1357);
   REGISTERS_reg_48_25_inst : DFF_X1 port map( D => n10739, CK => CLK, Q => 
                           n_1382, QN => n1358);
   REGISTERS_reg_48_24_inst : DFF_X1 port map( D => n10740, CK => CLK, Q => 
                           n_1383, QN => n1359);
   REGISTERS_reg_48_23_inst : DFF_X1 port map( D => n10741, CK => CLK, Q => 
                           n_1384, QN => n1360);
   REGISTERS_reg_48_22_inst : DFF_X1 port map( D => n10742, CK => CLK, Q => 
                           n_1385, QN => n1361);
   REGISTERS_reg_48_21_inst : DFF_X1 port map( D => n10743, CK => CLK, Q => 
                           n_1386, QN => n1362);
   REGISTERS_reg_48_20_inst : DFF_X1 port map( D => n10744, CK => CLK, Q => 
                           n_1387, QN => n1363);
   REGISTERS_reg_48_19_inst : DFF_X1 port map( D => n10745, CK => CLK, Q => 
                           n_1388, QN => n1364);
   REGISTERS_reg_48_18_inst : DFF_X1 port map( D => n10746, CK => CLK, Q => 
                           n_1389, QN => n1365);
   REGISTERS_reg_48_17_inst : DFF_X1 port map( D => n10747, CK => CLK, Q => 
                           n_1390, QN => n1366);
   REGISTERS_reg_48_16_inst : DFF_X1 port map( D => n10748, CK => CLK, Q => 
                           n_1391, QN => n1367);
   REGISTERS_reg_48_15_inst : DFF_X1 port map( D => n10749, CK => CLK, Q => 
                           n_1392, QN => n1368);
   REGISTERS_reg_48_14_inst : DFF_X1 port map( D => n10750, CK => CLK, Q => 
                           n_1393, QN => n1369);
   REGISTERS_reg_48_13_inst : DFF_X1 port map( D => n10751, CK => CLK, Q => 
                           n_1394, QN => n1370);
   REGISTERS_reg_48_12_inst : DFF_X1 port map( D => n10752, CK => CLK, Q => 
                           n_1395, QN => n1371);
   REGISTERS_reg_48_11_inst : DFF_X1 port map( D => n10753, CK => CLK, Q => 
                           n_1396, QN => n1372);
   REGISTERS_reg_48_10_inst : DFF_X1 port map( D => n10754, CK => CLK, Q => 
                           n_1397, QN => n1373);
   REGISTERS_reg_48_9_inst : DFF_X1 port map( D => n10755, CK => CLK, Q => 
                           n_1398, QN => n1374);
   REGISTERS_reg_48_8_inst : DFF_X1 port map( D => n10756, CK => CLK, Q => 
                           n_1399, QN => n1375);
   REGISTERS_reg_47_31_inst : DFF_X1 port map( D => n10701, CK => CLK, Q => 
                           n_1400, QN => n1376);
   REGISTERS_reg_47_30_inst : DFF_X1 port map( D => n10702, CK => CLK, Q => 
                           n_1401, QN => n1377);
   REGISTERS_reg_47_29_inst : DFF_X1 port map( D => n10703, CK => CLK, Q => 
                           n_1402, QN => n1378);
   REGISTERS_reg_47_28_inst : DFF_X1 port map( D => n10704, CK => CLK, Q => 
                           n_1403, QN => n1379);
   REGISTERS_reg_47_27_inst : DFF_X1 port map( D => n10705, CK => CLK, Q => 
                           n_1404, QN => n1380);
   REGISTERS_reg_47_26_inst : DFF_X1 port map( D => n10706, CK => CLK, Q => 
                           n_1405, QN => n1381);
   REGISTERS_reg_47_25_inst : DFF_X1 port map( D => n10707, CK => CLK, Q => 
                           n_1406, QN => n1382);
   REGISTERS_reg_47_24_inst : DFF_X1 port map( D => n10708, CK => CLK, Q => 
                           n_1407, QN => n1383);
   REGISTERS_reg_47_23_inst : DFF_X1 port map( D => n10709, CK => CLK, Q => 
                           n_1408, QN => n1384);
   REGISTERS_reg_47_22_inst : DFF_X1 port map( D => n10710, CK => CLK, Q => 
                           n_1409, QN => n1385);
   REGISTERS_reg_47_21_inst : DFF_X1 port map( D => n10711, CK => CLK, Q => 
                           n_1410, QN => n1386);
   REGISTERS_reg_47_20_inst : DFF_X1 port map( D => n10712, CK => CLK, Q => 
                           n_1411, QN => n1387);
   REGISTERS_reg_47_19_inst : DFF_X1 port map( D => n10713, CK => CLK, Q => 
                           n_1412, QN => n1388);
   REGISTERS_reg_47_18_inst : DFF_X1 port map( D => n10714, CK => CLK, Q => 
                           n_1413, QN => n1389);
   REGISTERS_reg_47_17_inst : DFF_X1 port map( D => n10715, CK => CLK, Q => 
                           n_1414, QN => n1390);
   REGISTERS_reg_47_16_inst : DFF_X1 port map( D => n10716, CK => CLK, Q => 
                           n_1415, QN => n1391);
   REGISTERS_reg_47_15_inst : DFF_X1 port map( D => n10717, CK => CLK, Q => 
                           n_1416, QN => n1392);
   REGISTERS_reg_47_14_inst : DFF_X1 port map( D => n10718, CK => CLK, Q => 
                           n_1417, QN => n1393);
   REGISTERS_reg_47_13_inst : DFF_X1 port map( D => n10719, CK => CLK, Q => 
                           n_1418, QN => n1394);
   REGISTERS_reg_47_12_inst : DFF_X1 port map( D => n10720, CK => CLK, Q => 
                           n_1419, QN => n1395);
   REGISTERS_reg_47_11_inst : DFF_X1 port map( D => n10721, CK => CLK, Q => 
                           n_1420, QN => n1396);
   REGISTERS_reg_47_10_inst : DFF_X1 port map( D => n10722, CK => CLK, Q => 
                           n_1421, QN => n1397);
   REGISTERS_reg_47_9_inst : DFF_X1 port map( D => n10723, CK => CLK, Q => 
                           n_1422, QN => n1398);
   REGISTERS_reg_47_8_inst : DFF_X1 port map( D => n10724, CK => CLK, Q => 
                           n_1423, QN => n1399);
   REGISTERS_reg_46_31_inst : DFF_X1 port map( D => n10669, CK => CLK, Q => 
                           n8482, QN => n1400);
   REGISTERS_reg_46_30_inst : DFF_X1 port map( D => n10670, CK => CLK, Q => 
                           n8483, QN => n1401);
   REGISTERS_reg_46_29_inst : DFF_X1 port map( D => n10671, CK => CLK, Q => 
                           n8484, QN => n1402);
   REGISTERS_reg_46_28_inst : DFF_X1 port map( D => n10672, CK => CLK, Q => 
                           n8485, QN => n1403);
   REGISTERS_reg_46_27_inst : DFF_X1 port map( D => n10673, CK => CLK, Q => 
                           n8486, QN => n1404);
   REGISTERS_reg_46_26_inst : DFF_X1 port map( D => n10674, CK => CLK, Q => 
                           n8487, QN => n1405);
   REGISTERS_reg_46_25_inst : DFF_X1 port map( D => n10675, CK => CLK, Q => 
                           n8488, QN => n1406);
   REGISTERS_reg_46_24_inst : DFF_X1 port map( D => n10676, CK => CLK, Q => 
                           n8489, QN => n1407);
   REGISTERS_reg_46_23_inst : DFF_X1 port map( D => n10677, CK => CLK, Q => 
                           n8490, QN => n1408);
   REGISTERS_reg_46_22_inst : DFF_X1 port map( D => n10678, CK => CLK, Q => 
                           n8491, QN => n1409);
   REGISTERS_reg_46_21_inst : DFF_X1 port map( D => n10679, CK => CLK, Q => 
                           n8492, QN => n1410);
   REGISTERS_reg_46_20_inst : DFF_X1 port map( D => n10680, CK => CLK, Q => 
                           n8493, QN => n1411);
   REGISTERS_reg_46_19_inst : DFF_X1 port map( D => n10681, CK => CLK, Q => 
                           n8494, QN => n1412);
   REGISTERS_reg_46_18_inst : DFF_X1 port map( D => n10682, CK => CLK, Q => 
                           n8495, QN => n1413);
   REGISTERS_reg_46_17_inst : DFF_X1 port map( D => n10683, CK => CLK, Q => 
                           n8496, QN => n1414);
   REGISTERS_reg_46_16_inst : DFF_X1 port map( D => n10684, CK => CLK, Q => 
                           n8497, QN => n1415);
   REGISTERS_reg_46_15_inst : DFF_X1 port map( D => n10685, CK => CLK, Q => 
                           n8498, QN => n1416);
   REGISTERS_reg_46_14_inst : DFF_X1 port map( D => n10686, CK => CLK, Q => 
                           n8499, QN => n1417);
   REGISTERS_reg_46_13_inst : DFF_X1 port map( D => n10687, CK => CLK, Q => 
                           n8500, QN => n1418);
   REGISTERS_reg_46_12_inst : DFF_X1 port map( D => n10688, CK => CLK, Q => 
                           n8501, QN => n1419);
   REGISTERS_reg_46_11_inst : DFF_X1 port map( D => n10689, CK => CLK, Q => 
                           n8502, QN => n1420);
   REGISTERS_reg_46_10_inst : DFF_X1 port map( D => n10690, CK => CLK, Q => 
                           n8503, QN => n1421);
   REGISTERS_reg_46_9_inst : DFF_X1 port map( D => n10691, CK => CLK, Q => 
                           n8504, QN => n1422);
   REGISTERS_reg_46_8_inst : DFF_X1 port map( D => n10692, CK => CLK, Q => 
                           n8505, QN => n1423);
   REGISTERS_reg_45_31_inst : DFF_X1 port map( D => n10637, CK => CLK, Q => 
                           n8450, QN => n1424);
   REGISTERS_reg_45_30_inst : DFF_X1 port map( D => n10638, CK => CLK, Q => 
                           n8451, QN => n1425);
   REGISTERS_reg_45_29_inst : DFF_X1 port map( D => n10639, CK => CLK, Q => 
                           n8452, QN => n1426);
   REGISTERS_reg_45_28_inst : DFF_X1 port map( D => n10640, CK => CLK, Q => 
                           n8453, QN => n1427);
   REGISTERS_reg_45_27_inst : DFF_X1 port map( D => n10641, CK => CLK, Q => 
                           n8454, QN => n1428);
   REGISTERS_reg_45_26_inst : DFF_X1 port map( D => n10642, CK => CLK, Q => 
                           n8455, QN => n1429);
   REGISTERS_reg_45_25_inst : DFF_X1 port map( D => n10643, CK => CLK, Q => 
                           n8456, QN => n1430);
   REGISTERS_reg_45_24_inst : DFF_X1 port map( D => n10644, CK => CLK, Q => 
                           n8457, QN => n1431);
   REGISTERS_reg_45_23_inst : DFF_X1 port map( D => n10645, CK => CLK, Q => 
                           n8458, QN => n1432);
   REGISTERS_reg_45_22_inst : DFF_X1 port map( D => n10646, CK => CLK, Q => 
                           n8459, QN => n1433);
   REGISTERS_reg_45_21_inst : DFF_X1 port map( D => n10647, CK => CLK, Q => 
                           n8460, QN => n1434);
   REGISTERS_reg_45_20_inst : DFF_X1 port map( D => n10648, CK => CLK, Q => 
                           n8461, QN => n1435);
   REGISTERS_reg_45_19_inst : DFF_X1 port map( D => n10649, CK => CLK, Q => 
                           n8462, QN => n1436);
   REGISTERS_reg_45_18_inst : DFF_X1 port map( D => n10650, CK => CLK, Q => 
                           n8463, QN => n1437);
   REGISTERS_reg_45_17_inst : DFF_X1 port map( D => n10651, CK => CLK, Q => 
                           n8464, QN => n1438);
   REGISTERS_reg_45_16_inst : DFF_X1 port map( D => n10652, CK => CLK, Q => 
                           n8465, QN => n1439);
   REGISTERS_reg_45_15_inst : DFF_X1 port map( D => n10653, CK => CLK, Q => 
                           n8466, QN => n1440);
   REGISTERS_reg_45_14_inst : DFF_X1 port map( D => n10654, CK => CLK, Q => 
                           n8467, QN => n1441);
   REGISTERS_reg_45_13_inst : DFF_X1 port map( D => n10655, CK => CLK, Q => 
                           n8468, QN => n1442);
   REGISTERS_reg_45_12_inst : DFF_X1 port map( D => n10656, CK => CLK, Q => 
                           n8469, QN => n1443);
   REGISTERS_reg_45_11_inst : DFF_X1 port map( D => n10657, CK => CLK, Q => 
                           n8470, QN => n1444);
   REGISTERS_reg_45_10_inst : DFF_X1 port map( D => n10658, CK => CLK, Q => 
                           n8471, QN => n1445);
   REGISTERS_reg_45_9_inst : DFF_X1 port map( D => n10659, CK => CLK, Q => 
                           n8472, QN => n1446);
   REGISTERS_reg_45_8_inst : DFF_X1 port map( D => n10660, CK => CLK, Q => 
                           n8473, QN => n1447);
   REGISTERS_reg_44_31_inst : DFF_X1 port map( D => n10605, CK => CLK, Q => 
                           n_1424, QN => n2119);
   REGISTERS_reg_44_30_inst : DFF_X1 port map( D => n10606, CK => CLK, Q => 
                           n_1425, QN => n2120);
   REGISTERS_reg_44_29_inst : DFF_X1 port map( D => n10607, CK => CLK, Q => 
                           n_1426, QN => n2121);
   REGISTERS_reg_44_28_inst : DFF_X1 port map( D => n10608, CK => CLK, Q => 
                           n_1427, QN => n2122);
   REGISTERS_reg_44_27_inst : DFF_X1 port map( D => n10609, CK => CLK, Q => 
                           n_1428, QN => n2123);
   REGISTERS_reg_44_26_inst : DFF_X1 port map( D => n10610, CK => CLK, Q => 
                           n_1429, QN => n2124);
   REGISTERS_reg_44_25_inst : DFF_X1 port map( D => n10611, CK => CLK, Q => 
                           n_1430, QN => n2125);
   REGISTERS_reg_44_24_inst : DFF_X1 port map( D => n10612, CK => CLK, Q => 
                           n_1431, QN => n2126);
   REGISTERS_reg_44_23_inst : DFF_X1 port map( D => n10613, CK => CLK, Q => 
                           n_1432, QN => n2127);
   REGISTERS_reg_44_22_inst : DFF_X1 port map( D => n10614, CK => CLK, Q => 
                           n_1433, QN => n2128);
   REGISTERS_reg_44_21_inst : DFF_X1 port map( D => n10615, CK => CLK, Q => 
                           n_1434, QN => n2129);
   REGISTERS_reg_44_20_inst : DFF_X1 port map( D => n10616, CK => CLK, Q => 
                           n_1435, QN => n2130);
   REGISTERS_reg_44_19_inst : DFF_X1 port map( D => n10617, CK => CLK, Q => 
                           n_1436, QN => n2131);
   REGISTERS_reg_44_18_inst : DFF_X1 port map( D => n10618, CK => CLK, Q => 
                           n_1437, QN => n2132);
   REGISTERS_reg_44_17_inst : DFF_X1 port map( D => n10619, CK => CLK, Q => 
                           n_1438, QN => n1448);
   REGISTERS_reg_44_16_inst : DFF_X1 port map( D => n10620, CK => CLK, Q => 
                           n_1439, QN => n1449);
   REGISTERS_reg_44_15_inst : DFF_X1 port map( D => n10621, CK => CLK, Q => 
                           n_1440, QN => n1450);
   REGISTERS_reg_44_14_inst : DFF_X1 port map( D => n10622, CK => CLK, Q => 
                           n_1441, QN => n1451);
   REGISTERS_reg_44_13_inst : DFF_X1 port map( D => n10623, CK => CLK, Q => 
                           n_1442, QN => n1452);
   REGISTERS_reg_44_12_inst : DFF_X1 port map( D => n10624, CK => CLK, Q => 
                           n_1443, QN => n2133);
   REGISTERS_reg_44_11_inst : DFF_X1 port map( D => n10625, CK => CLK, Q => 
                           n_1444, QN => n2134);
   REGISTERS_reg_44_10_inst : DFF_X1 port map( D => n10626, CK => CLK, Q => 
                           n_1445, QN => n2135);
   REGISTERS_reg_44_9_inst : DFF_X1 port map( D => n10627, CK => CLK, Q => 
                           n_1446, QN => n2136);
   REGISTERS_reg_44_8_inst : DFF_X1 port map( D => n10628, CK => CLK, Q => 
                           n_1447, QN => n2137);
   REGISTERS_reg_43_31_inst : DFF_X1 port map( D => n10573, CK => CLK, Q => 
                           n_1448, QN => n2138);
   REGISTERS_reg_43_30_inst : DFF_X1 port map( D => n10574, CK => CLK, Q => 
                           n_1449, QN => n2139);
   REGISTERS_reg_43_29_inst : DFF_X1 port map( D => n10575, CK => CLK, Q => 
                           n_1450, QN => n2140);
   REGISTERS_reg_43_28_inst : DFF_X1 port map( D => n10576, CK => CLK, Q => 
                           n_1451, QN => n2141);
   REGISTERS_reg_43_27_inst : DFF_X1 port map( D => n10577, CK => CLK, Q => 
                           n_1452, QN => n2142);
   REGISTERS_reg_43_26_inst : DFF_X1 port map( D => n10578, CK => CLK, Q => 
                           n_1453, QN => n2143);
   REGISTERS_reg_43_25_inst : DFF_X1 port map( D => n10579, CK => CLK, Q => 
                           n_1454, QN => n2144);
   REGISTERS_reg_43_24_inst : DFF_X1 port map( D => n10580, CK => CLK, Q => 
                           n_1455, QN => n2145);
   REGISTERS_reg_43_23_inst : DFF_X1 port map( D => n10581, CK => CLK, Q => 
                           n_1456, QN => n2146);
   REGISTERS_reg_43_22_inst : DFF_X1 port map( D => n10582, CK => CLK, Q => 
                           n_1457, QN => n2147);
   REGISTERS_reg_43_21_inst : DFF_X1 port map( D => n10583, CK => CLK, Q => 
                           n_1458, QN => n2148);
   REGISTERS_reg_43_20_inst : DFF_X1 port map( D => n10584, CK => CLK, Q => 
                           n_1459, QN => n2149);
   REGISTERS_reg_43_19_inst : DFF_X1 port map( D => n10585, CK => CLK, Q => 
                           n_1460, QN => n2278);
   REGISTERS_reg_43_18_inst : DFF_X1 port map( D => n10586, CK => CLK, Q => 
                           n_1461, QN => n2279);
   REGISTERS_reg_43_17_inst : DFF_X1 port map( D => n10587, CK => CLK, Q => 
                           n_1462, QN => n1453);
   REGISTERS_reg_43_16_inst : DFF_X1 port map( D => n10588, CK => CLK, Q => 
                           n_1463, QN => n1454);
   REGISTERS_reg_43_15_inst : DFF_X1 port map( D => n10589, CK => CLK, Q => 
                           n_1464, QN => n1455);
   REGISTERS_reg_43_14_inst : DFF_X1 port map( D => n10590, CK => CLK, Q => 
                           n_1465, QN => n1456);
   REGISTERS_reg_43_13_inst : DFF_X1 port map( D => n10591, CK => CLK, Q => 
                           n_1466, QN => n1457);
   REGISTERS_reg_43_12_inst : DFF_X1 port map( D => n10592, CK => CLK, Q => 
                           n_1467, QN => n1458);
   REGISTERS_reg_43_11_inst : DFF_X1 port map( D => n10593, CK => CLK, Q => 
                           n_1468, QN => n1459);
   REGISTERS_reg_43_10_inst : DFF_X1 port map( D => n10594, CK => CLK, Q => 
                           n_1469, QN => n1460);
   REGISTERS_reg_43_9_inst : DFF_X1 port map( D => n10595, CK => CLK, Q => 
                           n_1470, QN => n1461);
   REGISTERS_reg_43_8_inst : DFF_X1 port map( D => n10596, CK => CLK, Q => 
                           n_1471, QN => n1462);
   REGISTERS_reg_42_20_inst : DFF_X1 port map( D => n10552, CK => CLK, Q => 
                           n777, QN => n2291);
   REGISTERS_reg_41_31_inst : DFF_X1 port map( D => n10509, CK => CLK, Q => 
                           n8418, QN => n1463);
   REGISTERS_reg_41_30_inst : DFF_X1 port map( D => n10510, CK => CLK, Q => 
                           n8419, QN => n1464);
   REGISTERS_reg_41_29_inst : DFF_X1 port map( D => n10511, CK => CLK, Q => 
                           n8420, QN => n1465);
   REGISTERS_reg_41_28_inst : DFF_X1 port map( D => n10512, CK => CLK, Q => 
                           n8421, QN => n1466);
   REGISTERS_reg_41_27_inst : DFF_X1 port map( D => n10513, CK => CLK, Q => 
                           n8422, QN => n1467);
   REGISTERS_reg_41_26_inst : DFF_X1 port map( D => n10514, CK => CLK, Q => 
                           n8423, QN => n1468);
   REGISTERS_reg_41_25_inst : DFF_X1 port map( D => n10515, CK => CLK, Q => 
                           n8424, QN => n1469);
   REGISTERS_reg_41_24_inst : DFF_X1 port map( D => n10516, CK => CLK, Q => 
                           n8425, QN => n1470);
   REGISTERS_reg_41_23_inst : DFF_X1 port map( D => n10517, CK => CLK, Q => 
                           n8426, QN => n1471);
   REGISTERS_reg_41_22_inst : DFF_X1 port map( D => n10518, CK => CLK, Q => 
                           n8427, QN => n1472);
   REGISTERS_reg_41_21_inst : DFF_X1 port map( D => n10519, CK => CLK, Q => 
                           n8428, QN => n1473);
   REGISTERS_reg_41_20_inst : DFF_X1 port map( D => n10520, CK => CLK, Q => 
                           n8429, QN => n1474);
   REGISTERS_reg_41_19_inst : DFF_X1 port map( D => n10521, CK => CLK, Q => 
                           n8430, QN => n1475);
   REGISTERS_reg_41_18_inst : DFF_X1 port map( D => n10522, CK => CLK, Q => 
                           n8431, QN => n1476);
   REGISTERS_reg_41_17_inst : DFF_X1 port map( D => n10523, CK => CLK, Q => 
                           n8432, QN => n1477);
   REGISTERS_reg_41_16_inst : DFF_X1 port map( D => n10524, CK => CLK, Q => 
                           n8433, QN => n1478);
   REGISTERS_reg_41_15_inst : DFF_X1 port map( D => n10525, CK => CLK, Q => 
                           n8434, QN => n1479);
   REGISTERS_reg_41_14_inst : DFF_X1 port map( D => n10526, CK => CLK, Q => 
                           n8435, QN => n1480);
   REGISTERS_reg_41_13_inst : DFF_X1 port map( D => n10527, CK => CLK, Q => 
                           n8436, QN => n1481);
   REGISTERS_reg_41_12_inst : DFF_X1 port map( D => n10528, CK => CLK, Q => 
                           n8437, QN => n1482);
   REGISTERS_reg_41_11_inst : DFF_X1 port map( D => n10529, CK => CLK, Q => 
                           n8438, QN => n1483);
   REGISTERS_reg_41_10_inst : DFF_X1 port map( D => n10530, CK => CLK, Q => 
                           n8439, QN => n1484);
   REGISTERS_reg_41_9_inst : DFF_X1 port map( D => n10531, CK => CLK, Q => 
                           n8440, QN => n1485);
   REGISTERS_reg_41_8_inst : DFF_X1 port map( D => n10532, CK => CLK, Q => 
                           n8441, QN => n1486);
   REGISTERS_reg_40_31_inst : DFF_X1 port map( D => n10477, CK => CLK, Q => 
                           n8386, QN => n1487);
   REGISTERS_reg_40_30_inst : DFF_X1 port map( D => n10478, CK => CLK, Q => 
                           n8387, QN => n1488);
   REGISTERS_reg_40_29_inst : DFF_X1 port map( D => n10479, CK => CLK, Q => 
                           n8388, QN => n1489);
   REGISTERS_reg_40_28_inst : DFF_X1 port map( D => n10480, CK => CLK, Q => 
                           n8389, QN => n1490);
   REGISTERS_reg_40_27_inst : DFF_X1 port map( D => n10481, CK => CLK, Q => 
                           n8390, QN => n1491);
   REGISTERS_reg_40_26_inst : DFF_X1 port map( D => n10482, CK => CLK, Q => 
                           n8391, QN => n1492);
   REGISTERS_reg_40_25_inst : DFF_X1 port map( D => n10483, CK => CLK, Q => 
                           n8392, QN => n1493);
   REGISTERS_reg_40_24_inst : DFF_X1 port map( D => n10484, CK => CLK, Q => 
                           n8393, QN => n1494);
   REGISTERS_reg_40_23_inst : DFF_X1 port map( D => n10485, CK => CLK, Q => 
                           n8394, QN => n1495);
   REGISTERS_reg_40_22_inst : DFF_X1 port map( D => n10486, CK => CLK, Q => 
                           n8395, QN => n1496);
   REGISTERS_reg_40_21_inst : DFF_X1 port map( D => n10487, CK => CLK, Q => 
                           n8396, QN => n1497);
   REGISTERS_reg_40_20_inst : DFF_X1 port map( D => n10488, CK => CLK, Q => 
                           n8397, QN => n1498);
   REGISTERS_reg_40_19_inst : DFF_X1 port map( D => n10489, CK => CLK, Q => 
                           n8398, QN => n1499);
   REGISTERS_reg_40_18_inst : DFF_X1 port map( D => n10490, CK => CLK, Q => 
                           n8399, QN => n1500);
   REGISTERS_reg_40_17_inst : DFF_X1 port map( D => n10491, CK => CLK, Q => 
                           n8400, QN => n1501);
   REGISTERS_reg_40_16_inst : DFF_X1 port map( D => n10492, CK => CLK, Q => 
                           n8401, QN => n1502);
   REGISTERS_reg_40_15_inst : DFF_X1 port map( D => n10493, CK => CLK, Q => 
                           n8402, QN => n1503);
   REGISTERS_reg_40_14_inst : DFF_X1 port map( D => n10494, CK => CLK, Q => 
                           n8403, QN => n1504);
   REGISTERS_reg_40_13_inst : DFF_X1 port map( D => n10495, CK => CLK, Q => 
                           n8404, QN => n1505);
   REGISTERS_reg_40_12_inst : DFF_X1 port map( D => n10496, CK => CLK, Q => 
                           n8405, QN => n1506);
   REGISTERS_reg_40_11_inst : DFF_X1 port map( D => n10497, CK => CLK, Q => 
                           n8406, QN => n1507);
   REGISTERS_reg_40_10_inst : DFF_X1 port map( D => n10498, CK => CLK, Q => 
                           n8407, QN => n1508);
   REGISTERS_reg_40_9_inst : DFF_X1 port map( D => n10499, CK => CLK, Q => 
                           n8408, QN => n1509);
   REGISTERS_reg_40_8_inst : DFF_X1 port map( D => n10500, CK => CLK, Q => 
                           n8409, QN => n1510);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n10445, CK => CLK, Q => 
                           n831, QN => n1511);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n10456, CK => CLK, Q => 
                           n774, QN => n2314);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n10381, CK => CLK, Q => 
                           n8354, QN => n1512);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n10382, CK => CLK, Q => 
                           n_1472, QN => n1513);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n10383, CK => CLK, Q => 
                           n_1473, QN => n1514);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n10384, CK => CLK, Q => 
                           n_1474, QN => n1515);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n10385, CK => CLK, Q => 
                           n_1475, QN => n1516);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n10386, CK => CLK, Q => 
                           n_1476, QN => n1517);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n10387, CK => CLK, Q => 
                           n_1477, QN => n1518);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n10388, CK => CLK, Q => 
                           n_1478, QN => n1519);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n10389, CK => CLK, Q => 
                           n_1479, QN => n1520);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n10390, CK => CLK, Q => 
                           n_1480, QN => n1521);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n10391, CK => CLK, Q => 
                           n_1481, QN => n1522);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n10392, CK => CLK, Q => 
                           n_1482, QN => n1523);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n10393, CK => CLK, Q => 
                           n_1483, QN => n1524);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n10394, CK => CLK, Q => 
                           n_1484, QN => n1525);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n10395, CK => CLK, Q => 
                           n_1485, QN => n1526);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n10396, CK => CLK, Q => 
                           n_1486, QN => n1527);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n10397, CK => CLK, Q => 
                           n_1487, QN => n1528);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n10398, CK => CLK, Q => 
                           n_1488, QN => n1529);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n10399, CK => CLK, Q => 
                           n_1489, QN => n1530);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n10400, CK => CLK, Q => 
                           n_1490, QN => n1531);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n10401, CK => CLK, Q => 
                           n_1491, QN => n1532);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n10402, CK => CLK, Q => 
                           n_1492, QN => n1533);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n10403, CK => CLK, Q => 
                           n_1493, QN => n1534);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n10404, CK => CLK, Q => 
                           n_1494, QN => n1535);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n10349, CK => CLK, Q => 
                           n8322, QN => n1536);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n10350, CK => CLK, Q => 
                           n_1495, QN => n1537);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n10351, CK => CLK, Q => 
                           n_1496, QN => n1538);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n10352, CK => CLK, Q => 
                           n_1497, QN => n1539);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n10353, CK => CLK, Q => 
                           n_1498, QN => n1540);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n10354, CK => CLK, Q => 
                           n_1499, QN => n1541);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n10355, CK => CLK, Q => 
                           n_1500, QN => n1542);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n10356, CK => CLK, Q => 
                           n_1501, QN => n1543);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n10357, CK => CLK, Q => 
                           n_1502, QN => n1544);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n10358, CK => CLK, Q => 
                           n_1503, QN => n1545);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n10359, CK => CLK, Q => 
                           n_1504, QN => n1546);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n10360, CK => CLK, Q => 
                           n_1505, QN => n1547);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n10361, CK => CLK, Q => 
                           n_1506, QN => n1548);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n10362, CK => CLK, Q => 
                           n_1507, QN => n1549);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n10363, CK => CLK, Q => 
                           n_1508, QN => n1550);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n10364, CK => CLK, Q => 
                           n_1509, QN => n1551);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n10365, CK => CLK, Q => 
                           n_1510, QN => n1552);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n10366, CK => CLK, Q => 
                           n_1511, QN => n1553);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n10367, CK => CLK, Q => 
                           n_1512, QN => n1554);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n10368, CK => CLK, Q => 
                           n_1513, QN => n1555);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n10369, CK => CLK, Q => 
                           n_1514, QN => n1556);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n10370, CK => CLK, Q => 
                           n_1515, QN => n1557);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n10371, CK => CLK, Q => 
                           n_1516, QN => n1558);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n10372, CK => CLK, Q => 
                           n_1517, QN => n1559);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n10317, CK => CLK, Q => 
                           n_1518, QN => n2351);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n10318, CK => CLK, Q => 
                           n_1519, QN => n2352);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n10319, CK => CLK, Q => 
                           n_1520, QN => n2353);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n10320, CK => CLK, Q => 
                           n_1521, QN => n2354);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n10321, CK => CLK, Q => 
                           n_1522, QN => n2355);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n10322, CK => CLK, Q => 
                           n_1523, QN => n2356);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n10323, CK => CLK, Q => 
                           n_1524, QN => n2357);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n10324, CK => CLK, Q => 
                           n_1525, QN => n2358);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n10325, CK => CLK, Q => 
                           n_1526, QN => n2359);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n10326, CK => CLK, Q => 
                           n_1527, QN => n2360);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n10327, CK => CLK, Q => 
                           n_1528, QN => n2361);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n10328, CK => CLK, Q => 
                           n_1529, QN => n2362);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n10329, CK => CLK, Q => 
                           n_1530, QN => n2363);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n10330, CK => CLK, Q => 
                           n_1531, QN => n2364);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n10332, CK => CLK, Q => 
                           n_1532, QN => n1560);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n10333, CK => CLK, Q => 
                           n_1533, QN => n1561);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n10334, CK => CLK, Q => 
                           n_1534, QN => n1562);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n10335, CK => CLK, Q => 
                           n_1535, QN => n1563);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n10336, CK => CLK, Q => 
                           n_1536, QN => n1564);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n10285, CK => CLK, Q => 
                           n_1537, QN => n2365);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n10286, CK => CLK, Q => 
                           n_1538, QN => n2366);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n10287, CK => CLK, Q => 
                           n_1539, QN => n2367);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n10288, CK => CLK, Q => 
                           n_1540, QN => n2368);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n10289, CK => CLK, Q => 
                           n_1541, QN => n2369);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n10290, CK => CLK, Q => 
                           n_1542, QN => n2370);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n10291, CK => CLK, Q => 
                           n_1543, QN => n2371);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n10292, CK => CLK, Q => 
                           n_1544, QN => n2372);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n10293, CK => CLK, Q => 
                           n_1545, QN => n2373);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n10294, CK => CLK, Q => 
                           n_1546, QN => n2374);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n10295, CK => CLK, Q => 
                           n_1547, QN => n2375);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n10296, CK => CLK, Q => 
                           n_1548, QN => n2376);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n10297, CK => CLK, Q => 
                           n_1549, QN => n2377);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n10298, CK => CLK, Q => 
                           n_1550, QN => n2378);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n10299, CK => CLK, Q => 
                           n_1551, QN => n1565);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n10300, CK => CLK, Q => 
                           n_1552, QN => n1566);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n10301, CK => CLK, Q => 
                           n_1553, QN => n1567);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n10302, CK => CLK, Q => 
                           n_1554, QN => n1568);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n10303, CK => CLK, Q => 
                           n_1555, QN => n1569);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n10304, CK => CLK, Q => 
                           n_1556, QN => n1570);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n10305, CK => CLK, Q => 
                           n_1557, QN => n1571);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n10306, CK => CLK, Q => 
                           n_1558, QN => n1572);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n10307, CK => CLK, Q => 
                           n_1559, QN => n1573);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n10308, CK => CLK, Q => 
                           n_1560, QN => n1574);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n10264, CK => CLK, Q => 
                           n770, QN => n2390);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n10221, CK => CLK, Q => 
                           n8290, QN => n1575);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n10222, CK => CLK, Q => 
                           n8291, QN => n1576);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n10223, CK => CLK, Q => 
                           n8292, QN => n1577);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n10224, CK => CLK, Q => 
                           n8293, QN => n1578);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n10225, CK => CLK, Q => 
                           n8294, QN => n1579);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n10226, CK => CLK, Q => 
                           n8295, QN => n1580);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n10227, CK => CLK, Q => 
                           n8296, QN => n1581);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n10228, CK => CLK, Q => 
                           n8297, QN => n1582);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n10229, CK => CLK, Q => 
                           n8298, QN => n1583);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n10230, CK => CLK, Q => 
                           n8299, QN => n1584);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n10231, CK => CLK, Q => 
                           n8300, QN => n1585);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n10232, CK => CLK, Q => 
                           n8301, QN => n1586);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n10233, CK => CLK, Q => 
                           n8302, QN => n1587);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n10234, CK => CLK, Q => 
                           n8303, QN => n1588);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n10235, CK => CLK, Q => 
                           n8304, QN => n1589);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n10236, CK => CLK, Q => 
                           n8305, QN => n1590);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n10237, CK => CLK, Q => 
                           n8306, QN => n1591);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n10238, CK => CLK, Q => 
                           n8307, QN => n1592);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n10239, CK => CLK, Q => 
                           n8308, QN => n1593);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n10240, CK => CLK, Q => 
                           n8309, QN => n1594);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n10241, CK => CLK, Q => 
                           n8310, QN => n1595);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n10242, CK => CLK, Q => 
                           n8311, QN => n1596);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n10243, CK => CLK, Q => 
                           n8312, QN => n1597);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n10244, CK => CLK, Q => 
                           n8313, QN => n1598);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n9648, CK => CLK, Q => 
                           n8103, QN => n415);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n9936, CK => CLK, Q => 
                           n8167, QN => n1708);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n9904, CK => CLK, Q => 
                           n8135, QN => n1709);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n9808, CK => CLK, Q => 
                           n7080, QN => n1710);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n9776, CK => CLK, Q => 
                           n_1561, QN => n1711);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n9688, CK => CLK, Q => n752
                           , QN => n2418);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n9689, CK => CLK, Q => n816
                           , QN => n2419);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n10040, CK => CLK, Q => 
                           n763, QN => n2497);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n10041, CK => CLK, Q => 
                           n827, QN => n2519);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n10044, CK => CLK, Q => n94
                           , QN => n1712);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n10045, CK => CLK, Q => n88
                           , QN => n1713);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n10046, CK => CLK, Q => n82
                           , QN => n1714);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n10047, CK => CLK, Q => n76
                           , QN => n1715);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n9933, CK => CLK, Q => 
                           n8164, QN => n1608);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n9937, CK => CLK, Q => 
                           n8168, QN => n1609);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n9938, CK => CLK, Q => 
                           n8169, QN => n1610);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n9939, CK => CLK, Q => 
                           n8170, QN => n1611);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n9940, CK => CLK, Q => 
                           n8171, QN => n1612);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n9941, CK => CLK, Q => 
                           n8172, QN => n1613);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n9942, CK => CLK, Q => 
                           n8173, QN => n1614);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n9943, CK => CLK, Q => 
                           n8174, QN => n1615);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n9944, CK => CLK, Q => 
                           n8175, QN => n1616);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n9946, CK => CLK, Q => 
                           n8177, QN => n1618);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n9947, CK => CLK, Q => 
                           n8178, QN => n1619);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n9948, CK => CLK, Q => 
                           n8179, QN => n1620);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n9949, CK => CLK, Q => 
                           n8180, QN => n1621);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n9950, CK => CLK, Q => 
                           n8181, QN => n1622);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n9951, CK => CLK, Q => 
                           n8182, QN => n1623);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n9952, CK => CLK, Q => 
                           n8183, QN => n1624);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n9953, CK => CLK, Q => 
                           n8184, QN => n1625);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n9954, CK => CLK, Q => 
                           n8185, QN => n1626);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n9955, CK => CLK, Q => n8186
                           , QN => n1627);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n9956, CK => CLK, Q => n8187
                           , QN => n1628);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n9901, CK => CLK, Q => 
                           n8132, QN => n1629);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n9905, CK => CLK, Q => 
                           n8136, QN => n1630);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n9906, CK => CLK, Q => 
                           n8137, QN => n1631);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n9907, CK => CLK, Q => 
                           n8138, QN => n1632);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n9908, CK => CLK, Q => 
                           n8139, QN => n1633);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n9909, CK => CLK, Q => 
                           n8140, QN => n1634);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n9910, CK => CLK, Q => 
                           n8141, QN => n1635);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n9911, CK => CLK, Q => 
                           n8142, QN => n1636);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n9912, CK => CLK, Q => 
                           n8143, QN => n1637);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n9914, CK => CLK, Q => 
                           n8145, QN => n1639);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n9915, CK => CLK, Q => 
                           n8146, QN => n1640);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n9916, CK => CLK, Q => 
                           n8147, QN => n1641);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n9917, CK => CLK, Q => 
                           n8148, QN => n1642);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n9918, CK => CLK, Q => 
                           n8149, QN => n1643);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n9919, CK => CLK, Q => 
                           n8150, QN => n1644);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n9920, CK => CLK, Q => 
                           n8151, QN => n1645);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n9921, CK => CLK, Q => 
                           n8152, QN => n1646);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n9922, CK => CLK, Q => 
                           n8153, QN => n1647);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n9923, CK => CLK, Q => n8154
                           , QN => n1648);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n9924, CK => CLK, Q => n8155
                           , QN => n1649);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n9881, CK => CLK, Q => n822
                           , QN => n2447);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n9849, CK => CLK, Q => n821
                           , QN => n2468);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n9805, CK => CLK, Q => 
                           n7104, QN => n1650);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n9809, CK => CLK, Q => 
                           n7071, QN => n1651);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n9810, CK => CLK, Q => 
                           n7063, QN => n1652);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n9811, CK => CLK, Q => 
                           n7056, QN => n1653);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n9812, CK => CLK, Q => 
                           n7047, QN => n1654);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n9813, CK => CLK, Q => 
                           n7039, QN => n1655);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n9814, CK => CLK, Q => 
                           n7032, QN => n1656);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n9815, CK => CLK, Q => 
                           n7018, QN => n1657);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n9818, CK => CLK, Q => 
                           n6979, QN => n1660);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n9819, CK => CLK, Q => 
                           n6965, QN => n1661);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n9820, CK => CLK, Q => 
                           n6952, QN => n1662);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n9821, CK => CLK, Q => 
                           n6940, QN => n1663);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n9822, CK => CLK, Q => 
                           n6925, QN => n1664);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n9823, CK => CLK, Q => 
                           n6915, QN => n1665);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n9824, CK => CLK, Q => 
                           n6898, QN => n1666);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n9825, CK => CLK, Q => 
                           n6889, QN => n1667);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n9826, CK => CLK, Q => 
                           n6871, QN => n1668);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n9827, CK => CLK, Q => n6859
                           , QN => n1669);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n9828, CK => CLK, Q => n6845
                           , QN => n1670);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n9773, CK => CLK, Q => 
                           n_1562, QN => n1671);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n9777, CK => CLK, Q => 
                           n_1563, QN => n1672);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n9778, CK => CLK, Q => 
                           n_1564, QN => n1673);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n9779, CK => CLK, Q => 
                           n_1565, QN => n1674);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n9780, CK => CLK, Q => 
                           n_1566, QN => n1675);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n9781, CK => CLK, Q => 
                           n_1567, QN => n1676);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n9782, CK => CLK, Q => 
                           n_1568, QN => n1677);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n9783, CK => CLK, Q => 
                           n_1569, QN => n1678);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n9784, CK => CLK, Q => 
                           n_1570, QN => n1679);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n9785, CK => CLK, Q => 
                           n_1571, QN => n1680);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n9786, CK => CLK, Q => 
                           n_1572, QN => n1681);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n9787, CK => CLK, Q => 
                           n_1573, QN => n1682);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n9788, CK => CLK, Q => 
                           n_1574, QN => n1683);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n9789, CK => CLK, Q => 
                           n_1575, QN => n1684);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n9790, CK => CLK, Q => 
                           n_1576, QN => n1685);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n9791, CK => CLK, Q => 
                           n_1577, QN => n1686);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n9792, CK => CLK, Q => 
                           n_1578, QN => n1687);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n9793, CK => CLK, Q => 
                           n_1579, QN => n1688);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n9794, CK => CLK, Q => 
                           n_1580, QN => n1689);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n9795, CK => CLK, Q => 
                           n_1581, QN => n1690);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n9796, CK => CLK, Q => 
                           n_1582, QN => n1691);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n9752, CK => CLK, Q => 
                           n_1583, QN => n2480);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n9753, CK => CLK, Q => 
                           n_1584, QN => n2481);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n9756, CK => CLK, Q => 
                           n_1585, QN => n1692);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n9757, CK => CLK, Q => 
                           n_1586, QN => n1693);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n9758, CK => CLK, Q => 
                           n_1587, QN => n1694);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n9759, CK => CLK, Q => 
                           n_1588, QN => n1695);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n9760, CK => CLK, Q => 
                           n_1589, QN => n1696);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n9720, CK => CLK, Q => 
                           n_1590, QN => n2482);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n9721, CK => CLK, Q => 
                           n_1591, QN => n2483);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n9723, CK => CLK, Q => 
                           n_1592, QN => n1697);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n9724, CK => CLK, Q => 
                           n_1593, QN => n1698);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n9725, CK => CLK, Q => 
                           n_1594, QN => n1699);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n9726, CK => CLK, Q => 
                           n_1595, QN => n1700);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n9727, CK => CLK, Q => 
                           n_1596, QN => n1701);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n9728, CK => CLK, Q => 
                           n_1597, QN => n1702);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n9729, CK => CLK, Q => 
                           n_1598, QN => n1703);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n9730, CK => CLK, Q => 
                           n_1599, QN => n1704);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n9731, CK => CLK, Q => 
                           n_1600, QN => n1705);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n9732, CK => CLK, Q => 
                           n_1601, QN => n1706);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n10062, CK => CLK, Q => 
                           n_1602, QN => n1085);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n10063, CK => CLK, Q => 
                           n_1603, QN => n1086);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n9934, CK => CLK, Q => 
                           n8165, QN => n1599);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n9935, CK => CLK, Q => 
                           n8166, QN => n1600);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n9902, CK => CLK, Q => 
                           n8133, QN => n1601);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n9903, CK => CLK, Q => 
                           n8134, QN => n1602);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n9806, CK => CLK, Q => 
                           n7095, QN => n1603);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n9807, CK => CLK, Q => 
                           n7087, QN => n1604);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n9774, CK => CLK, Q => 
                           n_1604, QN => n1605);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n9775, CK => CLK, Q => 
                           n_1605, QN => n1606);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n10008, CK => CLK, Q => 
                           n762, QN => n2431);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n10009, CK => CLK, Q => 
                           n826, QN => n2432);
   REGISTERS_reg_71_21_inst : DFF_X1 port map( D => n11479, CK => CLK, Q => 
                           n736, QN => n2505);
   REGISTERS_reg_71_20_inst : DFF_X1 port map( D => n11480, CK => CLK, Q => 
                           n800, QN => n2506);
   REGISTERS_reg_70_0_inst : DFF_X1 port map( D => n11468, CK => CLK, Q => 
                           n1716, QN => n6727);
   REGISTERS_reg_69_7_inst : DFF_X1 port map( D => n11429, CK => CLK, Q => 
                           n1717, QN => n6896);
   REGISTERS_reg_69_6_inst : DFF_X1 port map( D => n11430, CK => CLK, Q => 
                           n1718, QN => n6872);
   REGISTERS_reg_69_5_inst : DFF_X1 port map( D => n11431, CK => CLK, Q => 
                           n1719, QN => n6848);
   REGISTERS_reg_69_4_inst : DFF_X1 port map( D => n11432, CK => CLK, Q => 
                           n1720, QN => n6824);
   REGISTERS_reg_69_3_inst : DFF_X1 port map( D => n11433, CK => CLK, Q => 
                           n1721, QN => n6800);
   REGISTERS_reg_69_2_inst : DFF_X1 port map( D => n11434, CK => CLK, Q => 
                           n1722, QN => n6776);
   REGISTERS_reg_69_1_inst : DFF_X1 port map( D => n11435, CK => CLK, Q => 
                           n1723, QN => n6752);
   REGISTERS_reg_69_0_inst : DFF_X1 port map( D => n11436, CK => CLK, Q => 
                           n1724, QN => n6728);
   REGISTERS_reg_60_7_inst : DFF_X1 port map( D => n11141, CK => CLK, Q => 
                           n1733, QN => n6899);
   REGISTERS_reg_60_6_inst : DFF_X1 port map( D => n11142, CK => CLK, Q => 
                           n1734, QN => n6875);
   REGISTERS_reg_60_5_inst : DFF_X1 port map( D => n11143, CK => CLK, Q => 
                           n1735, QN => n6851);
   REGISTERS_reg_60_4_inst : DFF_X1 port map( D => n11144, CK => CLK, Q => 
                           n1736, QN => n6827);
   REGISTERS_reg_60_3_inst : DFF_X1 port map( D => n11145, CK => CLK, Q => 
                           n1737, QN => n6803);
   REGISTERS_reg_60_2_inst : DFF_X1 port map( D => n11146, CK => CLK, Q => 
                           n1738, QN => n6779);
   REGISTERS_reg_60_1_inst : DFF_X1 port map( D => n11147, CK => CLK, Q => 
                           n1739, QN => n6755);
   REGISTERS_reg_60_0_inst : DFF_X1 port map( D => n11148, CK => CLK, Q => 
                           n1740, QN => n6731);
   REGISTERS_reg_53_7_inst : DFF_X1 port map( D => n10917, CK => CLK, Q => 
                           n_1606, QN => n6900);
   REGISTERS_reg_53_6_inst : DFF_X1 port map( D => n10918, CK => CLK, Q => 
                           n_1607, QN => n6876);
   REGISTERS_reg_53_5_inst : DFF_X1 port map( D => n10919, CK => CLK, Q => 
                           n_1608, QN => n6852);
   REGISTERS_reg_53_4_inst : DFF_X1 port map( D => n10920, CK => CLK, Q => 
                           n_1609, QN => n6828);
   REGISTERS_reg_53_3_inst : DFF_X1 port map( D => n10921, CK => CLK, Q => 
                           n_1610, QN => n6804);
   REGISTERS_reg_53_1_inst : DFF_X1 port map( D => n10923, CK => CLK, Q => 
                           n_1611, QN => n6756);
   REGISTERS_reg_51_7_inst : DFF_X1 port map( D => n10853, CK => CLK, Q => 
                           n1743, QN => n6902);
   REGISTERS_reg_51_6_inst : DFF_X1 port map( D => n10854, CK => CLK, Q => 
                           n1744, QN => n6878);
   REGISTERS_reg_51_5_inst : DFF_X1 port map( D => n10855, CK => CLK, Q => 
                           n1745, QN => n6854);
   REGISTERS_reg_51_4_inst : DFF_X1 port map( D => n10856, CK => CLK, Q => 
                           n1746, QN => n6830);
   REGISTERS_reg_51_3_inst : DFF_X1 port map( D => n10857, CK => CLK, Q => 
                           n1747, QN => n6806);
   REGISTERS_reg_51_2_inst : DFF_X1 port map( D => n10858, CK => CLK, Q => 
                           n1748, QN => n6782);
   REGISTERS_reg_51_1_inst : DFF_X1 port map( D => n10859, CK => CLK, Q => 
                           n1749, QN => n6758);
   REGISTERS_reg_51_0_inst : DFF_X1 port map( D => n10860, CK => CLK, Q => 
                           n1750, QN => n6734);
   REGISTERS_reg_42_7_inst : DFF_X1 port map( D => n10565, CK => CLK, Q => 
                           n1759, QN => n6905);
   REGISTERS_reg_42_6_inst : DFF_X1 port map( D => n10566, CK => CLK, Q => 
                           n1760, QN => n6881);
   REGISTERS_reg_42_5_inst : DFF_X1 port map( D => n10567, CK => CLK, Q => 
                           n1761, QN => n6857);
   REGISTERS_reg_42_4_inst : DFF_X1 port map( D => n10568, CK => CLK, Q => 
                           n1762, QN => n6833);
   REGISTERS_reg_42_3_inst : DFF_X1 port map( D => n10569, CK => CLK, Q => 
                           n1763, QN => n6809);
   REGISTERS_reg_42_2_inst : DFF_X1 port map( D => n10570, CK => CLK, Q => 
                           n1764, QN => n6785);
   REGISTERS_reg_42_1_inst : DFF_X1 port map( D => n10571, CK => CLK, Q => 
                           n1765, QN => n6761);
   REGISTERS_reg_42_0_inst : DFF_X1 port map( D => n10572, CK => CLK, Q => 
                           n1766, QN => n6737);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n10469, CK => CLK, Q => 
                           n1767, QN => n7785);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n10470, CK => CLK, Q => 
                           n1768, QN => n7789);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n10471, CK => CLK, Q => 
                           n1769, QN => n7793);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n10472, CK => CLK, Q => 
                           n1770, QN => n7797);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n10473, CK => CLK, Q => 
                           n1771, QN => n7801);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n10474, CK => CLK, Q => 
                           n1772, QN => n7805);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n10475, CK => CLK, Q => 
                           n1773, QN => n7809);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n10437, CK => CLK, Q => 
                           n1774, QN => n7784);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n10438, CK => CLK, Q => 
                           n1775, QN => n7788);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n10439, CK => CLK, Q => 
                           n1776, QN => n7792);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n10440, CK => CLK, Q => 
                           n1777, QN => n7796);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n10441, CK => CLK, Q => 
                           n1778, QN => n7800);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n10442, CK => CLK, Q => 
                           n1779, QN => n7804);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n10443, CK => CLK, Q => 
                           n1780, QN => n7808);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n10444, CK => CLK, Q => 
                           n1781, QN => n7812);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n10341, CK => CLK, Q => 
                           n_1612, QN => n6906);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n10342, CK => CLK, Q => 
                           n_1613, QN => n6882);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n10343, CK => CLK, Q => 
                           n_1614, QN => n6858);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n10344, CK => CLK, Q => 
                           n_1615, QN => n6834);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n10345, CK => CLK, Q => 
                           n_1616, QN => n6810);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n10346, CK => CLK, Q => 
                           n_1617, QN => n6786);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n10347, CK => CLK, Q => 
                           n_1618, QN => n6762);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n10277, CK => CLK, Q => 
                           n1784, QN => n6908);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n10278, CK => CLK, Q => 
                           n1785, QN => n6884);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n10279, CK => CLK, Q => 
                           n1786, QN => n6860);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n10280, CK => CLK, Q => 
                           n1787, QN => n6836);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n10281, CK => CLK, Q => 
                           n1788, QN => n6812);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n10282, CK => CLK, Q => 
                           n1789, QN => n6788);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n10283, CK => CLK, Q => 
                           n1790, QN => n6764);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n10284, CK => CLK, Q => 
                           n1791, QN => n6740);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n10181, CK => CLK, Q => 
                           n1792, QN => n7887);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n10182, CK => CLK, Q => 
                           n1793, QN => n7890);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n10183, CK => CLK, Q => 
                           n1794, QN => n7893);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n10184, CK => CLK, Q => 
                           n1795, QN => n7896);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n10185, CK => CLK, Q => 
                           n1796, QN => n7899);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n10186, CK => CLK, Q => 
                           n1797, QN => n7902);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n10187, CK => CLK, Q => 
                           n1798, QN => n7905);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n10149, CK => CLK, Q => 
                           n1799, QN => n7886);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n10150, CK => CLK, Q => 
                           n1800, QN => n7889);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n10151, CK => CLK, Q => 
                           n1801, QN => n7892);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n10152, CK => CLK, Q => 
                           n1802, QN => n7895);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n10153, CK => CLK, Q => 
                           n1803, QN => n7898);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n10154, CK => CLK, Q => 
                           n1804, QN => n7901);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n10155, CK => CLK, Q => 
                           n1805, QN => n7904);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n10156, CK => CLK, Q => 
                           n1806, QN => n8898);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n10032, CK => CLK, Q => 
                           n_1619, QN => n7413);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n9989, CK => CLK, Q => n1807
                           , QN => n6911);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n9990, CK => CLK, Q => n1808
                           , QN => n6887);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n9991, CK => CLK, Q => n1809
                           , QN => n6863);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n9992, CK => CLK, Q => n1810
                           , QN => n6839);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n9993, CK => CLK, Q => n1811
                           , QN => n6815);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n9994, CK => CLK, Q => n1812
                           , QN => n6791);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n9995, CK => CLK, Q => n1813
                           , QN => n6767);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n9996, CK => CLK, Q => n1814
                           , QN => n6743);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n9573, CK => CLK, Q => n1815
                           , QN => n7640);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n9574, CK => CLK, Q => n1816
                           , QN => n7646);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n9575, CK => CLK, Q => n1817
                           , QN => n7652);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n9576, CK => CLK, Q => n1818
                           , QN => n7658);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n9577, CK => CLK, Q => n1819
                           , QN => n7664);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n9578, CK => CLK, Q => n1820
                           , QN => n7670);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n9579, CK => CLK, Q => n1821
                           , QN => n7676);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n9580, CK => CLK, Q => n1822
                           , QN => n7682);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n9285, CK => CLK, Q => n1823,
                           QN => n7642);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n9286, CK => CLK, Q => n1824,
                           QN => n7648);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n9287, CK => CLK, Q => n1825,
                           QN => n7654);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n9288, CK => CLK, Q => n1826,
                           QN => n7660);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n9289, CK => CLK, Q => n1827,
                           QN => n7666);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n9290, CK => CLK, Q => n1828,
                           QN => n7672);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n9291, CK => CLK, Q => n1829,
                           QN => n7678);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n9292, CK => CLK, Q => n1830,
                           QN => n7684);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n10000, CK => CLK, Q => 
                           n_1620, QN => n7414);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n10033, CK => CLK, Q => 
                           n_1621, QN => n7389);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n10034, CK => CLK, Q => 
                           n_1622, QN => n7365);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n10035, CK => CLK, Q => 
                           n_1623, QN => n7341);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n10036, CK => CLK, Q => 
                           n_1624, QN => n7317);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n10037, CK => CLK, Q => 
                           n_1625, QN => n7293);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n10038, CK => CLK, Q => 
                           n_1626, QN => n7269);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n10039, CK => CLK, Q => 
                           n_1627, QN => n7245);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n9893, CK => CLK, Q => n1831
                           , QN => n7787);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n9894, CK => CLK, Q => n1832
                           , QN => n7791);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n9895, CK => CLK, Q => n1833
                           , QN => n7795);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n9896, CK => CLK, Q => n1834
                           , QN => n7799);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n9897, CK => CLK, Q => n1835
                           , QN => n7803);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n9898, CK => CLK, Q => n1836
                           , QN => n7807);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n9899, CK => CLK, Q => n1837
                           , QN => n7811);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n9900, CK => CLK, Q => n1838
                           , QN => n7815);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n9861, CK => CLK, Q => n1839
                           , QN => n7786);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n9862, CK => CLK, Q => n1840
                           , QN => n7790);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n9863, CK => CLK, Q => n1841
                           , QN => n7794);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n9864, CK => CLK, Q => n1842
                           , QN => n7798);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n9865, CK => CLK, Q => n1843
                           , QN => n7802);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n9866, CK => CLK, Q => n1844
                           , QN => n7806);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n9867, CK => CLK, Q => n1845
                           , QN => n7810);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n9868, CK => CLK, Q => n1846
                           , QN => n7814);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n9765, CK => CLK, Q => 
                           n_1628, QN => n6912);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n9766, CK => CLK, Q => 
                           n_1629, QN => n6888);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n9767, CK => CLK, Q => 
                           n_1630, QN => n6864);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n9768, CK => CLK, Q => 
                           n_1631, QN => n6840);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n9769, CK => CLK, Q => 
                           n_1632, QN => n6816);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n9770, CK => CLK, Q => 
                           n_1633, QN => n6792);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n9771, CK => CLK, Q => 
                           n_1634, QN => n6768);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n9772, CK => CLK, Q => 
                           n_1635, QN => n6744);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n9740, CK => CLK, Q => 
                           n_1636, QN => n6745);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n9701, CK => CLK, Q => n1847
                           , QN => n6914);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n9702, CK => CLK, Q => n1848
                           , QN => n6890);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n9703, CK => CLK, Q => n1849
                           , QN => n6866);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n9704, CK => CLK, Q => n1850
                           , QN => n6842);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n9705, CK => CLK, Q => n1851
                           , QN => n6818);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n9706, CK => CLK, Q => n1852
                           , QN => n6794);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n9707, CK => CLK, Q => n1853
                           , QN => n6770);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n9708, CK => CLK, Q => n1854
                           , QN => n6746);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n9677, CK => CLK, Q => 
                           n1855, QN => n7490);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n9678, CK => CLK, Q => 
                           n2403, QN => n7466);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n9679, CK => CLK, Q => 
                           n2404, QN => n7442);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n9657, CK => CLK, Q => n424
                           , QN => n815);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n9625, CK => CLK, Q => n448
                           , QN => n814);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n9549, CK => CLK, Q => 
                           n1856, QN => n7496);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n9550, CK => CLK, Q => 
                           n1857, QN => n7502);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n9551, CK => CLK, Q => 
                           n1858, QN => n7508);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n9552, CK => CLK, Q => 
                           n1859, QN => n7514);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n9553, CK => CLK, Q => 
                           n1860, QN => n7520);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n9554, CK => CLK, Q => 
                           n1861, QN => n7526);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n9555, CK => CLK, Q => 
                           n1862, QN => n7532);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n9556, CK => CLK, Q => 
                           n1863, QN => n7538);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n9557, CK => CLK, Q => 
                           n1864, QN => n7544);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n9558, CK => CLK, Q => 
                           n1865, QN => n7550);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n9559, CK => CLK, Q => 
                           n1866, QN => n7556);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n9560, CK => CLK, Q => 
                           n1867, QN => n7562);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n9562, CK => CLK, Q => 
                           n1869, QN => n7574);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n9563, CK => CLK, Q => 
                           n1870, QN => n7580);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n9564, CK => CLK, Q => 
                           n1871, QN => n7586);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n9565, CK => CLK, Q => 
                           n1872, QN => n7592);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n9566, CK => CLK, Q => 
                           n1873, QN => n7598);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n9567, CK => CLK, Q => 
                           n1874, QN => n7604);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n9568, CK => CLK, Q => 
                           n1875, QN => n7610);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n9569, CK => CLK, Q => 
                           n1876, QN => n7616);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n9570, CK => CLK, Q => 
                           n1877, QN => n7622);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n9571, CK => CLK, Q => n1878
                           , QN => n7628);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n9572, CK => CLK, Q => n1879
                           , QN => n7634);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n9529, CK => CLK, Q => n496
                           , QN => n811);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n9400, CK => CLK, Q => n1000
                           , QN => n743);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n9401, CK => CLK, Q => n1001
                           , QN => n807);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n9369, CK => CLK, Q => n1025
                           , QN => n806);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n9337, CK => CLK, Q => n544,
                           QN => n805);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n9261, CK => CLK, Q => n1880
                           , QN => n7498);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n9262, CK => CLK, Q => n1881
                           , QN => n7504);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n9263, CK => CLK, Q => n1882
                           , QN => n7510);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n9264, CK => CLK, Q => n1883
                           , QN => n7516);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n9265, CK => CLK, Q => n1884
                           , QN => n7522);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n9266, CK => CLK, Q => n1885
                           , QN => n7528);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n9267, CK => CLK, Q => n1886
                           , QN => n7534);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n9268, CK => CLK, Q => n1887
                           , QN => n7540);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n9269, CK => CLK, Q => n1888
                           , QN => n7546);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n9270, CK => CLK, Q => n1889
                           , QN => n7552);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n9271, CK => CLK, Q => n1890
                           , QN => n7558);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n9272, CK => CLK, Q => n1891
                           , QN => n7564);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n9274, CK => CLK, Q => n1893
                           , QN => n7576);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n9275, CK => CLK, Q => n1894
                           , QN => n7582);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n9276, CK => CLK, Q => n1895
                           , QN => n7588);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n9277, CK => CLK, Q => n1896
                           , QN => n7594);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n9278, CK => CLK, Q => n1897
                           , QN => n7600);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n9279, CK => CLK, Q => n1898
                           , QN => n7606);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n9280, CK => CLK, Q => n1899
                           , QN => n7612);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n9281, CK => CLK, Q => n1900
                           , QN => n7618);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n9282, CK => CLK, Q => n1901
                           , QN => n7624);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n9283, CK => CLK, Q => n1902,
                           QN => n7630);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n9284, CK => CLK, Q => n1903,
                           QN => n7636);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n9241, CK => CLK, Q => n592,
                           QN => n802);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n9191, CK => CLK, Q => n616,
                           QN => n801);
   REGISTERS_reg_70_31_inst : DFF_X1 port map( D => n11437, CK => CLK, Q => 
                           n1904, QN => n7471);
   REGISTERS_reg_70_30_inst : DFF_X1 port map( D => n11438, CK => CLK, Q => 
                           n1905, QN => n7447);
   REGISTERS_reg_70_29_inst : DFF_X1 port map( D => n11439, CK => CLK, Q => 
                           n1906, QN => n7423);
   REGISTERS_reg_70_28_inst : DFF_X1 port map( D => n11440, CK => CLK, Q => 
                           n1907, QN => n7399);
   REGISTERS_reg_70_27_inst : DFF_X1 port map( D => n11441, CK => CLK, Q => 
                           n1908, QN => n7375);
   REGISTERS_reg_70_26_inst : DFF_X1 port map( D => n11442, CK => CLK, Q => 
                           n1909, QN => n7351);
   REGISTERS_reg_70_25_inst : DFF_X1 port map( D => n11443, CK => CLK, Q => 
                           n1910, QN => n7327);
   REGISTERS_reg_70_24_inst : DFF_X1 port map( D => n11444, CK => CLK, Q => 
                           n1911, QN => n7303);
   REGISTERS_reg_70_23_inst : DFF_X1 port map( D => n11445, CK => CLK, Q => 
                           n1912, QN => n7279);
   REGISTERS_reg_70_22_inst : DFF_X1 port map( D => n11446, CK => CLK, Q => 
                           n1913, QN => n7255);
   REGISTERS_reg_70_19_inst : DFF_X1 port map( D => n11449, CK => CLK, Q => 
                           n1916, QN => n7183);
   REGISTERS_reg_70_18_inst : DFF_X1 port map( D => n11450, CK => CLK, Q => 
                           n1917, QN => n7159);
   REGISTERS_reg_69_31_inst : DFF_X1 port map( D => n11405, CK => CLK, Q => 
                           n1918, QN => n7472);
   REGISTERS_reg_69_30_inst : DFF_X1 port map( D => n11406, CK => CLK, Q => 
                           n1919, QN => n7448);
   REGISTERS_reg_69_29_inst : DFF_X1 port map( D => n11407, CK => CLK, Q => 
                           n1920, QN => n7424);
   REGISTERS_reg_69_28_inst : DFF_X1 port map( D => n11408, CK => CLK, Q => 
                           n1921, QN => n7400);
   REGISTERS_reg_69_27_inst : DFF_X1 port map( D => n11409, CK => CLK, Q => 
                           n1922, QN => n7376);
   REGISTERS_reg_69_26_inst : DFF_X1 port map( D => n11410, CK => CLK, Q => 
                           n1923, QN => n7352);
   REGISTERS_reg_69_25_inst : DFF_X1 port map( D => n11411, CK => CLK, Q => 
                           n1924, QN => n7328);
   REGISTERS_reg_69_24_inst : DFF_X1 port map( D => n11412, CK => CLK, Q => 
                           n1925, QN => n7304);
   REGISTERS_reg_69_23_inst : DFF_X1 port map( D => n11413, CK => CLK, Q => 
                           n1926, QN => n7280);
   REGISTERS_reg_69_22_inst : DFF_X1 port map( D => n11414, CK => CLK, Q => 
                           n1927, QN => n7256);
   REGISTERS_reg_69_19_inst : DFF_X1 port map( D => n11417, CK => CLK, Q => 
                           n1930, QN => n7184);
   REGISTERS_reg_69_18_inst : DFF_X1 port map( D => n11418, CK => CLK, Q => 
                           n1931, QN => n7160);
   REGISTERS_reg_69_17_inst : DFF_X1 port map( D => n11419, CK => CLK, Q => 
                           n1932, QN => n7136);
   REGISTERS_reg_69_16_inst : DFF_X1 port map( D => n11420, CK => CLK, Q => 
                           n1933, QN => n7112);
   REGISTERS_reg_69_15_inst : DFF_X1 port map( D => n11421, CK => CLK, Q => 
                           n1934, QN => n7088);
   REGISTERS_reg_69_14_inst : DFF_X1 port map( D => n11422, CK => CLK, Q => 
                           n1935, QN => n7064);
   REGISTERS_reg_69_13_inst : DFF_X1 port map( D => n11423, CK => CLK, Q => 
                           n1936, QN => n7040);
   REGISTERS_reg_69_12_inst : DFF_X1 port map( D => n11424, CK => CLK, Q => 
                           n1937, QN => n7016);
   REGISTERS_reg_69_11_inst : DFF_X1 port map( D => n11425, CK => CLK, Q => 
                           n1938, QN => n6992);
   REGISTERS_reg_69_10_inst : DFF_X1 port map( D => n11426, CK => CLK, Q => 
                           n1939, QN => n6968);
   REGISTERS_reg_69_9_inst : DFF_X1 port map( D => n11427, CK => CLK, Q => 
                           n1940, QN => n6944);
   REGISTERS_reg_69_8_inst : DFF_X1 port map( D => n11428, CK => CLK, Q => 
                           n1941, QN => n6920);
   REGISTERS_reg_66_21_inst : DFF_X1 port map( D => n11319, CK => CLK, Q => 
                           n696, QN => n731);
   REGISTERS_reg_66_20_inst : DFF_X1 port map( D => n11320, CK => CLK, Q => 
                           n697, QN => n795);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n9497, CK => CLK, Q => n788,
                           QN => n810);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n10158, CK => CLK, Q => 
                           n1942, QN => n7818);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n10159, CK => CLK, Q => 
                           n1943, QN => n7821);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n10160, CK => CLK, Q => 
                           n1944, QN => n7824);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n10161, CK => CLK, Q => 
                           n1945, QN => n7827);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n10162, CK => CLK, Q => 
                           n1946, QN => n7830);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n10163, CK => CLK, Q => 
                           n1947, QN => n7833);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n10164, CK => CLK, Q => 
                           n1948, QN => n7836);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n10165, CK => CLK, Q => 
                           n1949, QN => n7839);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n10166, CK => CLK, Q => 
                           n1950, QN => n7842);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n10167, CK => CLK, Q => 
                           n1951, QN => n7845);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n10168, CK => CLK, Q => 
                           n1952, QN => n7848);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n10169, CK => CLK, Q => 
                           n1953, QN => n7851);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n10170, CK => CLK, Q => 
                           n1954, QN => n7854);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n10171, CK => CLK, Q => 
                           n1955, QN => n7857);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n10172, CK => CLK, Q => 
                           n1956, QN => n7860);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n10173, CK => CLK, Q => 
                           n1957, QN => n7863);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n10174, CK => CLK, Q => 
                           n1958, QN => n7866);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n10175, CK => CLK, Q => 
                           n1959, QN => n7869);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n10176, CK => CLK, Q => 
                           n1960, QN => n7872);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n10177, CK => CLK, Q => 
                           n1961, QN => n7875);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n10178, CK => CLK, Q => 
                           n1962, QN => n7878);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n10179, CK => CLK, Q => 
                           n1963, QN => n7881);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n10180, CK => CLK, Q => 
                           n1964, QN => n7884);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n10125, CK => CLK, Q => 
                           n1965, QN => n7686);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n10126, CK => CLK, Q => 
                           n1966, QN => n7817);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n10127, CK => CLK, Q => 
                           n1967, QN => n7820);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n10128, CK => CLK, Q => 
                           n1968, QN => n7823);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n10129, CK => CLK, Q => 
                           n1969, QN => n7826);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n10130, CK => CLK, Q => 
                           n1970, QN => n7829);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n10131, CK => CLK, Q => 
                           n1971, QN => n7832);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n10132, CK => CLK, Q => 
                           n1972, QN => n7835);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n10133, CK => CLK, Q => 
                           n1973, QN => n7838);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n10134, CK => CLK, Q => 
                           n1974, QN => n7841);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n10135, CK => CLK, Q => 
                           n1975, QN => n7844);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n10136, CK => CLK, Q => 
                           n1976, QN => n7847);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n10137, CK => CLK, Q => 
                           n1977, QN => n7850);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n10138, CK => CLK, Q => 
                           n1978, QN => n7853);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n10139, CK => CLK, Q => 
                           n1979, QN => n7856);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n10140, CK => CLK, Q => 
                           n1980, QN => n7859);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n10141, CK => CLK, Q => 
                           n1981, QN => n7862);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n10142, CK => CLK, Q => 
                           n1982, QN => n7865);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n10143, CK => CLK, Q => 
                           n1983, QN => n7868);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n10144, CK => CLK, Q => 
                           n1984, QN => n7871);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n10145, CK => CLK, Q => 
                           n1985, QN => n7874);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n10146, CK => CLK, Q => 
                           n1986, QN => n7877);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n10147, CK => CLK, Q => 
                           n1987, QN => n7880);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n10148, CK => CLK, Q => 
                           n1988, QN => n7883);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n10105, CK => CLK, Q => 
                           n_1637, QN => n829);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n10073, CK => CLK, Q => 
                           n_1638, QN => n828);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n9968, CK => CLK, Q => 
                           n1989, QN => n7415);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n9969, CK => CLK, Q => 
                           n1990, QN => n7391);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n9970, CK => CLK, Q => 
                           n1991, QN => n7367);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n9971, CK => CLK, Q => 
                           n1992, QN => n7343);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n9972, CK => CLK, Q => 
                           n1993, QN => n7319);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n9973, CK => CLK, Q => 
                           n1994, QN => n7295);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n9974, CK => CLK, Q => 
                           n1995, QN => n7271);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n9975, CK => CLK, Q => 
                           n1996, QN => n7247);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n9978, CK => CLK, Q => 
                           n1999, QN => n7175);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n9979, CK => CLK, Q => 
                           n2000, QN => n7151);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n9980, CK => CLK, Q => 
                           n2001, QN => n7127);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n9981, CK => CLK, Q => 
                           n2002, QN => n7103);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n9982, CK => CLK, Q => 
                           n2003, QN => n7079);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n9983, CK => CLK, Q => 
                           n2004, QN => n7055);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n9984, CK => CLK, Q => 
                           n2005, QN => n7031);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n9985, CK => CLK, Q => 
                           n2006, QN => n7007);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n9986, CK => CLK, Q => 
                           n2007, QN => n6983);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n9987, CK => CLK, Q => n2008
                           , QN => n6959);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n9988, CK => CLK, Q => n2009
                           , QN => n6935);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n9742, CK => CLK, Q => 
                           n_1639, QN => n7464);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n9743, CK => CLK, Q => 
                           n_1640, QN => n7440);
   REGISTERS_reg_60_31_inst : DFF_X1 port map( D => n11117, CK => CLK, Q => 
                           n2043, QN => n7475);
   REGISTERS_reg_60_30_inst : DFF_X1 port map( D => n11118, CK => CLK, Q => 
                           n2044, QN => n7451);
   REGISTERS_reg_60_29_inst : DFF_X1 port map( D => n11119, CK => CLK, Q => 
                           n2045, QN => n7427);
   REGISTERS_reg_60_28_inst : DFF_X1 port map( D => n11120, CK => CLK, Q => 
                           n2046, QN => n7403);
   REGISTERS_reg_60_27_inst : DFF_X1 port map( D => n11121, CK => CLK, Q => 
                           n2047, QN => n7379);
   REGISTERS_reg_60_26_inst : DFF_X1 port map( D => n11122, CK => CLK, Q => 
                           n2048, QN => n7355);
   REGISTERS_reg_60_25_inst : DFF_X1 port map( D => n11123, CK => CLK, Q => 
                           n2049, QN => n7331);
   REGISTERS_reg_60_24_inst : DFF_X1 port map( D => n11124, CK => CLK, Q => 
                           n2050, QN => n7307);
   REGISTERS_reg_60_23_inst : DFF_X1 port map( D => n11125, CK => CLK, Q => 
                           n2051, QN => n7283);
   REGISTERS_reg_60_22_inst : DFF_X1 port map( D => n11126, CK => CLK, Q => 
                           n2052, QN => n7259);
   REGISTERS_reg_60_19_inst : DFF_X1 port map( D => n11129, CK => CLK, Q => 
                           n2055, QN => n7187);
   REGISTERS_reg_60_18_inst : DFF_X1 port map( D => n11130, CK => CLK, Q => 
                           n2056, QN => n7163);
   REGISTERS_reg_60_17_inst : DFF_X1 port map( D => n11131, CK => CLK, Q => 
                           n2057, QN => n7139);
   REGISTERS_reg_60_16_inst : DFF_X1 port map( D => n11132, CK => CLK, Q => 
                           n2058, QN => n7115);
   REGISTERS_reg_60_15_inst : DFF_X1 port map( D => n11133, CK => CLK, Q => 
                           n2059, QN => n7091);
   REGISTERS_reg_60_14_inst : DFF_X1 port map( D => n11134, CK => CLK, Q => 
                           n2060, QN => n7067);
   REGISTERS_reg_60_13_inst : DFF_X1 port map( D => n11135, CK => CLK, Q => 
                           n2061, QN => n7043);
   REGISTERS_reg_60_12_inst : DFF_X1 port map( D => n11136, CK => CLK, Q => 
                           n2062, QN => n7019);
   REGISTERS_reg_60_11_inst : DFF_X1 port map( D => n11137, CK => CLK, Q => 
                           n2063, QN => n6995);
   REGISTERS_reg_60_10_inst : DFF_X1 port map( D => n11138, CK => CLK, Q => 
                           n2064, QN => n6971);
   REGISTERS_reg_60_9_inst : DFF_X1 port map( D => n11139, CK => CLK, Q => 
                           n2065, QN => n6947);
   REGISTERS_reg_60_8_inst : DFF_X1 port map( D => n11140, CK => CLK, Q => 
                           n2066, QN => n6923);
   REGISTERS_reg_55_20_inst : DFF_X1 port map( D => n10968, CK => CLK, Q => 
                           n1252, QN => n786);
   REGISTERS_reg_53_12_inst : DFF_X1 port map( D => n10912, CK => CLK, Q => 
                           n_1641, QN => n7020);
   REGISTERS_reg_53_11_inst : DFF_X1 port map( D => n10913, CK => CLK, Q => 
                           n_1642, QN => n6996);
   REGISTERS_reg_53_10_inst : DFF_X1 port map( D => n10914, CK => CLK, Q => 
                           n_1643, QN => n6972);
   REGISTERS_reg_53_9_inst : DFF_X1 port map( D => n10915, CK => CLK, Q => 
                           n_1644, QN => n6948);
   REGISTERS_reg_53_8_inst : DFF_X1 port map( D => n10916, CK => CLK, Q => 
                           n_1645, QN => n6924);
   REGISTERS_reg_51_31_inst : DFF_X1 port map( D => n10829, CK => CLK, Q => 
                           n2095, QN => n7478);
   REGISTERS_reg_51_30_inst : DFF_X1 port map( D => n10830, CK => CLK, Q => 
                           n2096, QN => n7454);
   REGISTERS_reg_51_29_inst : DFF_X1 port map( D => n10831, CK => CLK, Q => 
                           n2097, QN => n7430);
   REGISTERS_reg_51_28_inst : DFF_X1 port map( D => n10832, CK => CLK, Q => 
                           n2098, QN => n7406);
   REGISTERS_reg_51_27_inst : DFF_X1 port map( D => n10833, CK => CLK, Q => 
                           n2099, QN => n7382);
   REGISTERS_reg_51_26_inst : DFF_X1 port map( D => n10834, CK => CLK, Q => 
                           n2100, QN => n7358);
   REGISTERS_reg_51_25_inst : DFF_X1 port map( D => n10835, CK => CLK, Q => 
                           n2101, QN => n7334);
   REGISTERS_reg_51_24_inst : DFF_X1 port map( D => n10836, CK => CLK, Q => 
                           n2102, QN => n7310);
   REGISTERS_reg_51_23_inst : DFF_X1 port map( D => n10837, CK => CLK, Q => 
                           n2103, QN => n7286);
   REGISTERS_reg_51_22_inst : DFF_X1 port map( D => n10838, CK => CLK, Q => 
                           n2104, QN => n7262);
   REGISTERS_reg_51_21_inst : DFF_X1 port map( D => n10839, CK => CLK, Q => 
                           n2105, QN => n7238);
   REGISTERS_reg_51_19_inst : DFF_X1 port map( D => n10841, CK => CLK, Q => 
                           n2107, QN => n7190);
   REGISTERS_reg_51_18_inst : DFF_X1 port map( D => n10842, CK => CLK, Q => 
                           n2108, QN => n7166);
   REGISTERS_reg_51_17_inst : DFF_X1 port map( D => n10843, CK => CLK, Q => 
                           n2109, QN => n7142);
   REGISTERS_reg_51_16_inst : DFF_X1 port map( D => n10844, CK => CLK, Q => 
                           n2110, QN => n7118);
   REGISTERS_reg_51_15_inst : DFF_X1 port map( D => n10845, CK => CLK, Q => 
                           n2111, QN => n7094);
   REGISTERS_reg_51_14_inst : DFF_X1 port map( D => n10846, CK => CLK, Q => 
                           n2112, QN => n7070);
   REGISTERS_reg_51_13_inst : DFF_X1 port map( D => n10847, CK => CLK, Q => 
                           n2113, QN => n7046);
   REGISTERS_reg_51_12_inst : DFF_X1 port map( D => n10848, CK => CLK, Q => 
                           n2114, QN => n7022);
   REGISTERS_reg_51_11_inst : DFF_X1 port map( D => n10849, CK => CLK, Q => 
                           n2115, QN => n6998);
   REGISTERS_reg_51_10_inst : DFF_X1 port map( D => n10850, CK => CLK, Q => 
                           n2116, QN => n6974);
   REGISTERS_reg_51_9_inst : DFF_X1 port map( D => n10851, CK => CLK, Q => 
                           n2117, QN => n6950);
   REGISTERS_reg_51_8_inst : DFF_X1 port map( D => n10852, CK => CLK, Q => 
                           n2118, QN => n6926);
   REGISTERS_reg_42_31_inst : DFF_X1 port map( D => n10541, CK => CLK, Q => 
                           n2280, QN => n7481);
   REGISTERS_reg_42_30_inst : DFF_X1 port map( D => n10542, CK => CLK, Q => 
                           n2281, QN => n7457);
   REGISTERS_reg_42_29_inst : DFF_X1 port map( D => n10543, CK => CLK, Q => 
                           n2282, QN => n7433);
   REGISTERS_reg_42_28_inst : DFF_X1 port map( D => n10544, CK => CLK, Q => 
                           n2283, QN => n7409);
   REGISTERS_reg_42_27_inst : DFF_X1 port map( D => n10545, CK => CLK, Q => 
                           n2284, QN => n7385);
   REGISTERS_reg_42_26_inst : DFF_X1 port map( D => n10546, CK => CLK, Q => 
                           n2285, QN => n7361);
   REGISTERS_reg_42_25_inst : DFF_X1 port map( D => n10547, CK => CLK, Q => 
                           n2286, QN => n7337);
   REGISTERS_reg_42_24_inst : DFF_X1 port map( D => n10548, CK => CLK, Q => 
                           n2287, QN => n7313);
   REGISTERS_reg_42_23_inst : DFF_X1 port map( D => n10549, CK => CLK, Q => 
                           n2288, QN => n7289);
   REGISTERS_reg_42_22_inst : DFF_X1 port map( D => n10550, CK => CLK, Q => 
                           n2289, QN => n7265);
   REGISTERS_reg_42_21_inst : DFF_X1 port map( D => n10551, CK => CLK, Q => 
                           n2290, QN => n7241);
   REGISTERS_reg_42_19_inst : DFF_X1 port map( D => n10553, CK => CLK, Q => 
                           n2292, QN => n7193);
   REGISTERS_reg_42_18_inst : DFF_X1 port map( D => n10554, CK => CLK, Q => 
                           n2293, QN => n7169);
   REGISTERS_reg_42_17_inst : DFF_X1 port map( D => n10555, CK => CLK, Q => 
                           n2294, QN => n7145);
   REGISTERS_reg_42_16_inst : DFF_X1 port map( D => n10556, CK => CLK, Q => 
                           n2295, QN => n7121);
   REGISTERS_reg_42_15_inst : DFF_X1 port map( D => n10557, CK => CLK, Q => 
                           n2296, QN => n7097);
   REGISTERS_reg_42_14_inst : DFF_X1 port map( D => n10558, CK => CLK, Q => 
                           n2297, QN => n7073);
   REGISTERS_reg_42_13_inst : DFF_X1 port map( D => n10559, CK => CLK, Q => 
                           n2298, QN => n7049);
   REGISTERS_reg_42_12_inst : DFF_X1 port map( D => n10560, CK => CLK, Q => 
                           n2299, QN => n7025);
   REGISTERS_reg_42_11_inst : DFF_X1 port map( D => n10561, CK => CLK, Q => 
                           n2300, QN => n7001);
   REGISTERS_reg_42_10_inst : DFF_X1 port map( D => n10562, CK => CLK, Q => 
                           n2301, QN => n6977);
   REGISTERS_reg_42_9_inst : DFF_X1 port map( D => n10563, CK => CLK, Q => 
                           n2302, QN => n6953);
   REGISTERS_reg_42_8_inst : DFF_X1 port map( D => n10564, CK => CLK, Q => 
                           n2303, QN => n6929);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n10446, CK => CLK, Q => 
                           n2304, QN => n7693);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n10447, CK => CLK, Q => 
                           n2305, QN => n7697);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n10448, CK => CLK, Q => 
                           n2306, QN => n7701);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n10449, CK => CLK, Q => 
                           n2307, QN => n7705);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n10450, CK => CLK, Q => 
                           n2308, QN => n7709);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n10451, CK => CLK, Q => 
                           n2309, QN => n7713);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n10452, CK => CLK, Q => 
                           n2310, QN => n7717);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n10453, CK => CLK, Q => 
                           n2311, QN => n7721);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n10454, CK => CLK, Q => 
                           n2312, QN => n7725);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n10455, CK => CLK, Q => 
                           n2313, QN => n7729);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n10457, CK => CLK, Q => 
                           n2315, QN => n7737);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n10458, CK => CLK, Q => 
                           n2316, QN => n7741);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n10459, CK => CLK, Q => 
                           n2317, QN => n7745);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n10460, CK => CLK, Q => 
                           n2318, QN => n7749);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n10461, CK => CLK, Q => 
                           n2319, QN => n7753);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n10462, CK => CLK, Q => 
                           n2320, QN => n7757);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n10463, CK => CLK, Q => 
                           n2321, QN => n7761);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n10464, CK => CLK, Q => 
                           n2322, QN => n7765);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n10465, CK => CLK, Q => 
                           n2323, QN => n7769);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n10466, CK => CLK, Q => 
                           n2324, QN => n7773);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n10467, CK => CLK, Q => 
                           n2325, QN => n7777);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n10468, CK => CLK, Q => 
                           n2326, QN => n7781);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n10413, CK => CLK, Q => 
                           n2327, QN => n7688);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n10414, CK => CLK, Q => 
                           n2328, QN => n7692);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n10415, CK => CLK, Q => 
                           n2329, QN => n7696);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n10416, CK => CLK, Q => 
                           n2330, QN => n7700);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n10417, CK => CLK, Q => 
                           n2331, QN => n7704);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n10418, CK => CLK, Q => 
                           n2332, QN => n7708);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n10419, CK => CLK, Q => 
                           n2333, QN => n7712);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n10420, CK => CLK, Q => 
                           n2334, QN => n7716);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n10421, CK => CLK, Q => 
                           n2335, QN => n7720);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n10422, CK => CLK, Q => 
                           n2336, QN => n7724);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n10423, CK => CLK, Q => 
                           n2337, QN => n7728);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n10424, CK => CLK, Q => 
                           n2338, QN => n7732);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n10425, CK => CLK, Q => 
                           n2339, QN => n7736);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n10426, CK => CLK, Q => 
                           n2340, QN => n7740);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n10427, CK => CLK, Q => 
                           n2341, QN => n7744);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n10428, CK => CLK, Q => 
                           n2342, QN => n7748);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n10429, CK => CLK, Q => 
                           n2343, QN => n7752);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n10430, CK => CLK, Q => 
                           n2344, QN => n7756);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n10431, CK => CLK, Q => 
                           n2345, QN => n7760);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n10432, CK => CLK, Q => 
                           n2346, QN => n7764);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n10433, CK => CLK, Q => 
                           n2347, QN => n7768);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n10434, CK => CLK, Q => 
                           n2348, QN => n7772);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n10435, CK => CLK, Q => 
                           n2349, QN => n7776);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n10436, CK => CLK, Q => 
                           n2350, QN => n7780);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n10331, CK => CLK, Q => 
                           n_1646, QN => n7146);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n10337, CK => CLK, Q => 
                           n_1647, QN => n7002);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n10338, CK => CLK, Q => 
                           n_1648, QN => n6978);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n10339, CK => CLK, Q => 
                           n_1649, QN => n6954);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n10340, CK => CLK, Q => 
                           n_1650, QN => n6930);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n10253, CK => CLK, Q => 
                           n2379, QN => n7484);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n10254, CK => CLK, Q => 
                           n2380, QN => n7460);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n10255, CK => CLK, Q => 
                           n2381, QN => n7436);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n10256, CK => CLK, Q => 
                           n2382, QN => n7412);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n10257, CK => CLK, Q => 
                           n2383, QN => n7388);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n10258, CK => CLK, Q => 
                           n2384, QN => n7364);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n10259, CK => CLK, Q => 
                           n2385, QN => n7340);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n10260, CK => CLK, Q => 
                           n2386, QN => n7316);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n10261, CK => CLK, Q => 
                           n2387, QN => n7292);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n10262, CK => CLK, Q => 
                           n2388, QN => n7268);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n10263, CK => CLK, Q => 
                           n2389, QN => n7244);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n10265, CK => CLK, Q => 
                           n2391, QN => n7196);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n10266, CK => CLK, Q => 
                           n2392, QN => n7172);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n10267, CK => CLK, Q => 
                           n2393, QN => n7148);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n10268, CK => CLK, Q => 
                           n2394, QN => n7124);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n10269, CK => CLK, Q => 
                           n2395, QN => n7100);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n10270, CK => CLK, Q => 
                           n2396, QN => n7076);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n10271, CK => CLK, Q => 
                           n2397, QN => n7052);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n10272, CK => CLK, Q => 
                           n2398, QN => n7028);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n10273, CK => CLK, Q => 
                           n2399, QN => n7004);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n10274, CK => CLK, Q => 
                           n2400, QN => n6980);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n10275, CK => CLK, Q => 
                           n2401, QN => n6956);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n10276, CK => CLK, Q => 
                           n2402, QN => n6932);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n9680, CK => CLK, Q => 
                           n2484, QN => n7418);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n9872, CK => CLK, Q => 
                           n2485, QN => n7703);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n9840, CK => CLK, Q => 
                           n2486, QN => n7702);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n9744, CK => CLK, Q => 
                           n_1651, QN => n7416);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n9712, CK => CLK, Q => 
                           n_1652, QN => n7417);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n10029, CK => CLK, Q => 
                           n_1653, QN => n7485);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n10051, CK => CLK, Q => 
                           n_1654, QN => n6957);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n10052, CK => CLK, Q => 
                           n_1655, QN => n6933);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n10053, CK => CLK, Q => 
                           n_1656, QN => n6909);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n10054, CK => CLK, Q => 
                           n_1657, QN => n6885);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n10055, CK => CLK, Q => 
                           n_1658, QN => n6861);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n10056, CK => CLK, Q => 
                           n_1659, QN => n6837);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n10057, CK => CLK, Q => 
                           n_1660, QN => n6813);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n10058, CK => CLK, Q => 
                           n_1661, QN => n6789);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n10059, CK => CLK, Q => 
                           n_1662, QN => n6765);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n9681, CK => CLK, Q => 
                           n2411, QN => n7394);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n9682, CK => CLK, Q => 
                           n2412, QN => n7370);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n9683, CK => CLK, Q => 
                           n2413, QN => n7346);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n9684, CK => CLK, Q => 
                           n2414, QN => n7322);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n9685, CK => CLK, Q => 
                           n2415, QN => n7298);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n9686, CK => CLK, Q => 
                           n2416, QN => n7274);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n9687, CK => CLK, Q => 
                           n2417, QN => n7250);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n9690, CK => CLK, Q => 
                           n2420, QN => n7178);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n9691, CK => CLK, Q => 
                           n2421, QN => n7154);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n9692, CK => CLK, Q => 
                           n2422, QN => n7130);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n9693, CK => CLK, Q => 
                           n2423, QN => n7106);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n9694, CK => CLK, Q => 
                           n2424, QN => n7082);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n9695, CK => CLK, Q => 
                           n2425, QN => n7058);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n9696, CK => CLK, Q => 
                           n2426, QN => n7034);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n9697, CK => CLK, Q => 
                           n2427, QN => n7010);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n9698, CK => CLK, Q => 
                           n2428, QN => n6986);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n9699, CK => CLK, Q => n2429
                           , QN => n6962);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n9700, CK => CLK, Q => n2430
                           , QN => n6938);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n10042, CK => CLK, Q => 
                           n_1663, QN => n7173);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n10043, CK => CLK, Q => 
                           n_1664, QN => n7149);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n10048, CK => CLK, Q => 
                           n_1665, QN => n7029);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n10049, CK => CLK, Q => 
                           n_1666, QN => n7005);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n10050, CK => CLK, Q => 
                           n_1667, QN => n6981);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n10060, CK => CLK, Q => 
                           n_1668, QN => n6741);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n9965, CK => CLK, Q => 
                           n2437, QN => n7487);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n9945, CK => CLK, Q => 
                           n1617, QN => n824);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n9913, CK => CLK, Q => 
                           n1638, QN => n823);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n9869, CK => CLK, Q => 
                           n2438, QN => n7691);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n9873, CK => CLK, Q => 
                           n2439, QN => n7707);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n9874, CK => CLK, Q => 
                           n2440, QN => n7711);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n9875, CK => CLK, Q => 
                           n2441, QN => n7715);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n9876, CK => CLK, Q => 
                           n2442, QN => n7719);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n9877, CK => CLK, Q => 
                           n2443, QN => n7723);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n9878, CK => CLK, Q => 
                           n2444, QN => n7727);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n9879, CK => CLK, Q => 
                           n2445, QN => n7731);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n9880, CK => CLK, Q => 
                           n2446, QN => n7735);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n9882, CK => CLK, Q => 
                           n2448, QN => n7743);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n9883, CK => CLK, Q => 
                           n2449, QN => n7747);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n9884, CK => CLK, Q => 
                           n2450, QN => n7751);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n9885, CK => CLK, Q => 
                           n2451, QN => n7755);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n9886, CK => CLK, Q => 
                           n2452, QN => n7759);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n9887, CK => CLK, Q => 
                           n2453, QN => n7763);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n9888, CK => CLK, Q => 
                           n2454, QN => n7767);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n9889, CK => CLK, Q => 
                           n2455, QN => n7771);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n9890, CK => CLK, Q => 
                           n2456, QN => n7775);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n9891, CK => CLK, Q => n2457
                           , QN => n7779);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n9892, CK => CLK, Q => n2458
                           , QN => n7783);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n9837, CK => CLK, Q => 
                           n2459, QN => n7690);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n9841, CK => CLK, Q => 
                           n2460, QN => n7706);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n9842, CK => CLK, Q => 
                           n2461, QN => n7710);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n9843, CK => CLK, Q => 
                           n2462, QN => n7714);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n9844, CK => CLK, Q => 
                           n2463, QN => n7718);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n9845, CK => CLK, Q => 
                           n2464, QN => n7722);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n9846, CK => CLK, Q => 
                           n2465, QN => n7726);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n9847, CK => CLK, Q => 
                           n2466, QN => n7730);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n9848, CK => CLK, Q => 
                           n2467, QN => n7734);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n9850, CK => CLK, Q => 
                           n2469, QN => n7742);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n9851, CK => CLK, Q => 
                           n2470, QN => n7746);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n9852, CK => CLK, Q => 
                           n2471, QN => n7750);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n9853, CK => CLK, Q => 
                           n2472, QN => n7754);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n9854, CK => CLK, Q => 
                           n2473, QN => n7758);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n9855, CK => CLK, Q => 
                           n2474, QN => n7762);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n9856, CK => CLK, Q => 
                           n2475, QN => n7766);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n9857, CK => CLK, Q => 
                           n2476, QN => n7770);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n9858, CK => CLK, Q => 
                           n2477, QN => n7774);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n9859, CK => CLK, Q => n2478
                           , QN => n7778);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n9860, CK => CLK, Q => n2479
                           , QN => n7782);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n9816, CK => CLK, Q => 
                           n1658, QN => n756);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n9817, CK => CLK, Q => 
                           n1659, QN => n820);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n9741, CK => CLK, Q => 
                           n_1669, QN => n7488);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n9745, CK => CLK, Q => 
                           n_1670, QN => n7392);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n9746, CK => CLK, Q => 
                           n_1671, QN => n7368);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n9747, CK => CLK, Q => 
                           n_1672, QN => n7344);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n9748, CK => CLK, Q => 
                           n_1673, QN => n7320);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n9749, CK => CLK, Q => 
                           n_1674, QN => n7296);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n9750, CK => CLK, Q => 
                           n_1675, QN => n7272);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n9751, CK => CLK, Q => 
                           n_1676, QN => n7248);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n9754, CK => CLK, Q => 
                           n_1677, QN => n7176);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n9755, CK => CLK, Q => 
                           n_1678, QN => n7152);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n9761, CK => CLK, Q => 
                           n_1679, QN => n7008);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n9762, CK => CLK, Q => 
                           n_1680, QN => n6984);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n9763, CK => CLK, Q => 
                           n_1681, QN => n6960);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n9764, CK => CLK, Q => 
                           n_1682, QN => n6936);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n9709, CK => CLK, Q => 
                           n_1683, QN => n7489);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n9713, CK => CLK, Q => 
                           n_1684, QN => n7393);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n9714, CK => CLK, Q => 
                           n_1685, QN => n7369);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n9715, CK => CLK, Q => 
                           n_1686, QN => n7345);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n9716, CK => CLK, Q => 
                           n_1687, QN => n7321);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n9717, CK => CLK, Q => 
                           n_1688, QN => n7297);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n9718, CK => CLK, Q => 
                           n_1689, QN => n7273);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n9719, CK => CLK, Q => 
                           n_1690, QN => n7249);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n9722, CK => CLK, Q => 
                           n_1691, QN => n7177);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n9966, CK => CLK, Q => 
                           n2405, QN => n7463);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n9967, CK => CLK, Q => 
                           n2406, QN => n7439);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n9870, CK => CLK, Q => 
                           n2407, QN => n7695);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n9871, CK => CLK, Q => 
                           n2408, QN => n7699);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n9838, CK => CLK, Q => 
                           n2409, QN => n7694);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n9839, CK => CLK, Q => 
                           n2410, QN => n7698);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n9710, CK => CLK, Q => 
                           n_1692, QN => n7465);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n9711, CK => CLK, Q => 
                           n_1693, QN => n7441);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n10001, CK => CLK, Q => 
                           n_1694, QN => n7390);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n10002, CK => CLK, Q => 
                           n_1695, QN => n7366);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n10003, CK => CLK, Q => 
                           n_1696, QN => n7342);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n10004, CK => CLK, Q => 
                           n_1697, QN => n7318);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n10005, CK => CLK, Q => 
                           n_1698, QN => n7294);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n10030, CK => CLK, Q => 
                           n_1699, QN => n7461);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n10031, CK => CLK, Q => 
                           n_1700, QN => n7437);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n9997, CK => CLK, Q => 
                           n_1701, QN => n7486);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n10020, CK => CLK, Q => 
                           n_1702, QN => n6934);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n10021, CK => CLK, Q => 
                           n_1703, QN => n6910);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n10022, CK => CLK, Q => 
                           n_1704, QN => n6886);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n10023, CK => CLK, Q => 
                           n_1705, QN => n6862);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n10024, CK => CLK, Q => 
                           n_1706, QN => n6838);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n10025, CK => CLK, Q => 
                           n_1707, QN => n6814);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n10026, CK => CLK, Q => 
                           n_1708, QN => n6790);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n10027, CK => CLK, Q => 
                           n_1709, QN => n6766);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n10028, CK => CLK, Q => 
                           n_1710, QN => n6742);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n10006, CK => CLK, Q => 
                           n_1711, QN => n7270);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n10007, CK => CLK, Q => 
                           n_1712, QN => n7246);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n10010, CK => CLK, Q => 
                           n_1713, QN => n7174);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n10011, CK => CLK, Q => 
                           n_1714, QN => n7150);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n10012, CK => CLK, Q => 
                           n2433, QN => n7126);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n10013, CK => CLK, Q => 
                           n2434, QN => n7102);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n10014, CK => CLK, Q => 
                           n2435, QN => n7078);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n10015, CK => CLK, Q => 
                           n2436, QN => n7054);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n10016, CK => CLK, Q => 
                           n_1715, QN => n7030);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n10017, CK => CLK, Q => 
                           n_1716, QN => n7006);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n10018, CK => CLK, Q => 
                           n_1717, QN => n6982);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n10019, CK => CLK, Q => 
                           n_1718, QN => n6958);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n9998, CK => CLK, Q => 
                           n_1719, QN => n7462);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n9999, CK => CLK, Q => 
                           n_1720, QN => n7438);
   REGISTERS_reg_71_7_inst : DFF_X1 port map( D => n11493, CK => CLK, Q => 
                           n2487, QN => n6894);
   REGISTERS_reg_71_6_inst : DFF_X1 port map( D => n11494, CK => CLK, Q => 
                           n2488, QN => n6870);
   REGISTERS_reg_71_5_inst : DFF_X1 port map( D => n11495, CK => CLK, Q => 
                           n2489, QN => n6846);
   REGISTERS_reg_71_4_inst : DFF_X1 port map( D => n11496, CK => CLK, Q => 
                           n2490, QN => n6822);
   REGISTERS_reg_71_3_inst : DFF_X1 port map( D => n11497, CK => CLK, Q => 
                           n2491, QN => n6798);
   REGISTERS_reg_71_2_inst : DFF_X1 port map( D => n11498, CK => CLK, Q => 
                           n2492, QN => n6774);
   REGISTERS_reg_71_1_inst : DFF_X1 port map( D => n11499, CK => CLK, Q => 
                           n2493, QN => n6750);
   REGISTERS_reg_71_0_inst : DFF_X1 port map( D => n11500, CK => CLK, Q => 
                           n2494, QN => n6726);
   REGISTERS_reg_71_28_inst : DFF_X1 port map( D => n11472, CK => CLK, Q => 
                           n2520, QN => n7398);
   REGISTERS_reg_71_31_inst : DFF_X1 port map( D => n11469, CK => CLK, Q => 
                           n2498, QN => n7470);
   REGISTERS_reg_71_27_inst : DFF_X1 port map( D => n11473, CK => CLK, Q => 
                           n2499, QN => n7374);
   REGISTERS_reg_71_26_inst : DFF_X1 port map( D => n11474, CK => CLK, Q => 
                           n2500, QN => n7350);
   REGISTERS_reg_71_25_inst : DFF_X1 port map( D => n11475, CK => CLK, Q => 
                           n2501, QN => n7326);
   REGISTERS_reg_71_24_inst : DFF_X1 port map( D => n11476, CK => CLK, Q => 
                           n2502, QN => n7302);
   REGISTERS_reg_71_23_inst : DFF_X1 port map( D => n11477, CK => CLK, Q => 
                           n2503, QN => n7278);
   REGISTERS_reg_71_22_inst : DFF_X1 port map( D => n11478, CK => CLK, Q => 
                           n2504, QN => n7254);
   REGISTERS_reg_71_19_inst : DFF_X1 port map( D => n11481, CK => CLK, Q => 
                           n2507, QN => n7182);
   REGISTERS_reg_71_18_inst : DFF_X1 port map( D => n11482, CK => CLK, Q => 
                           n2508, QN => n7158);
   REGISTERS_reg_71_17_inst : DFF_X1 port map( D => n11483, CK => CLK, Q => 
                           n2509, QN => n7134);
   REGISTERS_reg_71_16_inst : DFF_X1 port map( D => n11484, CK => CLK, Q => 
                           n2510, QN => n7110);
   REGISTERS_reg_71_15_inst : DFF_X1 port map( D => n11485, CK => CLK, Q => 
                           n2511, QN => n7086);
   REGISTERS_reg_71_14_inst : DFF_X1 port map( D => n11486, CK => CLK, Q => 
                           n2512, QN => n7062);
   REGISTERS_reg_71_13_inst : DFF_X1 port map( D => n11487, CK => CLK, Q => 
                           n2513, QN => n7038);
   REGISTERS_reg_71_12_inst : DFF_X1 port map( D => n11488, CK => CLK, Q => 
                           n2514, QN => n7014);
   REGISTERS_reg_71_11_inst : DFF_X1 port map( D => n11489, CK => CLK, Q => 
                           n2515, QN => n6990);
   REGISTERS_reg_71_10_inst : DFF_X1 port map( D => n11490, CK => CLK, Q => 
                           n2516, QN => n6966);
   REGISTERS_reg_71_9_inst : DFF_X1 port map( D => n11491, CK => CLK, Q => 
                           n2517, QN => n6942);
   REGISTERS_reg_71_8_inst : DFF_X1 port map( D => n11492, CK => CLK, Q => 
                           n2518, QN => n6918);
   REGISTERS_reg_71_30_inst : DFF_X1 port map( D => n11470, CK => CLK, Q => 
                           n2495, QN => n7446);
   REGISTERS_reg_71_29_inst : DFF_X1 port map( D => n11471, CK => CLK, Q => 
                           n2496, QN => n7422);
   OUT2_reg_6_inst : DFF_X1 port map( D => n9127, CK => CLK, Q => n_1721, QN =>
                           n2188);
   OUT2_reg_5_inst : DFF_X1 port map( D => n9128, CK => CLK, Q => n_1722, QN =>
                           n2187);
   OUT2_reg_4_inst : DFF_X1 port map( D => n9129, CK => CLK, Q => n_1723, QN =>
                           n2186);
   OUT2_reg_3_inst : DFF_X1 port map( D => n9130, CK => CLK, Q => n_1724, QN =>
                           n2185);
   OUT2_reg_2_inst : DFF_X1 port map( D => n9131, CK => CLK, Q => n_1725, QN =>
                           n2184);
   OUT2_reg_1_inst : DFF_X1 port map( D => n9132, CK => CLK, Q => n_1726, QN =>
                           n2183);
   OUT2_reg_0_inst : DFF_X1 port map( D => n9133, CK => CLK, Q => n_1727, QN =>
                           n2182);
   OUT1_reg_6_inst : DFF_X1 port map( D => n9160, CK => CLK, Q => n_1728, QN =>
                           n2156);
   OUT1_reg_5_inst : DFF_X1 port map( D => n9161, CK => CLK, Q => n_1729, QN =>
                           n2155);
   OUT1_reg_4_inst : DFF_X1 port map( D => n9162, CK => CLK, Q => n_1730, QN =>
                           n2154);
   OUT1_reg_3_inst : DFF_X1 port map( D => n9163, CK => CLK, Q => n_1731, QN =>
                           n2153);
   OUT1_reg_2_inst : DFF_X1 port map( D => n9164, CK => CLK, Q => n_1732, QN =>
                           n2152);
   OUT1_reg_1_inst : DFF_X1 port map( D => n9165, CK => CLK, Q => n_1733, QN =>
                           n2151);
   OUT1_reg_0_inst : DFF_X1 port map( D => n9166, CK => CLK, Q => n_1734, QN =>
                           n2150);
   OUT2_reg_7_inst : DFF_X1 port map( D => n9126, CK => CLK, Q => n_1735, QN =>
                           n2189);
   OUT1_reg_7_inst : DFF_X1 port map( D => n9159, CK => CLK, Q => n_1736, QN =>
                           n2157);
   OUT2_reg_19_inst : DFF_X1 port map( D => n9114, CK => CLK, Q => n_1737, QN 
                           => n2201);
   OUT1_reg_19_inst : DFF_X1 port map( D => n9147, CK => CLK, Q => n_1738, QN 
                           => n2169);
   OUT2_reg_18_inst : DFF_X1 port map( D => n9115, CK => CLK, Q => n_1739, QN 
                           => n2200);
   OUT2_reg_17_inst : DFF_X1 port map( D => n9116, CK => CLK, Q => n_1740, QN 
                           => n2199);
   OUT2_reg_16_inst : DFF_X1 port map( D => n9117, CK => CLK, Q => n_1741, QN 
                           => n2198);
   OUT2_reg_15_inst : DFF_X1 port map( D => n9118, CK => CLK, Q => n_1742, QN 
                           => n2197);
   OUT2_reg_14_inst : DFF_X1 port map( D => n9119, CK => CLK, Q => n_1743, QN 
                           => n2196);
   OUT2_reg_13_inst : DFF_X1 port map( D => n9120, CK => CLK, Q => n_1744, QN 
                           => n2195);
   OUT2_reg_12_inst : DFF_X1 port map( D => n9121, CK => CLK, Q => n_1745, QN 
                           => n2194);
   OUT2_reg_11_inst : DFF_X1 port map( D => n9122, CK => CLK, Q => n_1746, QN 
                           => n2193);
   OUT2_reg_10_inst : DFF_X1 port map( D => n9123, CK => CLK, Q => n_1747, QN 
                           => n2192);
   OUT2_reg_9_inst : DFF_X1 port map( D => n9124, CK => CLK, Q => n_1748, QN =>
                           n2191);
   OUT2_reg_8_inst : DFF_X1 port map( D => n9125, CK => CLK, Q => n_1749, QN =>
                           n2190);
   OUT1_reg_18_inst : DFF_X1 port map( D => n9148, CK => CLK, Q => n_1750, QN 
                           => n2168);
   OUT1_reg_17_inst : DFF_X1 port map( D => n9149, CK => CLK, Q => n_1751, QN 
                           => n2167);
   OUT1_reg_16_inst : DFF_X1 port map( D => n9150, CK => CLK, Q => n_1752, QN 
                           => n2166);
   OUT1_reg_15_inst : DFF_X1 port map( D => n9151, CK => CLK, Q => n_1753, QN 
                           => n2165);
   OUT1_reg_14_inst : DFF_X1 port map( D => n9152, CK => CLK, Q => n_1754, QN 
                           => n2164);
   OUT1_reg_13_inst : DFF_X1 port map( D => n9153, CK => CLK, Q => n_1755, QN 
                           => n2163);
   OUT1_reg_12_inst : DFF_X1 port map( D => n9154, CK => CLK, Q => n_1756, QN 
                           => n2162);
   OUT1_reg_11_inst : DFF_X1 port map( D => n9155, CK => CLK, Q => n_1757, QN 
                           => n2161);
   OUT1_reg_10_inst : DFF_X1 port map( D => n9156, CK => CLK, Q => n_1758, QN 
                           => n2160);
   OUT1_reg_9_inst : DFF_X1 port map( D => n9157, CK => CLK, Q => n_1759, QN =>
                           n2159);
   OUT1_reg_8_inst : DFF_X1 port map( D => n9158, CK => CLK, Q => n_1760, QN =>
                           n2158);
   OUT2_reg_31_inst : DFF_X1 port map( D => n9102, CK => CLK, Q => n_1761, QN 
                           => n2213);
   OUT2_reg_30_inst : DFF_X1 port map( D => n9103, CK => CLK, Q => n_1762, QN 
                           => n2212);
   OUT2_reg_29_inst : DFF_X1 port map( D => n9104, CK => CLK, Q => n_1763, QN 
                           => n2211);
   OUT2_reg_28_inst : DFF_X1 port map( D => n9105, CK => CLK, Q => n_1764, QN 
                           => n2210);
   OUT2_reg_27_inst : DFF_X1 port map( D => n9106, CK => CLK, Q => n_1765, QN 
                           => n2209);
   OUT2_reg_26_inst : DFF_X1 port map( D => n9107, CK => CLK, Q => n_1766, QN 
                           => n2208);
   OUT2_reg_25_inst : DFF_X1 port map( D => n9108, CK => CLK, Q => n_1767, QN 
                           => n2207);
   OUT2_reg_24_inst : DFF_X1 port map( D => n9109, CK => CLK, Q => n_1768, QN 
                           => n2206);
   OUT2_reg_23_inst : DFF_X1 port map( D => n9110, CK => CLK, Q => n_1769, QN 
                           => n2205);
   OUT2_reg_22_inst : DFF_X1 port map( D => n9111, CK => CLK, Q => n_1770, QN 
                           => n2204);
   OUT2_reg_21_inst : DFF_X1 port map( D => n9112, CK => CLK, Q => n_1771, QN 
                           => n2203);
   OUT2_reg_20_inst : DFF_X1 port map( D => n9113, CK => CLK, Q => n_1772, QN 
                           => n2202);
   OUT1_reg_31_inst : DFF_X1 port map( D => n9135, CK => CLK, Q => n_1773, QN 
                           => n2181);
   OUT1_reg_30_inst : DFF_X1 port map( D => n9136, CK => CLK, Q => n_1774, QN 
                           => n2180);
   OUT1_reg_29_inst : DFF_X1 port map( D => n9137, CK => CLK, Q => n_1775, QN 
                           => n2179);
   OUT1_reg_28_inst : DFF_X1 port map( D => n9138, CK => CLK, Q => n_1776, QN 
                           => n2178);
   OUT1_reg_27_inst : DFF_X1 port map( D => n9139, CK => CLK, Q => n_1777, QN 
                           => n2177);
   OUT1_reg_26_inst : DFF_X1 port map( D => n9140, CK => CLK, Q => n_1778, QN 
                           => n2176);
   OUT1_reg_25_inst : DFF_X1 port map( D => n9141, CK => CLK, Q => n_1779, QN 
                           => n2175);
   OUT1_reg_24_inst : DFF_X1 port map( D => n9142, CK => CLK, Q => n_1780, QN 
                           => n2174);
   OUT1_reg_23_inst : DFF_X1 port map( D => n9143, CK => CLK, Q => n_1781, QN 
                           => n2173);
   U3 : NOR3_X1 port map( A1 => n2551, A2 => ADD_RD2(4), A3 => n2549, ZN => 
                           n6538);
   U4 : NOR3_X1 port map( A1 => n2550, A2 => ADD_RD2(3), A3 => n2549, ZN => 
                           n6536);
   U5 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), A3 => n2551, ZN 
                           => n6509);
   U6 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n2549, ZN 
                           => n6526);
   U7 : NOR3_X1 port map( A1 => n2553, A2 => ADD_RD2(0), A3 => n2552, ZN => 
                           n6513);
   U8 : NOR3_X1 port map( A1 => n2551, A2 => ADD_RD2(5), A3 => n2550, ZN => 
                           n6527);
   U9 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(5), A3 => n2550, ZN 
                           => n6507);
   U10 : NOR3_X1 port map( A1 => n2545, A2 => ADD_RD1(4), A3 => n2543, ZN => 
                           n5217);
   U11 : NOR3_X1 port map( A1 => n2544, A2 => ADD_RD1(3), A3 => n2543, ZN => 
                           n5215);
   U12 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), A3 => n2545, ZN 
                           => n5188);
   U13 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => ADD_RD1(0)
                           , ZN => n5187);
   U14 : NOR3_X1 port map( A1 => n2545, A2 => ADD_RD1(5), A3 => n2544, ZN => 
                           n5206);
   U15 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(5), A3 => n2544, ZN 
                           => n5186);
   U16 : NAND2_X1 port map( A1 => n6591, A2 => n6680, ZN => n2660);
   U17 : NAND2_X1 port map( A1 => n6582, A2 => n6680, ZN => n6684);
   U18 : NAND2_X1 port map( A1 => n6569, A2 => n6680, ZN => n6633);
   U19 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n2543, ZN 
                           => n5205);
   U20 : NOR2_X1 port map( A1 => n2563, A2 => ADD_SF(6), ZN => n2744);
   U85 : NOR2_X2 port map( A1 => n2569, A2 => ADD_SF(5), ZN => n6591);
   U86 : AND2_X1 port map( A1 => n5205, A2 => n5194, ZN => n13220);
   U87 : AND2_X1 port map( A1 => n2744, A2 => n2573, ZN => n13221);
   U88 : AND3_X1 port map( A1 => n2534, A2 => n2533, A3 => n3953, ZN => n2710);
   U89 : NOR3_X1 port map( A1 => n2548, A2 => ADD_RD1(1), A3 => n2546, ZN => 
                           n5191);
   U90 : NOR3_X1 port map( A1 => n2554, A2 => ADD_RD2(1), A3 => n2552, ZN => 
                           n6512);
   U91 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n2548, ZN 
                           => n5190);
   U92 : AND3_X1 port map( A1 => n3953, A2 => n2533, A3 => ADD_WR(4), ZN => 
                           n2663);
   U93 : BUF_X1 port map( A => n2625, Z => n14705);
   U94 : BUF_X1 port map( A => n2625, Z => n14704);
   U95 : BUF_X1 port map( A => n6821, Z => n13232);
   U96 : BUF_X1 port map( A => n6748, Z => n13296);
   U97 : BUF_X1 port map( A => n6748, Z => n13295);
   U98 : BUF_X1 port map( A => n6738, Z => n13304);
   U99 : BUF_X1 port map( A => n6732, Z => n13313);
   U100 : BUF_X1 port map( A => n6716, Z => n13341);
   U101 : BUF_X1 port map( A => n6716, Z => n13340);
   U102 : BUF_X1 port map( A => n6710, Z => n13350);
   U103 : BUF_X1 port map( A => n6698, Z => n13377);
   U104 : BUF_X1 port map( A => n6698, Z => n13376);
   U105 : BUF_X1 port map( A => n6695, Z => n13385);
   U106 : BUF_X1 port map( A => n6692, Z => n13394);
   U107 : BUF_X1 port map( A => n6668, Z => n13458);
   U108 : BUF_X1 port map( A => n6668, Z => n13457);
   U109 : BUF_X1 port map( A => n6665, Z => n13466);
   U110 : BUF_X1 port map( A => n6662, Z => n13475);
   U111 : BUF_X1 port map( A => n6641, Z => n13539);
   U112 : BUF_X1 port map( A => n6641, Z => n13538);
   U113 : BUF_X1 port map( A => n6638, Z => n13547);
   U114 : BUF_X1 port map( A => n6635, Z => n13556);
   U115 : BUF_X1 port map( A => n6753, Z => n13287);
   U116 : BUF_X1 port map( A => n6753, Z => n13286);
   U117 : BUF_X1 port map( A => n6738, Z => n13305);
   U118 : BUF_X1 port map( A => n6732, Z => n13314);
   U119 : BUF_X1 port map( A => n6725, Z => n13323);
   U120 : BUF_X1 port map( A => n6725, Z => n13322);
   U121 : BUF_X1 port map( A => n6721, Z => n13332);
   U122 : BUF_X1 port map( A => n6721, Z => n13331);
   U123 : BUF_X1 port map( A => n6710, Z => n13349);
   U124 : BUF_X1 port map( A => n6704, Z => n13359);
   U125 : BUF_X1 port map( A => n6704, Z => n13358);
   U126 : BUF_X1 port map( A => n6701, Z => n13368);
   U127 : BUF_X1 port map( A => n6701, Z => n13367);
   U128 : BUF_X1 port map( A => n6695, Z => n13386);
   U129 : BUF_X1 port map( A => n6692, Z => n13395);
   U130 : BUF_X1 port map( A => n6689, Z => n13404);
   U131 : BUF_X1 port map( A => n6689, Z => n13403);
   U132 : BUF_X1 port map( A => n6686, Z => n13413);
   U133 : BUF_X1 port map( A => n6686, Z => n13412);
   U134 : BUF_X1 port map( A => n6681, Z => n13422);
   U135 : BUF_X1 port map( A => n6681, Z => n13421);
   U136 : BUF_X1 port map( A => n6677, Z => n13431);
   U137 : BUF_X1 port map( A => n6677, Z => n13430);
   U138 : BUF_X1 port map( A => n6674, Z => n13440);
   U139 : BUF_X1 port map( A => n6674, Z => n13439);
   U140 : BUF_X1 port map( A => n6671, Z => n13449);
   U141 : BUF_X1 port map( A => n6671, Z => n13448);
   U142 : BUF_X1 port map( A => n6665, Z => n13467);
   U143 : BUF_X1 port map( A => n6662, Z => n13476);
   U144 : BUF_X1 port map( A => n6659, Z => n13485);
   U145 : BUF_X1 port map( A => n6659, Z => n13484);
   U146 : BUF_X1 port map( A => n6656, Z => n13494);
   U147 : BUF_X1 port map( A => n6656, Z => n13493);
   U148 : BUF_X1 port map( A => n6653, Z => n13503);
   U149 : BUF_X1 port map( A => n6653, Z => n13502);
   U150 : BUF_X1 port map( A => n6650, Z => n13512);
   U151 : BUF_X1 port map( A => n6650, Z => n13511);
   U152 : BUF_X1 port map( A => n6647, Z => n13521);
   U153 : BUF_X1 port map( A => n6647, Z => n13520);
   U154 : BUF_X1 port map( A => n6644, Z => n13530);
   U155 : BUF_X1 port map( A => n6644, Z => n13529);
   U156 : BUF_X1 port map( A => n6638, Z => n13548);
   U157 : BUF_X1 port map( A => n6635, Z => n13557);
   U158 : BUF_X1 port map( A => n6630, Z => n13566);
   U159 : BUF_X1 port map( A => n6630, Z => n13565);
   U160 : BUF_X1 port map( A => n2679, Z => n14480);
   U161 : BUF_X1 port map( A => n2674, Z => n14489);
   U162 : BUF_X1 port map( A => n2704, Z => n14435);
   U163 : BUF_X1 port map( A => n2699, Z => n14443);
   U164 : BUF_X1 port map( A => n2679, Z => n14479);
   U165 : BUF_X1 port map( A => n2674, Z => n14488);
   U166 : BUF_X1 port map( A => n2694, Z => n14452);
   U167 : BUF_X1 port map( A => n2628, Z => n14690);
   U168 : BUF_X1 port map( A => n2628, Z => n14689);
   U169 : BUF_X1 port map( A => n6793, Z => n13260);
   U170 : BUF_X1 port map( A => n6793, Z => n13259);
   U171 : BUF_X1 port map( A => n6780, Z => n13269);
   U172 : BUF_X1 port map( A => n2726, Z => n14399);
   U173 : BUF_X1 port map( A => n2726, Z => n14398);
   U174 : BUF_X1 port map( A => n2704, Z => n14434);
   U175 : BUF_X1 port map( A => n6821, Z => n13233);
   U176 : BUF_X1 port map( A => n2699, Z => n14444);
   U177 : BUF_X1 port map( A => n2694, Z => n14453);
   U178 : BUF_X1 port map( A => n2689, Z => n14462);
   U179 : BUF_X1 port map( A => n2684, Z => n14471);
   U180 : BUF_X1 port map( A => n2669, Z => n14498);
   U181 : BUF_X1 port map( A => n2664, Z => n14507);
   U182 : BUF_X1 port map( A => n2689, Z => n14461);
   U183 : BUF_X1 port map( A => n2684, Z => n14470);
   U184 : BUF_X1 port map( A => n2669, Z => n14497);
   U185 : BUF_X1 port map( A => n2664, Z => n14506);
   U186 : BUF_X1 port map( A => n6808, Z => n13242);
   U187 : BUF_X1 port map( A => n6808, Z => n13241);
   U188 : BUF_X1 port map( A => n6801, Z => n13251);
   U189 : BUF_X1 port map( A => n6801, Z => n13250);
   U190 : BUF_X1 port map( A => n6780, Z => n13268);
   U191 : BUF_X1 port map( A => n6763, Z => n13278);
   U192 : BUF_X1 port map( A => n6763, Z => n13277);
   U193 : BUF_X1 port map( A => n2741, Z => n14372);
   U194 : BUF_X1 port map( A => n2741, Z => n14371);
   U195 : BUF_X1 port map( A => n2736, Z => n14381);
   U196 : BUF_X1 port map( A => n2736, Z => n14380);
   U197 : BUF_X1 port map( A => n2731, Z => n14390);
   U198 : BUF_X1 port map( A => n2731, Z => n14389);
   U199 : BUF_X1 port map( A => n2721, Z => n14408);
   U200 : BUF_X1 port map( A => n2721, Z => n14407);
   U201 : BUF_X1 port map( A => n2716, Z => n14417);
   U202 : BUF_X1 port map( A => n2716, Z => n14416);
   U203 : BUF_X1 port map( A => n2711, Z => n14426);
   U204 : BUF_X1 port map( A => n2711, Z => n14425);
   U205 : BUF_X1 port map( A => n2625, Z => n14706);
   U206 : BUF_X1 port map( A => n6748, Z => n13297);
   U207 : BUF_X1 port map( A => n6732, Z => n13315);
   U208 : BUF_X1 port map( A => n6716, Z => n13342);
   U209 : BUF_X1 port map( A => n6698, Z => n13378);
   U210 : BUF_X1 port map( A => n6668, Z => n13459);
   U211 : BUF_X1 port map( A => n6641, Z => n13540);
   U212 : BUF_X1 port map( A => n6753, Z => n13288);
   U213 : BUF_X1 port map( A => n6738, Z => n13306);
   U214 : BUF_X1 port map( A => n6725, Z => n13324);
   U215 : BUF_X1 port map( A => n6721, Z => n13333);
   U216 : BUF_X1 port map( A => n6710, Z => n13351);
   U217 : BUF_X1 port map( A => n6704, Z => n13360);
   U218 : BUF_X1 port map( A => n6701, Z => n13369);
   U219 : BUF_X1 port map( A => n6695, Z => n13387);
   U220 : BUF_X1 port map( A => n6692, Z => n13396);
   U221 : BUF_X1 port map( A => n6689, Z => n13405);
   U222 : BUF_X1 port map( A => n6686, Z => n13414);
   U223 : BUF_X1 port map( A => n6681, Z => n13423);
   U224 : BUF_X1 port map( A => n6677, Z => n13432);
   U225 : BUF_X1 port map( A => n6674, Z => n13441);
   U226 : BUF_X1 port map( A => n6671, Z => n13450);
   U227 : BUF_X1 port map( A => n6665, Z => n13468);
   U228 : BUF_X1 port map( A => n6662, Z => n13477);
   U229 : BUF_X1 port map( A => n6659, Z => n13486);
   U230 : BUF_X1 port map( A => n6656, Z => n13495);
   U231 : BUF_X1 port map( A => n6653, Z => n13504);
   U232 : BUF_X1 port map( A => n6650, Z => n13513);
   U233 : BUF_X1 port map( A => n6647, Z => n13522);
   U234 : BUF_X1 port map( A => n6644, Z => n13531);
   U235 : BUF_X1 port map( A => n6638, Z => n13549);
   U236 : BUF_X1 port map( A => n6635, Z => n13558);
   U237 : BUF_X1 port map( A => n6630, Z => n13567);
   U238 : BUF_X1 port map( A => n6821, Z => n13234);
   U239 : BUF_X1 port map( A => n2704, Z => n14436);
   U240 : BUF_X1 port map( A => n2694, Z => n14454);
   U241 : BUF_X1 port map( A => n2679, Z => n14481);
   U242 : BUF_X1 port map( A => n2674, Z => n14490);
   U243 : BUF_X1 port map( A => n2726, Z => n14400);
   U244 : BUF_X1 port map( A => n2628, Z => n14691);
   U245 : BUF_X1 port map( A => n6793, Z => n13261);
   U246 : BUF_X1 port map( A => n2699, Z => n14445);
   U247 : BUF_X1 port map( A => n2689, Z => n14463);
   U248 : BUF_X1 port map( A => n2684, Z => n14472);
   U249 : BUF_X1 port map( A => n2669, Z => n14499);
   U250 : BUF_X1 port map( A => n2664, Z => n14508);
   U251 : BUF_X1 port map( A => n2741, Z => n14373);
   U252 : BUF_X1 port map( A => n2736, Z => n14382);
   U253 : BUF_X1 port map( A => n2731, Z => n14391);
   U254 : BUF_X1 port map( A => n2721, Z => n14409);
   U255 : BUF_X1 port map( A => n2716, Z => n14418);
   U256 : BUF_X1 port map( A => n2711, Z => n14427);
   U257 : BUF_X1 port map( A => n6808, Z => n13243);
   U258 : BUF_X1 port map( A => n6801, Z => n13252);
   U259 : BUF_X1 port map( A => n6780, Z => n13270);
   U260 : BUF_X1 port map( A => n6763, Z => n13279);
   U261 : INV_X1 port map( A => n14965, ZN => n14943);
   U262 : INV_X1 port map( A => n14965, ZN => n14944);
   U263 : INV_X1 port map( A => n14965, ZN => n14945);
   U264 : INV_X1 port map( A => n14965, ZN => n14946);
   U265 : INV_X1 port map( A => n13871, ZN => n13870);
   U266 : INV_X1 port map( A => n14149, ZN => n14148);
   U267 : INV_X1 port map( A => n14964, ZN => n14942);
   U268 : INV_X1 port map( A => n13220, ZN => n13868);
   U269 : INV_X1 port map( A => n13220, ZN => n13869);
   U270 : INV_X1 port map( A => n14147, ZN => n14146);
   U271 : INV_X1 port map( A => n13221, ZN => n14354);
   U272 : INV_X1 port map( A => n13221, ZN => n14355);
   U273 : BUF_X1 port map( A => n2868, Z => n14110);
   U274 : BUF_X1 port map( A => n2874, Z => n14095);
   U275 : BUF_X1 port map( A => n2868, Z => n14109);
   U276 : BUF_X1 port map( A => n2874, Z => n14094);
   U277 : BUF_X1 port map( A => n4049, Z => n13905);
   U278 : BUF_X1 port map( A => n2559, Z => n14726);
   U279 : BUF_X1 port map( A => n2556, Z => n14732);
   U280 : BUF_X1 port map( A => n2559, Z => n14725);
   U281 : BUF_X1 port map( A => n2556, Z => n14731);
   U282 : BUF_X1 port map( A => n4049, Z => n13906);
   U283 : BUF_X1 port map( A => n2743, Z => n14366);
   U284 : BUF_X1 port map( A => n2705, Z => n14431);
   U285 : BUF_X1 port map( A => n2629, Z => n14686);
   U286 : BUF_X1 port map( A => n2622, Z => n14716);
   U287 : BUF_X1 port map( A => n2559, Z => n14727);
   U288 : BUF_X1 port map( A => n2680, Z => n14476);
   U289 : BUF_X1 port map( A => n2675, Z => n14485);
   U290 : BUF_X1 port map( A => n2727, Z => n14395);
   U291 : BUF_X1 port map( A => n2622, Z => n14717);
   U292 : BUF_X1 port map( A => n2706, Z => n14430);
   U293 : BUF_X1 port map( A => n2768, Z => n14311);
   U294 : BUF_X1 port map( A => n2728, Z => n14394);
   U295 : BUF_X1 port map( A => n2776, Z => n14289);
   U296 : BUF_X1 port map( A => n2772, Z => n14300);
   U297 : BUF_X1 port map( A => n2764, Z => n14320);
   U298 : BUF_X1 port map( A => n2760, Z => n14329);
   U299 : BUF_X1 port map( A => n2756, Z => n14338);
   U300 : BUF_X1 port map( A => n2752, Z => n14347);
   U301 : BUF_X1 port map( A => n2747, Z => n14358);
   U302 : BUF_X1 port map( A => n2738, Z => n14376);
   U303 : BUF_X1 port map( A => n2733, Z => n14385);
   U304 : BUF_X1 port map( A => n2723, Z => n14403);
   U305 : BUF_X1 port map( A => n2718, Z => n14412);
   U306 : BUF_X1 port map( A => n2713, Z => n14421);
   U307 : BUF_X1 port map( A => n2705, Z => n14432);
   U308 : BUF_X1 port map( A => n2695, Z => n14450);
   U309 : BUF_X1 port map( A => n2680, Z => n14477);
   U310 : BUF_X1 port map( A => n2675, Z => n14486);
   U311 : BUF_X1 port map( A => n2727, Z => n14396);
   U312 : BUF_X1 port map( A => n2629, Z => n14687);
   U313 : INV_X1 port map( A => n14286, ZN => n14276);
   U314 : INV_X1 port map( A => n14286, ZN => n14277);
   U315 : BUF_X1 port map( A => n2742, Z => n14369);
   U316 : BUF_X1 port map( A => n2742, Z => n14368);
   U317 : BUF_X1 port map( A => n2690, Z => n14459);
   U318 : BUF_X1 port map( A => n2690, Z => n14458);
   U319 : BUF_X1 port map( A => n2722, Z => n14405);
   U320 : BUF_X1 port map( A => n2722, Z => n14404);
   U321 : BUF_X1 port map( A => n2700, Z => n14440);
   U322 : BUF_X1 port map( A => n2685, Z => n14468);
   U323 : BUF_X1 port map( A => n2685, Z => n14467);
   U324 : BUF_X1 port map( A => n2670, Z => n14495);
   U325 : BUF_X1 port map( A => n2670, Z => n14494);
   U326 : BUF_X1 port map( A => n2665, Z => n14504);
   U327 : BUF_X1 port map( A => n2665, Z => n14503);
   U328 : BUF_X1 port map( A => n2737, Z => n14378);
   U329 : BUF_X1 port map( A => n2737, Z => n14377);
   U330 : BUF_X1 port map( A => n2732, Z => n14387);
   U331 : BUF_X1 port map( A => n2732, Z => n14386);
   U332 : BUF_X1 port map( A => n2717, Z => n14414);
   U333 : BUF_X1 port map( A => n2717, Z => n14413);
   U334 : BUF_X1 port map( A => n2712, Z => n14423);
   U335 : BUF_X1 port map( A => n2712, Z => n14422);
   U336 : BUF_X1 port map( A => n2867, Z => n14113);
   U337 : BUF_X1 port map( A => n2873, Z => n14098);
   U338 : BUF_X1 port map( A => n2867, Z => n14112);
   U339 : BUF_X1 port map( A => n2873, Z => n14097);
   U340 : BUF_X1 port map( A => n2542, Z => n14737);
   U341 : BUF_X1 port map( A => n2565, Z => n14722);
   U342 : BUF_X1 port map( A => n2542, Z => n14738);
   U343 : BUF_X1 port map( A => n2565, Z => n14723);
   U344 : BUF_X1 port map( A => n2700, Z => n14441);
   U345 : BUF_X1 port map( A => n2695, Z => n14449);
   U346 : BUF_X1 port map( A => n2558, Z => n14728);
   U347 : BUF_X1 port map( A => n2566, Z => n14719);
   U348 : BUF_X1 port map( A => n2566, Z => n14720);
   U349 : BUF_X1 port map( A => n2541, Z => n14740);
   U350 : BUF_X1 port map( A => n2541, Z => n14741);
   U351 : BUF_X1 port map( A => n5372, Z => n13673);
   U352 : BUF_X1 port map( A => n5372, Z => n13674);
   U353 : BUF_X1 port map( A => n2555, Z => n14735);
   U354 : BUF_X1 port map( A => n2558, Z => n14729);
   U355 : BUF_X1 port map( A => n2555, Z => n14734);
   U356 : BUF_X1 port map( A => n2743, Z => n14365);
   U357 : BUF_X1 port map( A => n2768, Z => n14309);
   U358 : BUF_X1 port map( A => n2728, Z => n14392);
   U359 : BUF_X1 port map( A => n2706, Z => n14428);
   U360 : BUF_X1 port map( A => n2756, Z => n14336);
   U361 : BUF_X1 port map( A => n2752, Z => n14345);
   U362 : BUF_X1 port map( A => n2738, Z => n14374);
   U363 : BUF_X1 port map( A => n2776, Z => n14287);
   U364 : BUF_X1 port map( A => n2772, Z => n14298);
   U365 : BUF_X1 port map( A => n2764, Z => n14318);
   U366 : BUF_X1 port map( A => n2760, Z => n14327);
   U367 : BUF_X1 port map( A => n2747, Z => n14356);
   U368 : BUF_X1 port map( A => n2733, Z => n14383);
   U369 : BUF_X1 port map( A => n2723, Z => n14401);
   U370 : BUF_X1 port map( A => n2718, Z => n14410);
   U371 : BUF_X1 port map( A => n2713, Z => n14419);
   U372 : BUF_X1 port map( A => n2706, Z => n14429);
   U373 : BUF_X1 port map( A => n2768, Z => n14310);
   U374 : BUF_X1 port map( A => n2728, Z => n14393);
   U375 : BUF_X1 port map( A => n2756, Z => n14337);
   U376 : BUF_X1 port map( A => n2752, Z => n14346);
   U377 : BUF_X1 port map( A => n2738, Z => n14375);
   U378 : BUF_X1 port map( A => n2776, Z => n14288);
   U379 : BUF_X1 port map( A => n2772, Z => n14299);
   U380 : BUF_X1 port map( A => n2764, Z => n14319);
   U381 : BUF_X1 port map( A => n2760, Z => n14328);
   U382 : BUF_X1 port map( A => n2747, Z => n14357);
   U383 : BUF_X1 port map( A => n2733, Z => n14384);
   U384 : BUF_X1 port map( A => n2723, Z => n14402);
   U385 : BUF_X1 port map( A => n2718, Z => n14411);
   U386 : BUF_X1 port map( A => n2713, Z => n14420);
   U387 : BUF_X1 port map( A => n2558, Z => n14730);
   U388 : BUF_X1 port map( A => n6823, Z => n13229);
   U389 : BUF_X1 port map( A => n6796, Z => n13257);
   U390 : BUF_X1 port map( A => n6796, Z => n13256);
   U391 : BUF_X1 port map( A => n6783, Z => n13266);
   U392 : BUF_X1 port map( A => n6823, Z => n13230);
   U393 : BUF_X1 port map( A => n6811, Z => n13239);
   U394 : BUF_X1 port map( A => n6811, Z => n13238);
   U395 : BUF_X1 port map( A => n6802, Z => n13248);
   U396 : BUF_X1 port map( A => n6802, Z => n13247);
   U397 : BUF_X1 port map( A => n6783, Z => n13265);
   U398 : BUF_X1 port map( A => n6769, Z => n13275);
   U399 : BUF_X1 port map( A => n6769, Z => n13274);
   U400 : BUF_X1 port map( A => n2742, Z => n14370);
   U401 : BUF_X1 port map( A => n6757, Z => n13284);
   U402 : BUF_X1 port map( A => n6757, Z => n13283);
   U403 : BUF_X1 port map( A => n6678, Z => n13428);
   U404 : BUF_X1 port map( A => n6678, Z => n13427);
   U405 : BUF_X1 port map( A => n2690, Z => n14460);
   U406 : BUF_X1 port map( A => n2722, Z => n14406);
   U407 : BUF_X1 port map( A => n6749, Z => n13293);
   U408 : BUF_X1 port map( A => n6749, Z => n13292);
   U409 : BUF_X1 port map( A => n6739, Z => n13301);
   U410 : BUF_X1 port map( A => n6733, Z => n13310);
   U411 : BUF_X1 port map( A => n6717, Z => n13338);
   U412 : BUF_X1 port map( A => n6717, Z => n13337);
   U413 : BUF_X1 port map( A => n6711, Z => n13347);
   U414 : BUF_X1 port map( A => n6699, Z => n13374);
   U415 : BUF_X1 port map( A => n6699, Z => n13373);
   U416 : BUF_X1 port map( A => n6696, Z => n13382);
   U417 : BUF_X1 port map( A => n6693, Z => n13391);
   U418 : BUF_X1 port map( A => n6669, Z => n13455);
   U419 : BUF_X1 port map( A => n6669, Z => n13454);
   U420 : BUF_X1 port map( A => n6666, Z => n13463);
   U421 : BUF_X1 port map( A => n6663, Z => n13472);
   U422 : BUF_X1 port map( A => n6642, Z => n13536);
   U423 : BUF_X1 port map( A => n6642, Z => n13535);
   U424 : BUF_X1 port map( A => n6639, Z => n13544);
   U425 : BUF_X1 port map( A => n6636, Z => n13553);
   U426 : BUF_X1 port map( A => n6739, Z => n13302);
   U427 : BUF_X1 port map( A => n6733, Z => n13311);
   U428 : BUF_X1 port map( A => n6729, Z => n13320);
   U429 : BUF_X1 port map( A => n6729, Z => n13319);
   U430 : BUF_X1 port map( A => n6722, Z => n13329);
   U431 : BUF_X1 port map( A => n6722, Z => n13328);
   U432 : BUF_X1 port map( A => n6711, Z => n13346);
   U433 : BUF_X1 port map( A => n6705, Z => n13356);
   U434 : BUF_X1 port map( A => n6705, Z => n13355);
   U435 : BUF_X1 port map( A => n6702, Z => n13365);
   U436 : BUF_X1 port map( A => n6702, Z => n13364);
   U437 : BUF_X1 port map( A => n6696, Z => n13383);
   U438 : BUF_X1 port map( A => n6693, Z => n13392);
   U439 : BUF_X1 port map( A => n6690, Z => n13401);
   U440 : BUF_X1 port map( A => n6690, Z => n13400);
   U441 : BUF_X1 port map( A => n6687, Z => n13410);
   U442 : BUF_X1 port map( A => n6687, Z => n13409);
   U443 : BUF_X1 port map( A => n6682, Z => n13419);
   U444 : BUF_X1 port map( A => n6682, Z => n13418);
   U445 : BUF_X1 port map( A => n6675, Z => n13437);
   U446 : BUF_X1 port map( A => n6675, Z => n13436);
   U447 : BUF_X1 port map( A => n6672, Z => n13446);
   U448 : BUF_X1 port map( A => n6672, Z => n13445);
   U449 : BUF_X1 port map( A => n6666, Z => n13464);
   U450 : BUF_X1 port map( A => n6663, Z => n13473);
   U451 : BUF_X1 port map( A => n6660, Z => n13482);
   U452 : BUF_X1 port map( A => n6660, Z => n13481);
   U453 : BUF_X1 port map( A => n6657, Z => n13491);
   U454 : BUF_X1 port map( A => n6657, Z => n13490);
   U455 : BUF_X1 port map( A => n6654, Z => n13500);
   U456 : BUF_X1 port map( A => n6654, Z => n13499);
   U457 : BUF_X1 port map( A => n6651, Z => n13509);
   U458 : BUF_X1 port map( A => n6651, Z => n13508);
   U459 : BUF_X1 port map( A => n6648, Z => n13518);
   U460 : BUF_X1 port map( A => n6648, Z => n13517);
   U461 : BUF_X1 port map( A => n6645, Z => n13527);
   U462 : BUF_X1 port map( A => n6645, Z => n13526);
   U463 : BUF_X1 port map( A => n6639, Z => n13545);
   U464 : BUF_X1 port map( A => n6636, Z => n13554);
   U465 : BUF_X1 port map( A => n6631, Z => n13563);
   U466 : BUF_X1 port map( A => n6631, Z => n13562);
   U467 : BUF_X1 port map( A => n2762, Z => n14325);
   U468 : BUF_X1 port map( A => n2762, Z => n14324);
   U469 : BUF_X1 port map( A => n6612, Z => n13620);
   U470 : BUF_X1 port map( A => n6612, Z => n13619);
   U471 : BUF_X1 port map( A => n6609, Z => n13628);
   U472 : BUF_X1 port map( A => n2750, Z => n14352);
   U473 : BUF_X1 port map( A => n2750, Z => n14351);
   U474 : BUF_X1 port map( A => n6627, Z => n13575);
   U475 : BUF_X1 port map( A => n6627, Z => n13574);
   U476 : BUF_X1 port map( A => n6624, Z => n13584);
   U477 : BUF_X1 port map( A => n6624, Z => n13583);
   U478 : BUF_X1 port map( A => n6621, Z => n13593);
   U479 : BUF_X1 port map( A => n6621, Z => n13592);
   U480 : BUF_X1 port map( A => n6618, Z => n13602);
   U481 : BUF_X1 port map( A => n6618, Z => n13601);
   U482 : BUF_X1 port map( A => n6615, Z => n13611);
   U483 : BUF_X1 port map( A => n6615, Z => n13610);
   U484 : BUF_X1 port map( A => n6609, Z => n13629);
   U485 : BUF_X1 port map( A => n2758, Z => n14334);
   U486 : BUF_X1 port map( A => n2758, Z => n14333);
   U487 : BUF_X1 port map( A => n2754, Z => n14343);
   U488 : BUF_X1 port map( A => n2754, Z => n14342);
   U489 : BUF_X1 port map( A => n2766, Z => n14316);
   U490 : BUF_X1 port map( A => n2766, Z => n14315);
   U491 : BUF_X1 port map( A => n2774, Z => n14294);
   U492 : BUF_X1 port map( A => n2774, Z => n14293);
   U493 : BUF_X1 port map( A => n2770, Z => n14305);
   U494 : BUF_X1 port map( A => n2770, Z => n14304);
   U495 : BUF_X1 port map( A => n2745, Z => n14363);
   U496 : BUF_X1 port map( A => n2745, Z => n14362);
   U497 : BUF_X1 port map( A => n6605, Z => n13635);
   U498 : BUF_X1 port map( A => n6605, Z => n13634);
   U499 : BUF_X1 port map( A => n2743, Z => n14367);
   U500 : BUF_X1 port map( A => n5277, Z => n13862);
   U501 : BUF_X1 port map( A => n3956, Z => n14082);
   U502 : BUF_X1 port map( A => n3956, Z => n14083);
   U503 : BUF_X1 port map( A => n5277, Z => n13863);
   U504 : BUF_X1 port map( A => n2670, Z => n14496);
   U505 : BUF_X1 port map( A => n2665, Z => n14505);
   U506 : BUF_X1 port map( A => n2737, Z => n14379);
   U507 : BUF_X1 port map( A => n2732, Z => n14388);
   U508 : BUF_X1 port map( A => n2717, Z => n14415);
   U509 : BUF_X1 port map( A => n2712, Z => n14424);
   U510 : BUF_X1 port map( A => n2685, Z => n14469);
   U511 : BUF_X1 port map( A => n2556, Z => n14733);
   U512 : BUF_X1 port map( A => n2867, Z => n14114);
   U513 : BUF_X1 port map( A => n2873, Z => n14099);
   U514 : BUF_X1 port map( A => n2868, Z => n14111);
   U515 : BUF_X1 port map( A => n2874, Z => n14096);
   U516 : BUF_X1 port map( A => n5372, Z => n13675);
   U517 : BUF_X1 port map( A => n6823, Z => n13231);
   U518 : BUF_X1 port map( A => n6796, Z => n13258);
   U519 : BUF_X1 port map( A => n6811, Z => n13240);
   U520 : BUF_X1 port map( A => n6802, Z => n13249);
   U521 : BUF_X1 port map( A => n6783, Z => n13267);
   U522 : BUF_X1 port map( A => n6769, Z => n13276);
   U523 : BUF_X1 port map( A => n6757, Z => n13285);
   U524 : BUF_X1 port map( A => n6678, Z => n13429);
   U525 : BUF_X1 port map( A => n2700, Z => n14442);
   U526 : BUF_X1 port map( A => n6749, Z => n13294);
   U527 : BUF_X1 port map( A => n6733, Z => n13312);
   U528 : BUF_X1 port map( A => n6717, Z => n13339);
   U529 : BUF_X1 port map( A => n6699, Z => n13375);
   U530 : BUF_X1 port map( A => n6669, Z => n13456);
   U531 : BUF_X1 port map( A => n6642, Z => n13537);
   U532 : BUF_X1 port map( A => n6739, Z => n13303);
   U533 : BUF_X1 port map( A => n6729, Z => n13321);
   U534 : BUF_X1 port map( A => n6722, Z => n13330);
   U535 : BUF_X1 port map( A => n6711, Z => n13348);
   U536 : BUF_X1 port map( A => n6705, Z => n13357);
   U537 : BUF_X1 port map( A => n6702, Z => n13366);
   U538 : BUF_X1 port map( A => n6696, Z => n13384);
   U539 : BUF_X1 port map( A => n6693, Z => n13393);
   U540 : BUF_X1 port map( A => n6690, Z => n13402);
   U541 : BUF_X1 port map( A => n6687, Z => n13411);
   U542 : BUF_X1 port map( A => n6682, Z => n13420);
   U543 : BUF_X1 port map( A => n6675, Z => n13438);
   U544 : BUF_X1 port map( A => n6672, Z => n13447);
   U545 : BUF_X1 port map( A => n6666, Z => n13465);
   U546 : BUF_X1 port map( A => n6663, Z => n13474);
   U547 : BUF_X1 port map( A => n6660, Z => n13483);
   U548 : BUF_X1 port map( A => n6657, Z => n13492);
   U549 : BUF_X1 port map( A => n6654, Z => n13501);
   U550 : BUF_X1 port map( A => n6651, Z => n13510);
   U551 : BUF_X1 port map( A => n6648, Z => n13519);
   U552 : BUF_X1 port map( A => n6645, Z => n13528);
   U553 : BUF_X1 port map( A => n6639, Z => n13546);
   U554 : BUF_X1 port map( A => n6636, Z => n13555);
   U555 : BUF_X1 port map( A => n6631, Z => n13564);
   U556 : INV_X1 port map( A => n2708, ZN => n2581);
   U557 : BUF_X1 port map( A => n2762, Z => n14326);
   U558 : BUF_X1 port map( A => n6612, Z => n13621);
   U559 : BUF_X1 port map( A => n2750, Z => n14353);
   U560 : BUF_X1 port map( A => n2758, Z => n14335);
   U561 : BUF_X1 port map( A => n6627, Z => n13576);
   U562 : BUF_X1 port map( A => n6624, Z => n13585);
   U563 : BUF_X1 port map( A => n6621, Z => n13594);
   U564 : BUF_X1 port map( A => n6618, Z => n13603);
   U565 : BUF_X1 port map( A => n6615, Z => n13612);
   U566 : BUF_X1 port map( A => n6609, Z => n13630);
   U567 : BUF_X1 port map( A => n2754, Z => n14344);
   U568 : BUF_X1 port map( A => n2766, Z => n14317);
   U569 : BUF_X1 port map( A => n2774, Z => n14295);
   U570 : BUF_X1 port map( A => n2770, Z => n14306);
   U571 : BUF_X1 port map( A => n2745, Z => n14364);
   U572 : BUF_X1 port map( A => n6605, Z => n13636);
   U573 : BUF_X1 port map( A => n3956, Z => n14084);
   U574 : BUF_X1 port map( A => n5277, Z => n13864);
   U575 : BUF_X1 port map( A => n2555, Z => n14736);
   U576 : BUF_X1 port map( A => n2695, Z => n14451);
   U577 : BUF_X1 port map( A => n2542, Z => n14739);
   U578 : BUF_X1 port map( A => n2622, Z => n14718);
   U579 : BUF_X1 port map( A => n2680, Z => n14478);
   U580 : BUF_X1 port map( A => n2675, Z => n14487);
   U581 : BUF_X1 port map( A => n2705, Z => n14433);
   U582 : BUF_X1 port map( A => n2629, Z => n14688);
   U583 : BUF_X1 port map( A => n2727, Z => n14397);
   U584 : BUF_X1 port map( A => n2541, Z => n14742);
   U585 : BUF_X1 port map( A => n4049, Z => n13907);
   U586 : BUF_X1 port map( A => n2565, Z => n14724);
   U587 : BUF_X1 port map( A => n2566, Z => n14721);
   U588 : INV_X1 port map( A => n13223, ZN => n14115);
   U589 : INV_X1 port map( A => n13222, ZN => n14296);
   U590 : INV_X1 port map( A => n13224, ZN => n14308);
   U591 : OAI221_X1 port map( B1 => n2660, B2 => n2739, C1 => n14964, C2 => 
                           n14709, A => n14743, ZN => n2622);
   U592 : OAI221_X1 port map( B1 => n2660, B2 => n2719, C1 => n14963, C2 => 
                           n13253, A => n14743, ZN => n6796);
   U593 : OAI221_X1 port map( B1 => n2660, B2 => n2734, C1 => n14964, C2 => 
                           n13226, A => n14743, ZN => n6823);
   U594 : OAI221_X1 port map( B1 => n2660, B2 => n2729, C1 => n14964, C2 => 
                           n13235, A => n14743, ZN => n6811);
   U595 : OAI221_X1 port map( B1 => n2660, B2 => n2724, C1 => n14964, C2 => 
                           n13244, A => n14743, ZN => n6802);
   U596 : OAI221_X1 port map( B1 => n2660, B2 => n2714, C1 => n14963, C2 => 
                           n13262, A => n14743, ZN => n6783);
   U597 : OAI221_X1 port map( B1 => n2660, B2 => n2708, C1 => n14963, C2 => 
                           n13271, A => n14743, ZN => n6769);
   U598 : INV_X1 port map( A => n13225, ZN => n14117);
   U599 : OAI221_X1 port map( B1 => n2702, B2 => n6684, C1 => n14963, C2 => 
                           n13280, A => n14743, ZN => n6757);
   U600 : OAI221_X1 port map( B1 => n2702, B2 => n6633, C1 => n14962, C2 => 
                           n13424, A => n14744, ZN => n6678);
   U601 : OAI221_X1 port map( B1 => n2661, B2 => n2707, C1 => n14962, C2 => 
                           n14365, A => n14747, ZN => n2742);
   U602 : OAI221_X1 port map( B1 => n14949, B2 => n14428, C1 => n2707, C2 => 
                           n2708, A => n14748, ZN => n2705);
   U603 : OAI221_X1 port map( B1 => n14947, B2 => n14473, C1 => n2660, C2 => 
                           n2682, A => n14748, ZN => n2680);
   U604 : OAI221_X1 port map( B1 => n14947, B2 => n14482, C1 => n2660, C2 => 
                           n2677, A => n14748, ZN => n2675);
   U605 : OAI221_X1 port map( B1 => n14950, B2 => n14392, C1 => n2707, C2 => 
                           n2729, A => n14747, ZN => n2727);
   U606 : OAI221_X1 port map( B1 => n14956, B2 => n14685, C1 => n2660, C2 => 
                           n2661, A => n14748, ZN => n2629);
   U607 : OAI221_X1 port map( B1 => n14962, B2 => n13289, C1 => n2697, C2 => 
                           n6684, A => n14743, ZN => n6749);
   U608 : OAI221_X1 port map( B1 => n14961, B2 => n13334, C1 => n2672, C2 => 
                           n6684, A => n14744, ZN => n6717);
   U609 : OAI221_X1 port map( B1 => n14960, B2 => n13370, C1 => n2734, C2 => 
                           n6684, A => n14744, ZN => n6699);
   U610 : OAI221_X1 port map( B1 => n14957, B2 => n13451, C1 => n2687, C2 => 
                           n6633, A => n14745, ZN => n6669);
   U611 : OAI221_X1 port map( B1 => n14955, B2 => n13532, C1 => n2724, C2 => 
                           n6633, A => n14745, ZN => n6642);
   U612 : OAI221_X1 port map( B1 => n14948, B2 => n14446, C1 => n2660, C2 => 
                           n2697, A => n14748, ZN => n2695);
   U613 : OAI221_X1 port map( B1 => n14961, B2 => n13307, C1 => n2687, C2 => 
                           n6684, A => n14743, ZN => n6733);
   U614 : OAI221_X1 port map( B1 => n14948, B2 => n14437, C1 => n2660, C2 => 
                           n2702, A => n14748, ZN => n2700);
   U615 : OAI221_X1 port map( B1 => n14948, B2 => n14455, C1 => n2660, C2 => 
                           n2692, A => n14748, ZN => n2690);
   U616 : OAI221_X1 port map( B1 => n14948, B2 => n14464, C1 => n2660, C2 => 
                           n2687, A => n14748, ZN => n2685);
   U617 : OAI221_X1 port map( B1 => n14947, B2 => n14491, C1 => n2660, C2 => 
                           n2672, A => n14748, ZN => n2670);
   U618 : OAI221_X1 port map( B1 => n14947, B2 => n14500, C1 => n2660, C2 => 
                           n2667, A => n14748, ZN => n2665);
   U619 : OAI221_X1 port map( B1 => n14950, B2 => n14374, C1 => n2739, C2 => 
                           n2707, A => n14747, ZN => n2737);
   U620 : OAI221_X1 port map( B1 => n14950, B2 => n14383, C1 => n2707, C2 => 
                           n2734, A => n14747, ZN => n2732);
   U621 : OAI221_X1 port map( B1 => n14949, B2 => n14401, C1 => n2707, C2 => 
                           n2724, A => n14747, ZN => n2722);
   U622 : OAI221_X1 port map( B1 => n14949, B2 => n14410, C1 => n2707, C2 => 
                           n2719, A => n14748, ZN => n2717);
   U623 : OAI221_X1 port map( B1 => n14949, B2 => n14419, C1 => n2707, C2 => 
                           n2714, A => n14748, ZN => n2712);
   U624 : OAI221_X1 port map( B1 => n14960, B2 => n13298, C1 => n2692, C2 => 
                           n6684, A => n14743, ZN => n6739);
   U625 : OAI221_X1 port map( B1 => n14961, B2 => n13316, C1 => n2682, C2 => 
                           n6684, A => n14743, ZN => n6729);
   U626 : OAI221_X1 port map( B1 => n14960, B2 => n13325, C1 => n2677, C2 => 
                           n6684, A => n14744, ZN => n6722);
   U627 : OAI221_X1 port map( B1 => n14961, B2 => n13343, C1 => n2667, C2 => 
                           n6684, A => n14744, ZN => n6711);
   U628 : OAI221_X1 port map( B1 => n14958, B2 => n13352, C1 => n2661, C2 => 
                           n6684, A => n14744, ZN => n6705);
   U629 : OAI221_X1 port map( B1 => n14960, B2 => n13361, C1 => n2739, C2 => 
                           n6684, A => n14744, ZN => n6702);
   U630 : OAI221_X1 port map( B1 => n14959, B2 => n13379, C1 => n2729, C2 => 
                           n6684, A => n14744, ZN => n6696);
   U631 : OAI221_X1 port map( B1 => n14959, B2 => n13388, C1 => n2724, C2 => 
                           n6684, A => n14744, ZN => n6693);
   U632 : OAI221_X1 port map( B1 => n14959, B2 => n13397, C1 => n2719, C2 => 
                           n6684, A => n14744, ZN => n6690);
   U633 : OAI221_X1 port map( B1 => n14958, B2 => n13406, C1 => n2714, C2 => 
                           n6684, A => n14744, ZN => n6687);
   U634 : OAI221_X1 port map( B1 => n14959, B2 => n13415, C1 => n2708, C2 => 
                           n6684, A => n14744, ZN => n6682);
   U635 : OAI221_X1 port map( B1 => n14958, B2 => n13433, C1 => n2697, C2 => 
                           n6633, A => n14745, ZN => n6675);
   U636 : OAI221_X1 port map( B1 => n14958, B2 => n13442, C1 => n2692, C2 => 
                           n6633, A => n14745, ZN => n6672);
   U637 : OAI221_X1 port map( B1 => n14957, B2 => n13460, C1 => n2682, C2 => 
                           n6633, A => n14745, ZN => n6666);
   U638 : OAI221_X1 port map( B1 => n14957, B2 => n13469, C1 => n2677, C2 => 
                           n6633, A => n14745, ZN => n6663);
   U639 : OAI221_X1 port map( B1 => n14957, B2 => n13478, C1 => n2672, C2 => 
                           n6633, A => n14745, ZN => n6660);
   U640 : OAI221_X1 port map( B1 => n14956, B2 => n13487, C1 => n2667, C2 => 
                           n6633, A => n14745, ZN => n6657);
   U641 : OAI221_X1 port map( B1 => n14956, B2 => n13496, C1 => n2661, C2 => 
                           n6633, A => n14745, ZN => n6654);
   U642 : OAI221_X1 port map( B1 => n14956, B2 => n13505, C1 => n2739, C2 => 
                           n6633, A => n14745, ZN => n6651);
   U643 : OAI221_X1 port map( B1 => n14955, B2 => n13514, C1 => n2734, C2 => 
                           n6633, A => n14745, ZN => n6648);
   U644 : OAI221_X1 port map( B1 => n14955, B2 => n13523, C1 => n2729, C2 => 
                           n6633, A => n14745, ZN => n6645);
   U645 : OAI221_X1 port map( B1 => n14955, B2 => n13541, C1 => n2719, C2 => 
                           n6633, A => n14746, ZN => n6639);
   U646 : OAI221_X1 port map( B1 => n14954, B2 => n13550, C1 => n2714, C2 => 
                           n6633, A => n14746, ZN => n6636);
   U647 : OAI221_X1 port map( B1 => n14954, B2 => n13559, C1 => n2708, C2 => 
                           n6633, A => n14746, ZN => n6631);
   U648 : INV_X1 port map( A => n6684, ZN => n2525);
   U649 : INV_X1 port map( A => n6633, ZN => n2526);
   U650 : INV_X1 port map( A => n2660, ZN => n2524);
   U651 : INV_X1 port map( A => n13225, ZN => n14118);
   U652 : BUF_X1 port map( A => n2814, Z => n14213);
   U653 : INV_X1 port map( A => n2677, ZN => n2572);
   U654 : INV_X1 port map( A => n2682, ZN => n2576);
   U655 : BUF_X1 port map( A => n3993, Z => n14016);
   U656 : BUF_X1 port map( A => n4019, Z => n13962);
   U657 : BUF_X1 port map( A => n4030, Z => n13935);
   U658 : BUF_X1 port map( A => n4025, Z => n13947);
   U659 : BUF_X1 port map( A => n4054, Z => n13893);
   U660 : BUF_X1 port map( A => n4060, Z => n13878);
   U661 : INV_X1 port map( A => n2672, ZN => n2577);
   U662 : NOR2_X1 port map( A1 => n2708, A2 => n2563, ZN => n2867);
   U663 : NOR2_X1 port map( A1 => n2719, A2 => n2563, ZN => n2873);
   U664 : BUF_X1 port map( A => n2788, Z => n14267);
   U665 : BUF_X1 port map( A => n2794, Z => n14253);
   U666 : BUF_X1 port map( A => n2825, Z => n14187);
   U667 : BUF_X1 port map( A => n2820, Z => n14199);
   U668 : BUF_X1 port map( A => n2831, Z => n14172);
   U669 : BUF_X1 port map( A => n2855, Z => n14126);
   U670 : BUF_X1 port map( A => n2788, Z => n14268);
   U671 : BUF_X1 port map( A => n2794, Z => n14252);
   U672 : BUF_X1 port map( A => n2825, Z => n14186);
   U673 : BUF_X1 port map( A => n2820, Z => n14198);
   U674 : BUF_X1 port map( A => n2831, Z => n14171);
   U675 : BUF_X1 port map( A => n2855, Z => n14125);
   U676 : BUF_X1 port map( A => n3993, Z => n14017);
   U677 : BUF_X1 port map( A => n4019, Z => n13963);
   U678 : BUF_X1 port map( A => n4030, Z => n13936);
   U679 : BUF_X1 port map( A => n4025, Z => n13948);
   U680 : BUF_X1 port map( A => n4054, Z => n13894);
   U681 : BUF_X1 port map( A => n4060, Z => n13879);
   U682 : BUF_X1 port map( A => n2814, Z => n14214);
   U683 : NAND2_X1 port map( A1 => n6576, A2 => n6775, ZN => n2708);
   U684 : BUF_X1 port map( A => n2833, Z => n14169);
   U685 : BUF_X1 port map( A => n2857, Z => n14123);
   U686 : BUF_X1 port map( A => n3997, Z => n14007);
   U687 : BUF_X1 port map( A => n4023, Z => n13953);
   U688 : BUF_X1 port map( A => n4034, Z => n13926);
   U689 : BUF_X1 port map( A => n4058, Z => n13884);
   U690 : BUF_X1 port map( A => n5278, Z => n13859);
   U691 : BUF_X1 port map( A => n5278, Z => n13860);
   U692 : BUF_X1 port map( A => n3957, Z => n14079);
   U693 : BUF_X1 port map( A => n3957, Z => n14080);
   U694 : BUF_X1 port map( A => n3997, Z => n14008);
   U695 : BUF_X1 port map( A => n4023, Z => n13954);
   U696 : BUF_X1 port map( A => n4034, Z => n13927);
   U697 : BUF_X1 port map( A => n4058, Z => n13885);
   U698 : BUF_X1 port map( A => n6797, Z => n13254);
   U699 : BUF_X1 port map( A => n6784, Z => n13263);
   U700 : BUF_X1 port map( A => n6825, Z => n13227);
   U701 : BUF_X1 port map( A => n6759, Z => n13281);
   U702 : BUF_X1 port map( A => n6679, Z => n13425);
   U703 : BUF_X1 port map( A => n6819, Z => n13236);
   U704 : BUF_X1 port map( A => n6807, Z => n13245);
   U705 : BUF_X1 port map( A => n6772, Z => n13272);
   U706 : BUF_X1 port map( A => n6629, Z => n13569);
   U707 : BUF_X1 port map( A => n5307, Z => n13805);
   U708 : BUF_X1 port map( A => n3986, Z => n14025);
   U709 : BUF_X1 port map( A => n3986, Z => n14026);
   U710 : BUF_X1 port map( A => n5307, Z => n13806);
   U711 : BUF_X1 port map( A => n5296, Z => n13832);
   U712 : BUF_X1 port map( A => n3975, Z => n14052);
   U713 : BUF_X1 port map( A => n4012, Z => n13971);
   U714 : BUF_X1 port map( A => n4001, Z => n13998);
   U715 : BUF_X1 port map( A => n3975, Z => n14053);
   U716 : BUF_X1 port map( A => n4001, Z => n13999);
   U717 : BUF_X1 port map( A => n4012, Z => n13972);
   U718 : BUF_X1 port map( A => n5322, Z => n13778);
   U719 : BUF_X1 port map( A => n5333, Z => n13751);
   U720 : BUF_X1 port map( A => n4062, Z => n13875);
   U721 : BUF_X1 port map( A => n4062, Z => n13876);
   U722 : BUF_X1 port map( A => n5296, Z => n13833);
   U723 : BUF_X1 port map( A => n5359, Z => n13697);
   U724 : BUF_X1 port map( A => n5322, Z => n13779);
   U725 : BUF_X1 port map( A => n5333, Z => n13752);
   U726 : BUF_X1 port map( A => n2876, Z => n14092);
   U727 : BUF_X1 port map( A => n2876, Z => n14091);
   U728 : BUF_X1 port map( A => n5359, Z => n13698);
   U729 : BUF_X1 port map( A => n5348, Z => n13724);
   U730 : BUF_X1 port map( A => n5385, Z => n13643);
   U731 : BUF_X1 port map( A => n4027, Z => n13944);
   U732 : BUF_X1 port map( A => n4027, Z => n13945);
   U733 : BUF_X1 port map( A => n5348, Z => n13725);
   U734 : BUF_X1 port map( A => n5385, Z => n13644);
   U735 : BUF_X1 port map( A => n2857, Z => n14122);
   U736 : BUF_X1 port map( A => n2833, Z => n14168);
   U737 : BUF_X1 port map( A => n2767, Z => n14312);
   U738 : BUF_X1 port map( A => n2852, Z => n14134);
   U739 : BUF_X1 port map( A => n3957, Z => n14076);
   U740 : BUF_X1 port map( A => n5278, Z => n13856);
   U741 : BUF_X1 port map( A => n3957, Z => n14077);
   U742 : BUF_X1 port map( A => n5278, Z => n13857);
   U743 : BUF_X1 port map( A => n2630, Z => n14683);
   U744 : BUF_X1 port map( A => n2630, Z => n14684);
   U745 : BUF_X1 port map( A => n2853, Z => n14131);
   U746 : BUF_X1 port map( A => n2853, Z => n14132);
   U747 : BUF_X1 port map( A => n2792, Z => n14259);
   U748 : BUF_X1 port map( A => n2818, Z => n14205);
   U749 : BUF_X1 port map( A => n2829, Z => n14178);
   U750 : BUF_X1 port map( A => n2792, Z => n14258);
   U751 : BUF_X1 port map( A => n2818, Z => n14204);
   U752 : BUF_X1 port map( A => n2829, Z => n14177);
   U753 : BUF_X1 port map( A => n3995, Z => n14013);
   U754 : BUF_X1 port map( A => n4032, Z => n13932);
   U755 : BUF_X1 port map( A => n4056, Z => n13890);
   U756 : BUF_X1 port map( A => n4021, Z => n13959);
   U757 : BUF_X1 port map( A => n6606, Z => n13633);
   U758 : BUF_X1 port map( A => n2681, Z => n14475);
   U759 : BUF_X1 port map( A => n2676, Z => n14484);
   U760 : BUF_X1 port map( A => n6751, Z => n13291);
   U761 : BUF_X1 port map( A => n6718, Z => n13336);
   U762 : BUF_X1 port map( A => n6700, Z => n13372);
   U763 : BUF_X1 port map( A => n6670, Z => n13453);
   U764 : BUF_X1 port map( A => n6643, Z => n13534);
   U765 : BUF_X1 port map( A => n6614, Z => n13615);
   U766 : BUF_X1 port map( A => n2696, Z => n14448);
   U767 : BUF_X1 port map( A => n6735, Z => n13309);
   U768 : BUF_X1 port map( A => n2701, Z => n14439);
   U769 : BUF_X1 port map( A => n2691, Z => n14457);
   U770 : BUF_X1 port map( A => n2686, Z => n14466);
   U771 : BUF_X1 port map( A => n2671, Z => n14493);
   U772 : BUF_X1 port map( A => n2666, Z => n14502);
   U773 : BUF_X1 port map( A => n6747, Z => n13300);
   U774 : BUF_X1 port map( A => n6730, Z => n13318);
   U775 : BUF_X1 port map( A => n6723, Z => n13327);
   U776 : BUF_X1 port map( A => n6712, Z => n13345);
   U777 : BUF_X1 port map( A => n6706, Z => n13354);
   U778 : BUF_X1 port map( A => n6703, Z => n13363);
   U779 : BUF_X1 port map( A => n6697, Z => n13381);
   U780 : BUF_X1 port map( A => n6694, Z => n13390);
   U781 : BUF_X1 port map( A => n6691, Z => n13399);
   U782 : BUF_X1 port map( A => n6688, Z => n13408);
   U783 : BUF_X1 port map( A => n6683, Z => n13417);
   U784 : BUF_X1 port map( A => n6676, Z => n13435);
   U785 : BUF_X1 port map( A => n6673, Z => n13444);
   U786 : BUF_X1 port map( A => n6667, Z => n13462);
   U787 : BUF_X1 port map( A => n6664, Z => n13471);
   U788 : BUF_X1 port map( A => n6661, Z => n13480);
   U789 : BUF_X1 port map( A => n6658, Z => n13489);
   U790 : BUF_X1 port map( A => n6655, Z => n13498);
   U791 : BUF_X1 port map( A => n6652, Z => n13507);
   U792 : BUF_X1 port map( A => n6649, Z => n13516);
   U793 : BUF_X1 port map( A => n6646, Z => n13525);
   U794 : BUF_X1 port map( A => n6640, Z => n13543);
   U795 : BUF_X1 port map( A => n6637, Z => n13552);
   U796 : BUF_X1 port map( A => n6632, Z => n13561);
   U797 : BUF_X1 port map( A => n6626, Z => n13579);
   U798 : BUF_X1 port map( A => n6623, Z => n13588);
   U799 : BUF_X1 port map( A => n6620, Z => n13597);
   U800 : BUF_X1 port map( A => n6617, Z => n13606);
   U801 : BUF_X1 port map( A => n6611, Z => n13624);
   U802 : BUF_X1 port map( A => n2767, Z => n14313);
   U803 : INV_X1 port map( A => n13223, ZN => n14116);
   U804 : BUF_X1 port map( A => n5308, Z => n13802);
   U805 : BUF_X1 port map( A => n5349, Z => n13721);
   U806 : BUF_X1 port map( A => n4028, Z => n13941);
   U807 : BUF_X1 port map( A => n4028, Z => n13942);
   U808 : BUF_X1 port map( A => n5308, Z => n13803);
   U809 : BUF_X1 port map( A => n5349, Z => n13722);
   U810 : BUF_X1 port map( A => n5386, Z => n13640);
   U811 : BUF_X1 port map( A => n3987, Z => n14022);
   U812 : BUF_X1 port map( A => n3987, Z => n14023);
   U813 : BUF_X1 port map( A => n5386, Z => n13641);
   U814 : BUF_X1 port map( A => n5297, Z => n13829);
   U815 : BUF_X1 port map( A => n3976, Z => n14049);
   U816 : BUF_X1 port map( A => n5323, Z => n13775);
   U817 : BUF_X1 port map( A => n5334, Z => n13748);
   U818 : BUF_X1 port map( A => n5360, Z => n13694);
   U819 : BUF_X1 port map( A => n4013, Z => n13968);
   U820 : BUF_X1 port map( A => n4002, Z => n13995);
   U821 : BUF_X1 port map( A => n3976, Z => n14050);
   U822 : BUF_X1 port map( A => n4002, Z => n13996);
   U823 : BUF_X1 port map( A => n4013, Z => n13969);
   U824 : BUF_X1 port map( A => n5297, Z => n13830);
   U825 : BUF_X1 port map( A => n5323, Z => n13776);
   U826 : BUF_X1 port map( A => n5334, Z => n13749);
   U827 : BUF_X1 port map( A => n5360, Z => n13695);
   U828 : BUF_X1 port map( A => n2877, Z => n14089);
   U829 : BUF_X1 port map( A => n2877, Z => n14088);
   U830 : BUF_X1 port map( A => n4063, Z => n13872);
   U831 : BUF_X1 port map( A => n4063, Z => n13873);
   U832 : BUF_X1 port map( A => n2763, Z => n14322);
   U833 : BUF_X1 port map( A => n2763, Z => n14321);
   U834 : BUF_X1 port map( A => n2746, Z => n14360);
   U835 : BUF_X1 port map( A => n2746, Z => n14359);
   U836 : BUF_X1 port map( A => n2775, Z => n14291);
   U837 : BUF_X1 port map( A => n2775, Z => n14290);
   U838 : BUF_X1 port map( A => n2771, Z => n14302);
   U839 : BUF_X1 port map( A => n2771, Z => n14301);
   U840 : BUF_X1 port map( A => n2759, Z => n14331);
   U841 : BUF_X1 port map( A => n2759, Z => n14330);
   U842 : BUF_X1 port map( A => n2755, Z => n14340);
   U843 : BUF_X1 port map( A => n2755, Z => n14339);
   U844 : BUF_X1 port map( A => n2751, Z => n14349);
   U845 : BUF_X1 port map( A => n2751, Z => n14348);
   U846 : BUF_X1 port map( A => n3995, Z => n14014);
   U847 : BUF_X1 port map( A => n4032, Z => n13933);
   U848 : BUF_X1 port map( A => n4056, Z => n13891);
   U849 : BUF_X1 port map( A => n4021, Z => n13960);
   U850 : BUF_X1 port map( A => n2852, Z => n14135);
   U851 : BUF_X1 port map( A => n2624, Z => n14707);
   U852 : INV_X1 port map( A => n13224, ZN => n14307);
   U853 : BUF_X1 port map( A => n2624, Z => n14708);
   U854 : BUF_X1 port map( A => n2791, Z => n14262);
   U855 : BUF_X1 port map( A => n2828, Z => n14181);
   U856 : BUF_X1 port map( A => n2791, Z => n14261);
   U857 : BUF_X1 port map( A => n2828, Z => n14180);
   U858 : INV_X1 port map( A => n13222, ZN => n14297);
   U859 : INV_X1 port map( A => n2739, ZN => n2578);
   U860 : INV_X1 port map( A => n2692, ZN => n2575);
   U861 : BUF_X1 port map( A => n5278, Z => n13858);
   U862 : BUF_X1 port map( A => n3957, Z => n14078);
   U863 : INV_X1 port map( A => n2702, ZN => n2574);
   U864 : INV_X1 port map( A => n2729, ZN => n2579);
   U865 : BUF_X1 port map( A => n2851, Z => n14137);
   U866 : BUF_X1 port map( A => n2851, Z => n14138);
   U867 : BUF_X1 port map( A => n2790, Z => n14265);
   U868 : BUF_X1 port map( A => n2801, Z => n14238);
   U869 : BUF_X1 port map( A => n2816, Z => n14211);
   U870 : BUF_X1 port map( A => n2827, Z => n14184);
   U871 : BUF_X1 port map( A => n2790, Z => n14264);
   U872 : BUF_X1 port map( A => n2801, Z => n14237);
   U873 : BUF_X1 port map( A => n2816, Z => n14210);
   U874 : BUF_X1 port map( A => n2827, Z => n14183);
   U875 : BUF_X1 port map( A => n5298, Z => n13826);
   U876 : BUF_X1 port map( A => n5304, Z => n13811);
   U877 : BUF_X1 port map( A => n3977, Z => n14046);
   U878 : BUF_X1 port map( A => n3983, Z => n14031);
   U879 : BUF_X1 port map( A => n3977, Z => n14047);
   U880 : BUF_X1 port map( A => n3983, Z => n14032);
   U881 : BUF_X1 port map( A => n5298, Z => n13827);
   U882 : BUF_X1 port map( A => n5304, Z => n13812);
   U883 : BUF_X1 port map( A => n5293, Z => n13838);
   U884 : BUF_X1 port map( A => n5287, Z => n13853);
   U885 : BUF_X1 port map( A => n5313, Z => n13799);
   U886 : BUF_X1 port map( A => n5319, Z => n13784);
   U887 : BUF_X1 port map( A => n5330, Z => n13757);
   U888 : BUF_X1 port map( A => n5324, Z => n13772);
   U889 : BUF_X1 port map( A => n5339, Z => n13745);
   U890 : BUF_X1 port map( A => n5350, Z => n13718);
   U891 : BUF_X1 port map( A => n5345, Z => n13730);
   U892 : BUF_X1 port map( A => n5356, Z => n13703);
   U893 : BUF_X1 port map( A => n5376, Z => n13664);
   U894 : BUF_X1 port map( A => n5382, Z => n13649);
   U895 : BUF_X1 port map( A => n3972, Z => n14058);
   U896 : BUF_X1 port map( A => n3966, Z => n14073);
   U897 : BUF_X1 port map( A => n4009, Z => n13977);
   U898 : BUF_X1 port map( A => n4003, Z => n13992);
   U899 : BUF_X1 port map( A => n2787, Z => n14270);
   U900 : BUF_X1 port map( A => n2813, Z => n14216);
   U901 : BUF_X1 port map( A => n2824, Z => n14189);
   U902 : BUF_X1 port map( A => n2848, Z => n14143);
   U903 : BUF_X1 port map( A => n3992, Z => n14019);
   U904 : BUF_X1 port map( A => n3998, Z => n14004);
   U905 : BUF_X1 port map( A => n4018, Z => n13965);
   U906 : BUF_X1 port map( A => n4029, Z => n13938);
   U907 : BUF_X1 port map( A => n4024, Z => n13950);
   U908 : BUF_X1 port map( A => n4053, Z => n13896);
   U909 : BUF_X1 port map( A => n4059, Z => n13881);
   U910 : BUF_X1 port map( A => n3966, Z => n14074);
   U911 : BUF_X1 port map( A => n3972, Z => n14059);
   U912 : BUF_X1 port map( A => n3992, Z => n14020);
   U913 : BUF_X1 port map( A => n3998, Z => n14005);
   U914 : BUF_X1 port map( A => n4009, Z => n13978);
   U915 : BUF_X1 port map( A => n4003, Z => n13993);
   U916 : BUF_X1 port map( A => n4018, Z => n13966);
   U917 : BUF_X1 port map( A => n4029, Z => n13939);
   U918 : BUF_X1 port map( A => n4024, Z => n13951);
   U919 : BUF_X1 port map( A => n4053, Z => n13897);
   U920 : BUF_X1 port map( A => n4059, Z => n13882);
   U921 : BUF_X1 port map( A => n5287, Z => n13854);
   U922 : BUF_X1 port map( A => n5293, Z => n13839);
   U923 : BUF_X1 port map( A => n5313, Z => n13800);
   U924 : BUF_X1 port map( A => n5319, Z => n13785);
   U925 : BUF_X1 port map( A => n5330, Z => n13758);
   U926 : BUF_X1 port map( A => n5324, Z => n13773);
   U927 : BUF_X1 port map( A => n5339, Z => n13746);
   U928 : BUF_X1 port map( A => n5350, Z => n13719);
   U929 : BUF_X1 port map( A => n5345, Z => n13731);
   U930 : BUF_X1 port map( A => n5356, Z => n13704);
   U931 : BUF_X1 port map( A => n5376, Z => n13665);
   U932 : BUF_X1 port map( A => n5382, Z => n13650);
   U933 : BUF_X1 port map( A => n2839, Z => n14163);
   U934 : BUF_X1 port map( A => n2813, Z => n14217);
   U935 : BUF_X1 port map( A => n2824, Z => n14190);
   U936 : BUF_X1 port map( A => n2848, Z => n14144);
   U937 : BUF_X1 port map( A => n2787, Z => n14271);
   U938 : BUF_X1 port map( A => n2839, Z => n14162);
   U939 : BUF_X1 port map( A => n2797, Z => n14247);
   U940 : BUF_X1 port map( A => n2823, Z => n14193);
   U941 : BUF_X1 port map( A => n2834, Z => n14166);
   U942 : BUF_X1 port map( A => n2858, Z => n14120);
   U943 : BUF_X1 port map( A => n2797, Z => n14246);
   U944 : BUF_X1 port map( A => n2823, Z => n14192);
   U945 : BUF_X1 port map( A => n2834, Z => n14165);
   U946 : BUF_X1 port map( A => n2858, Z => n14119);
   U947 : BUF_X1 port map( A => n5299, Z => n13823);
   U948 : BUF_X1 port map( A => n5305, Z => n13808);
   U949 : BUF_X1 port map( A => n3978, Z => n14043);
   U950 : BUF_X1 port map( A => n3984, Z => n14028);
   U951 : BUF_X1 port map( A => n3978, Z => n14044);
   U952 : BUF_X1 port map( A => n3984, Z => n14029);
   U953 : BUF_X1 port map( A => n5299, Z => n13824);
   U954 : BUF_X1 port map( A => n5305, Z => n13809);
   U955 : BUF_X1 port map( A => n5294, Z => n13835);
   U956 : BUF_X1 port map( A => n5288, Z => n13850);
   U957 : BUF_X1 port map( A => n5314, Z => n13796);
   U958 : BUF_X1 port map( A => n5320, Z => n13781);
   U959 : BUF_X1 port map( A => n5331, Z => n13754);
   U960 : BUF_X1 port map( A => n5325, Z => n13769);
   U961 : BUF_X1 port map( A => n5340, Z => n13742);
   U962 : BUF_X1 port map( A => n5351, Z => n13715);
   U963 : BUF_X1 port map( A => n5346, Z => n13727);
   U964 : BUF_X1 port map( A => n5357, Z => n13700);
   U965 : BUF_X1 port map( A => n5377, Z => n13661);
   U966 : BUF_X1 port map( A => n5383, Z => n13646);
   U967 : BUF_X1 port map( A => n3973, Z => n14055);
   U968 : BUF_X1 port map( A => n3967, Z => n14070);
   U969 : BUF_X1 port map( A => n3999, Z => n14001);
   U970 : BUF_X1 port map( A => n4010, Z => n13974);
   U971 : BUF_X1 port map( A => n4004, Z => n13989);
   U972 : BUF_X1 port map( A => n3967, Z => n14071);
   U973 : BUF_X1 port map( A => n3973, Z => n14056);
   U974 : BUF_X1 port map( A => n3999, Z => n14002);
   U975 : BUF_X1 port map( A => n4010, Z => n13975);
   U976 : BUF_X1 port map( A => n4004, Z => n13990);
   U977 : BUF_X1 port map( A => n5288, Z => n13851);
   U978 : BUF_X1 port map( A => n5294, Z => n13836);
   U979 : BUF_X1 port map( A => n5314, Z => n13797);
   U980 : BUF_X1 port map( A => n5320, Z => n13782);
   U981 : BUF_X1 port map( A => n5331, Z => n13755);
   U982 : BUF_X1 port map( A => n5325, Z => n13770);
   U983 : BUF_X1 port map( A => n5340, Z => n13743);
   U984 : BUF_X1 port map( A => n5351, Z => n13716);
   U985 : BUF_X1 port map( A => n5346, Z => n13728);
   U986 : BUF_X1 port map( A => n5357, Z => n13701);
   U987 : BUF_X1 port map( A => n5377, Z => n13662);
   U988 : BUF_X1 port map( A => n5383, Z => n13647);
   U989 : BUF_X1 port map( A => n2849, Z => n14141);
   U990 : BUF_X1 port map( A => n2840, Z => n14160);
   U991 : BUF_X1 port map( A => n2849, Z => n14140);
   U992 : BUF_X1 port map( A => n2840, Z => n14159);
   U993 : BUF_X1 port map( A => n2794, Z => n14254);
   U994 : BUF_X1 port map( A => n2825, Z => n14188);
   U995 : BUF_X1 port map( A => n2820, Z => n14200);
   U996 : BUF_X1 port map( A => n2831, Z => n14173);
   U997 : BUF_X1 port map( A => n2855, Z => n14127);
   U998 : BUF_X1 port map( A => n2793, Z => n14256);
   U999 : BUF_X1 port map( A => n2819, Z => n14202);
   U1000 : BUF_X1 port map( A => n2830, Z => n14175);
   U1001 : BUF_X1 port map( A => n2854, Z => n14129);
   U1002 : BUF_X1 port map( A => n2793, Z => n14255);
   U1003 : BUF_X1 port map( A => n2819, Z => n14201);
   U1004 : BUF_X1 port map( A => n2830, Z => n14174);
   U1005 : BUF_X1 port map( A => n2854, Z => n14128);
   U1006 : BUF_X1 port map( A => n2796, Z => n14250);
   U1007 : BUF_X1 port map( A => n2822, Z => n14196);
   U1008 : BUF_X1 port map( A => n2796, Z => n14249);
   U1009 : BUF_X1 port map( A => n2822, Z => n14195);
   U1010 : BUF_X1 port map( A => n2788, Z => n14269);
   U1011 : BUF_X1 port map( A => n6825, Z => n13226);
   U1012 : BUF_X1 port map( A => n6797, Z => n13253);
   U1013 : BUF_X1 port map( A => n6759, Z => n13280);
   U1014 : BUF_X1 port map( A => n6679, Z => n13424);
   U1015 : BUF_X1 port map( A => n6819, Z => n13235);
   U1016 : BUF_X1 port map( A => n6807, Z => n13244);
   U1017 : BUF_X1 port map( A => n6784, Z => n13262);
   U1018 : BUF_X1 port map( A => n6772, Z => n13271);
   U1019 : BUF_X1 port map( A => n6629, Z => n13568);
   U1020 : BUF_X1 port map( A => n6606, Z => n13631);
   U1021 : BUF_X1 port map( A => n2701, Z => n14437);
   U1022 : BUF_X1 port map( A => n2681, Z => n14473);
   U1023 : BUF_X1 port map( A => n2676, Z => n14482);
   U1024 : BUF_X1 port map( A => n6751, Z => n13289);
   U1025 : BUF_X1 port map( A => n6747, Z => n13298);
   U1026 : BUF_X1 port map( A => n6735, Z => n13307);
   U1027 : BUF_X1 port map( A => n6718, Z => n13334);
   U1028 : BUF_X1 port map( A => n6700, Z => n13370);
   U1029 : BUF_X1 port map( A => n6697, Z => n13379);
   U1030 : BUF_X1 port map( A => n6694, Z => n13388);
   U1031 : BUF_X1 port map( A => n6670, Z => n13451);
   U1032 : BUF_X1 port map( A => n6667, Z => n13460);
   U1033 : BUF_X1 port map( A => n6664, Z => n13469);
   U1034 : BUF_X1 port map( A => n6643, Z => n13532);
   U1035 : BUF_X1 port map( A => n6640, Z => n13541);
   U1036 : BUF_X1 port map( A => n6637, Z => n13550);
   U1037 : BUF_X1 port map( A => n2696, Z => n14446);
   U1038 : BUF_X1 port map( A => n6614, Z => n13613);
   U1039 : BUF_X1 port map( A => n6611, Z => n13622);
   U1040 : BUF_X1 port map( A => n2691, Z => n14455);
   U1041 : BUF_X1 port map( A => n2686, Z => n14464);
   U1042 : BUF_X1 port map( A => n2671, Z => n14491);
   U1043 : BUF_X1 port map( A => n2666, Z => n14500);
   U1044 : BUF_X1 port map( A => n6730, Z => n13316);
   U1045 : BUF_X1 port map( A => n6723, Z => n13325);
   U1046 : BUF_X1 port map( A => n6712, Z => n13343);
   U1047 : BUF_X1 port map( A => n6706, Z => n13352);
   U1048 : BUF_X1 port map( A => n6703, Z => n13361);
   U1049 : BUF_X1 port map( A => n6691, Z => n13397);
   U1050 : BUF_X1 port map( A => n6688, Z => n13406);
   U1051 : BUF_X1 port map( A => n6683, Z => n13415);
   U1052 : BUF_X1 port map( A => n6676, Z => n13433);
   U1053 : BUF_X1 port map( A => n6673, Z => n13442);
   U1054 : BUF_X1 port map( A => n6661, Z => n13478);
   U1055 : BUF_X1 port map( A => n6658, Z => n13487);
   U1056 : BUF_X1 port map( A => n6655, Z => n13496);
   U1057 : BUF_X1 port map( A => n6652, Z => n13505);
   U1058 : BUF_X1 port map( A => n6649, Z => n13514);
   U1059 : BUF_X1 port map( A => n6646, Z => n13523);
   U1060 : BUF_X1 port map( A => n6632, Z => n13559);
   U1061 : BUF_X1 port map( A => n6626, Z => n13577);
   U1062 : BUF_X1 port map( A => n6623, Z => n13586);
   U1063 : BUF_X1 port map( A => n6620, Z => n13595);
   U1064 : BUF_X1 port map( A => n6617, Z => n13604);
   U1065 : BUF_X1 port map( A => n5292, Z => n13841);
   U1066 : BUF_X1 port map( A => n3971, Z => n14061);
   U1067 : BUF_X1 port map( A => n3971, Z => n14062);
   U1068 : BUF_X1 port map( A => n5292, Z => n13842);
   U1069 : BUF_X1 port map( A => n5303, Z => n13814);
   U1070 : BUF_X1 port map( A => n3982, Z => n14034);
   U1071 : BUF_X1 port map( A => n3982, Z => n14035);
   U1072 : BUF_X1 port map( A => n5303, Z => n13815);
   U1073 : BUF_X1 port map( A => n5318, Z => n13787);
   U1074 : BUF_X1 port map( A => n5329, Z => n13760);
   U1075 : BUF_X1 port map( A => n5344, Z => n13733);
   U1076 : BUF_X1 port map( A => n5355, Z => n13706);
   U1077 : BUF_X1 port map( A => n5318, Z => n13788);
   U1078 : BUF_X1 port map( A => n5329, Z => n13761);
   U1079 : BUF_X1 port map( A => n5344, Z => n13734);
   U1080 : BUF_X1 port map( A => n2844, Z => n14151);
   U1081 : BUF_X1 port map( A => n2844, Z => n14150);
   U1082 : BUF_X1 port map( A => n5381, Z => n13652);
   U1083 : BUF_X1 port map( A => n5355, Z => n13707);
   U1084 : BUF_X1 port map( A => n4008, Z => n13980);
   U1085 : BUF_X1 port map( A => n4008, Z => n13981);
   U1086 : BUF_X1 port map( A => n5381, Z => n13653);
   U1087 : BUF_X1 port map( A => n2872, Z => n14101);
   U1088 : BUF_X1 port map( A => n2872, Z => n14100);
   U1089 : BUF_X1 port map( A => n6606, Z => n13632);
   U1090 : BUF_X1 port map( A => n2681, Z => n14474);
   U1091 : BUF_X1 port map( A => n2676, Z => n14483);
   U1092 : BUF_X1 port map( A => n6751, Z => n13290);
   U1093 : BUF_X1 port map( A => n6718, Z => n13335);
   U1094 : BUF_X1 port map( A => n6712, Z => n13344);
   U1095 : BUF_X1 port map( A => n6700, Z => n13371);
   U1096 : BUF_X1 port map( A => n6670, Z => n13452);
   U1097 : BUF_X1 port map( A => n6643, Z => n13533);
   U1098 : BUF_X1 port map( A => n6614, Z => n13614);
   U1099 : BUF_X1 port map( A => n2701, Z => n14438);
   U1100 : BUF_X1 port map( A => n2696, Z => n14447);
   U1101 : BUF_X1 port map( A => n2691, Z => n14456);
   U1102 : BUF_X1 port map( A => n2686, Z => n14465);
   U1103 : BUF_X1 port map( A => n2671, Z => n14492);
   U1104 : BUF_X1 port map( A => n2666, Z => n14501);
   U1105 : BUF_X1 port map( A => n6747, Z => n13299);
   U1106 : BUF_X1 port map( A => n6735, Z => n13308);
   U1107 : BUF_X1 port map( A => n6730, Z => n13317);
   U1108 : BUF_X1 port map( A => n6723, Z => n13326);
   U1109 : BUF_X1 port map( A => n6706, Z => n13353);
   U1110 : BUF_X1 port map( A => n6703, Z => n13362);
   U1111 : BUF_X1 port map( A => n6697, Z => n13380);
   U1112 : BUF_X1 port map( A => n6694, Z => n13389);
   U1113 : BUF_X1 port map( A => n6691, Z => n13398);
   U1114 : BUF_X1 port map( A => n6688, Z => n13407);
   U1115 : BUF_X1 port map( A => n6683, Z => n13416);
   U1116 : BUF_X1 port map( A => n6676, Z => n13434);
   U1117 : BUF_X1 port map( A => n6673, Z => n13443);
   U1118 : BUF_X1 port map( A => n6667, Z => n13461);
   U1119 : BUF_X1 port map( A => n6664, Z => n13470);
   U1120 : BUF_X1 port map( A => n6661, Z => n13479);
   U1121 : BUF_X1 port map( A => n6658, Z => n13488);
   U1122 : BUF_X1 port map( A => n6655, Z => n13497);
   U1123 : BUF_X1 port map( A => n6652, Z => n13506);
   U1124 : BUF_X1 port map( A => n6649, Z => n13515);
   U1125 : BUF_X1 port map( A => n6646, Z => n13524);
   U1126 : BUF_X1 port map( A => n6640, Z => n13542);
   U1127 : BUF_X1 port map( A => n6637, Z => n13551);
   U1128 : BUF_X1 port map( A => n6632, Z => n13560);
   U1129 : BUF_X1 port map( A => n6626, Z => n13578);
   U1130 : BUF_X1 port map( A => n6623, Z => n13587);
   U1131 : BUF_X1 port map( A => n6620, Z => n13596);
   U1132 : BUF_X1 port map( A => n6617, Z => n13605);
   U1133 : BUF_X1 port map( A => n6611, Z => n13623);
   U1134 : INV_X1 port map( A => n2687, ZN => n2571);
   U1135 : BUF_X1 port map( A => n3986, Z => n14027);
   U1136 : BUF_X1 port map( A => n5307, Z => n13807);
   U1137 : BUF_X1 port map( A => n3975, Z => n14054);
   U1138 : BUF_X1 port map( A => n4012, Z => n13973);
   U1139 : BUF_X1 port map( A => n5296, Z => n13834);
   U1140 : BUF_X1 port map( A => n5322, Z => n13780);
   U1141 : BUF_X1 port map( A => n5333, Z => n13753);
   U1142 : BUF_X1 port map( A => n2876, Z => n14093);
   U1143 : BUF_X1 port map( A => n5359, Z => n13699);
   U1144 : BUF_X1 port map( A => n5348, Z => n13726);
   U1145 : BUF_X1 port map( A => n5385, Z => n13645);
   U1146 : INV_X1 port map( A => n2661, ZN => n2585);
   U1147 : BUF_X1 port map( A => n6628, Z => n13572);
   U1148 : BUF_X1 port map( A => n6628, Z => n13571);
   U1149 : BUF_X1 port map( A => n6604, Z => n13638);
   U1150 : BUF_X1 port map( A => n6604, Z => n13637);
   U1151 : BUF_X1 port map( A => n2763, Z => n14323);
   U1152 : BUF_X1 port map( A => n2746, Z => n14361);
   U1153 : BUF_X1 port map( A => n6613, Z => n13617);
   U1154 : BUF_X1 port map( A => n6613, Z => n13616);
   U1155 : BUF_X1 port map( A => n6610, Z => n13625);
   U1156 : BUF_X1 port map( A => n6625, Z => n13581);
   U1157 : BUF_X1 port map( A => n6625, Z => n13580);
   U1158 : BUF_X1 port map( A => n6622, Z => n13590);
   U1159 : BUF_X1 port map( A => n6622, Z => n13589);
   U1160 : BUF_X1 port map( A => n6619, Z => n13599);
   U1161 : BUF_X1 port map( A => n6619, Z => n13598);
   U1162 : BUF_X1 port map( A => n6616, Z => n13608);
   U1163 : BUF_X1 port map( A => n6616, Z => n13607);
   U1164 : BUF_X1 port map( A => n6610, Z => n13626);
   U1165 : INV_X1 port map( A => n2667, ZN => n2573);
   U1166 : BUF_X1 port map( A => n2792, Z => n14260);
   U1167 : BUF_X1 port map( A => n2818, Z => n14206);
   U1168 : BUF_X1 port map( A => n2829, Z => n14179);
   U1169 : BUF_X1 port map( A => n5301, Z => n13820);
   U1170 : BUF_X1 port map( A => n3980, Z => n14040);
   U1171 : BUF_X1 port map( A => n3980, Z => n14041);
   U1172 : BUF_X1 port map( A => n5301, Z => n13821);
   U1173 : BUF_X1 port map( A => n5379, Z => n13658);
   U1174 : BUF_X1 port map( A => n5379, Z => n13659);
   U1175 : BUF_X1 port map( A => n5290, Z => n13847);
   U1176 : BUF_X1 port map( A => n5316, Z => n13793);
   U1177 : BUF_X1 port map( A => n5327, Z => n13766);
   U1178 : BUF_X1 port map( A => n5353, Z => n13712);
   U1179 : BUF_X1 port map( A => n4006, Z => n13986);
   U1180 : BUF_X1 port map( A => n4006, Z => n13987);
   U1181 : BUF_X1 port map( A => n5290, Z => n13848);
   U1182 : BUF_X1 port map( A => n5327, Z => n13767);
   U1183 : BUF_X1 port map( A => n5353, Z => n13713);
   U1184 : BUF_X1 port map( A => n2842, Z => n14157);
   U1185 : BUF_X1 port map( A => n2842, Z => n14156);
   U1186 : BUF_X1 port map( A => n6797, Z => n13255);
   U1187 : BUF_X1 port map( A => n6819, Z => n13237);
   U1188 : BUF_X1 port map( A => n6807, Z => n13246);
   U1189 : BUF_X1 port map( A => n6784, Z => n13264);
   U1190 : BUF_X1 port map( A => n6772, Z => n13273);
   U1191 : BUF_X1 port map( A => n5316, Z => n13794);
   U1192 : BUF_X1 port map( A => n6759, Z => n13282);
   U1193 : BUF_X1 port map( A => n6679, Z => n13426);
   U1194 : BUF_X1 port map( A => n6629, Z => n13570);
   U1195 : BUF_X1 port map( A => n5342, Z => n13739);
   U1196 : BUF_X1 port map( A => n3969, Z => n14067);
   U1197 : BUF_X1 port map( A => n3969, Z => n14068);
   U1198 : BUF_X1 port map( A => n5342, Z => n13740);
   U1199 : BUF_X1 port map( A => n5328, Z => n13763);
   U1200 : BUF_X1 port map( A => n4007, Z => n13983);
   U1201 : BUF_X1 port map( A => n4007, Z => n13984);
   U1202 : BUF_X1 port map( A => n5328, Z => n13764);
   U1203 : BUF_X1 port map( A => n2870, Z => n14107);
   U1204 : BUF_X1 port map( A => n2870, Z => n14106);
   U1205 : BUF_X1 port map( A => n5302, Z => n13817);
   U1206 : BUF_X1 port map( A => n3981, Z => n14037);
   U1207 : BUF_X1 port map( A => n3981, Z => n14038);
   U1208 : BUF_X1 port map( A => n5302, Z => n13818);
   U1209 : BUF_X1 port map( A => n4022, Z => n13956);
   U1210 : BUF_X1 port map( A => n5354, Z => n13709);
   U1211 : BUF_X1 port map( A => n4057, Z => n13887);
   U1212 : BUF_X1 port map( A => n4022, Z => n13957);
   U1213 : BUF_X1 port map( A => n5317, Z => n13790);
   U1214 : BUF_X1 port map( A => n4057, Z => n13888);
   U1215 : BUF_X1 port map( A => n5343, Z => n13736);
   U1216 : BUF_X1 port map( A => n5380, Z => n13655);
   U1217 : BUF_X1 port map( A => n4033, Z => n13929);
   U1218 : BUF_X1 port map( A => n4033, Z => n13930);
   U1219 : BUF_X1 port map( A => n5317, Z => n13791);
   U1220 : BUF_X1 port map( A => n5343, Z => n13737);
   U1221 : BUF_X1 port map( A => n5354, Z => n13710);
   U1222 : BUF_X1 port map( A => n5380, Z => n13656);
   U1223 : BUF_X1 port map( A => n2843, Z => n14154);
   U1224 : BUF_X1 port map( A => n2843, Z => n14153);
   U1225 : BUF_X1 port map( A => n3996, Z => n14010);
   U1226 : BUF_X1 port map( A => n3996, Z => n14011);
   U1227 : BUF_X1 port map( A => n5291, Z => n13844);
   U1228 : BUF_X1 port map( A => n3970, Z => n14064);
   U1229 : BUF_X1 port map( A => n3970, Z => n14065);
   U1230 : BUF_X1 port map( A => n5291, Z => n13845);
   U1231 : BUF_X1 port map( A => n2817, Z => n14208);
   U1232 : BUF_X1 port map( A => n2871, Z => n14104);
   U1233 : BUF_X1 port map( A => n2817, Z => n14207);
   U1234 : BUF_X1 port map( A => n2871, Z => n14103);
   U1235 : BUF_X1 port map( A => n5308, Z => n13804);
   U1236 : BUF_X1 port map( A => n5349, Z => n13723);
   U1237 : BUF_X1 port map( A => n5386, Z => n13642);
   U1238 : BUF_X1 port map( A => n3987, Z => n14024);
   U1239 : BUF_X1 port map( A => n2755, Z => n14341);
   U1240 : BUF_X1 port map( A => n2775, Z => n14292);
   U1241 : BUF_X1 port map( A => n2771, Z => n14303);
   U1242 : BUF_X1 port map( A => n2759, Z => n14332);
   U1243 : BUF_X1 port map( A => n3976, Z => n14051);
   U1244 : BUF_X1 port map( A => n4013, Z => n13970);
   U1245 : BUF_X1 port map( A => n5297, Z => n13831);
   U1246 : BUF_X1 port map( A => n5334, Z => n13750);
   U1247 : BUF_X1 port map( A => n5323, Z => n13777);
   U1248 : BUF_X1 port map( A => n5360, Z => n13696);
   U1249 : BUF_X1 port map( A => n2877, Z => n14090);
   U1250 : BUF_X1 port map( A => n4001, Z => n14000);
   U1251 : BUF_X1 port map( A => n4062, Z => n13877);
   U1252 : BUF_X1 port map( A => n4027, Z => n13946);
   U1253 : BUF_X1 port map( A => n2853, Z => n14133);
   U1254 : INV_X1 port map( A => n2697, ZN => n2570);
   U1255 : BUF_X1 port map( A => n6825, Z => n13228);
   U1256 : BUF_X1 port map( A => n2791, Z => n14263);
   U1257 : BUF_X1 port map( A => n2828, Z => n14182);
   U1258 : INV_X1 port map( A => n2714, ZN => n2584);
   U1259 : INV_X1 port map( A => n2734, ZN => n2582);
   U1260 : BUF_X1 port map( A => n2751, Z => n14350);
   U1261 : BUF_X1 port map( A => n4028, Z => n13943);
   U1262 : BUF_X1 port map( A => n4002, Z => n13997);
   U1263 : BUF_X1 port map( A => n4063, Z => n13874);
   U1264 : BUF_X1 port map( A => n2790, Z => n14266);
   U1265 : BUF_X1 port map( A => n2801, Z => n14239);
   U1266 : BUF_X1 port map( A => n2816, Z => n14212);
   U1267 : BUF_X1 port map( A => n2827, Z => n14185);
   U1268 : BUF_X1 port map( A => n3977, Z => n14048);
   U1269 : BUF_X1 port map( A => n3983, Z => n14033);
   U1270 : BUF_X1 port map( A => n5298, Z => n13828);
   U1271 : BUF_X1 port map( A => n5304, Z => n13813);
   U1272 : BUF_X1 port map( A => n3966, Z => n14075);
   U1273 : BUF_X1 port map( A => n3972, Z => n14060);
   U1274 : BUF_X1 port map( A => n4009, Z => n13979);
   U1275 : BUF_X1 port map( A => n4003, Z => n13994);
   U1276 : BUF_X1 port map( A => n5287, Z => n13855);
   U1277 : BUF_X1 port map( A => n5293, Z => n13840);
   U1278 : BUF_X1 port map( A => n5313, Z => n13801);
   U1279 : BUF_X1 port map( A => n5319, Z => n13786);
   U1280 : BUF_X1 port map( A => n5330, Z => n13759);
   U1281 : BUF_X1 port map( A => n5324, Z => n13774);
   U1282 : BUF_X1 port map( A => n5339, Z => n13747);
   U1283 : BUF_X1 port map( A => n5350, Z => n13720);
   U1284 : BUF_X1 port map( A => n5345, Z => n13732);
   U1285 : BUF_X1 port map( A => n5356, Z => n13705);
   U1286 : BUF_X1 port map( A => n5376, Z => n13666);
   U1287 : BUF_X1 port map( A => n5382, Z => n13651);
   U1288 : BUF_X1 port map( A => n2839, Z => n14164);
   U1289 : INV_X1 port map( A => n2707, ZN => n2528);
   U1290 : BUF_X1 port map( A => n2813, Z => n14218);
   U1291 : BUF_X1 port map( A => n2824, Z => n14191);
   U1292 : BUF_X1 port map( A => n2848, Z => n14145);
   U1293 : BUF_X1 port map( A => n3992, Z => n14021);
   U1294 : BUF_X1 port map( A => n3998, Z => n14006);
   U1295 : BUF_X1 port map( A => n4018, Z => n13967);
   U1296 : BUF_X1 port map( A => n4029, Z => n13940);
   U1297 : BUF_X1 port map( A => n4024, Z => n13952);
   U1298 : BUF_X1 port map( A => n4053, Z => n13898);
   U1299 : BUF_X1 port map( A => n4059, Z => n13883);
   U1300 : BUF_X1 port map( A => n2787, Z => n14272);
   U1301 : BUF_X1 port map( A => n2851, Z => n14139);
   U1302 : BUF_X1 port map( A => n2797, Z => n14248);
   U1303 : BUF_X1 port map( A => n2823, Z => n14194);
   U1304 : BUF_X1 port map( A => n2834, Z => n14167);
   U1305 : BUF_X1 port map( A => n2858, Z => n14121);
   U1306 : BUF_X1 port map( A => n3978, Z => n14045);
   U1307 : BUF_X1 port map( A => n3984, Z => n14030);
   U1308 : BUF_X1 port map( A => n5299, Z => n13825);
   U1309 : BUF_X1 port map( A => n5305, Z => n13810);
   U1310 : BUF_X1 port map( A => n3967, Z => n14072);
   U1311 : BUF_X1 port map( A => n3973, Z => n14057);
   U1312 : BUF_X1 port map( A => n3999, Z => n14003);
   U1313 : BUF_X1 port map( A => n4010, Z => n13976);
   U1314 : BUF_X1 port map( A => n4004, Z => n13991);
   U1315 : BUF_X1 port map( A => n5288, Z => n13852);
   U1316 : BUF_X1 port map( A => n5294, Z => n13837);
   U1317 : BUF_X1 port map( A => n5314, Z => n13798);
   U1318 : BUF_X1 port map( A => n5320, Z => n13783);
   U1319 : BUF_X1 port map( A => n5331, Z => n13756);
   U1320 : BUF_X1 port map( A => n5325, Z => n13771);
   U1321 : BUF_X1 port map( A => n5340, Z => n13744);
   U1322 : BUF_X1 port map( A => n5351, Z => n13717);
   U1323 : BUF_X1 port map( A => n5346, Z => n13729);
   U1324 : BUF_X1 port map( A => n5357, Z => n13702);
   U1325 : BUF_X1 port map( A => n5377, Z => n13663);
   U1326 : BUF_X1 port map( A => n5383, Z => n13648);
   U1327 : BUF_X1 port map( A => n2849, Z => n14142);
   U1328 : BUF_X1 port map( A => n2840, Z => n14161);
   U1329 : BUF_X1 port map( A => n2793, Z => n14257);
   U1330 : BUF_X1 port map( A => n2819, Z => n14203);
   U1331 : BUF_X1 port map( A => n2830, Z => n14176);
   U1332 : BUF_X1 port map( A => n2854, Z => n14130);
   U1333 : BUF_X1 port map( A => n2796, Z => n14251);
   U1334 : BUF_X1 port map( A => n2822, Z => n14197);
   U1335 : BUF_X1 port map( A => n6628, Z => n13573);
   U1336 : BUF_X1 port map( A => n3971, Z => n14063);
   U1337 : BUF_X1 port map( A => n5292, Z => n13843);
   U1338 : BUF_X1 port map( A => n3982, Z => n14036);
   U1339 : BUF_X1 port map( A => n5303, Z => n13816);
   U1340 : BUF_X1 port map( A => n6604, Z => n13639);
   U1341 : BUF_X1 port map( A => n5318, Z => n13789);
   U1342 : BUF_X1 port map( A => n5329, Z => n13762);
   U1343 : BUF_X1 port map( A => n5344, Z => n13735);
   U1344 : BUF_X1 port map( A => n5355, Z => n13708);
   U1345 : BUF_X1 port map( A => n2844, Z => n14152);
   U1346 : BUF_X1 port map( A => n4008, Z => n13982);
   U1347 : BUF_X1 port map( A => n5381, Z => n13654);
   U1348 : BUF_X1 port map( A => n2872, Z => n14102);
   U1349 : BUF_X1 port map( A => n6613, Z => n13618);
   U1350 : BUF_X1 port map( A => n6625, Z => n13582);
   U1351 : BUF_X1 port map( A => n6622, Z => n13591);
   U1352 : BUF_X1 port map( A => n6619, Z => n13600);
   U1353 : BUF_X1 port map( A => n6616, Z => n13609);
   U1354 : BUF_X1 port map( A => n6610, Z => n13627);
   U1355 : BUF_X1 port map( A => n3980, Z => n14042);
   U1356 : BUF_X1 port map( A => n5301, Z => n13822);
   U1357 : BUF_X1 port map( A => n5379, Z => n13660);
   U1358 : BUF_X1 port map( A => n4007, Z => n13985);
   U1359 : BUF_X1 port map( A => n5328, Z => n13765);
   U1360 : BUF_X1 port map( A => n4006, Z => n13988);
   U1361 : BUF_X1 port map( A => n5290, Z => n13849);
   U1362 : BUF_X1 port map( A => n5327, Z => n13768);
   U1363 : BUF_X1 port map( A => n5353, Z => n13714);
   U1364 : BUF_X1 port map( A => n2842, Z => n14158);
   U1365 : BUF_X1 port map( A => n5302, Z => n13819);
   U1366 : BUF_X1 port map( A => n5316, Z => n13795);
   U1367 : BUF_X1 port map( A => n3981, Z => n14039);
   U1368 : BUF_X1 port map( A => n3969, Z => n14069);
   U1369 : BUF_X1 port map( A => n5342, Z => n13741);
   U1370 : BUF_X1 port map( A => n2870, Z => n14108);
   U1371 : BUF_X1 port map( A => n4022, Z => n13958);
   U1372 : BUF_X1 port map( A => n4033, Z => n13931);
   U1373 : BUF_X1 port map( A => n4057, Z => n13889);
   U1374 : BUF_X1 port map( A => n5317, Z => n13792);
   U1375 : BUF_X1 port map( A => n5354, Z => n13711);
   U1376 : BUF_X1 port map( A => n5343, Z => n13738);
   U1377 : BUF_X1 port map( A => n5380, Z => n13657);
   U1378 : BUF_X1 port map( A => n2843, Z => n14155);
   U1379 : BUF_X1 port map( A => n3996, Z => n14012);
   U1380 : BUF_X1 port map( A => n3970, Z => n14066);
   U1381 : BUF_X1 port map( A => n5291, Z => n13846);
   U1382 : BUF_X1 port map( A => n2817, Z => n14209);
   U1383 : BUF_X1 port map( A => n2871, Z => n14105);
   U1384 : INV_X1 port map( A => n2724, ZN => n2583);
   U1385 : BUF_X1 port map( A => n2624, Z => n14709);
   U1386 : INV_X1 port map( A => n2719, ZN => n2580);
   U1387 : BUF_X1 port map( A => n2630, Z => n14685);
   U1388 : BUF_X1 port map( A => n2833, Z => n14170);
   U1389 : BUF_X1 port map( A => n2857, Z => n14124);
   U1390 : NOR2_X1 port map( A1 => n2714, A2 => n2563, ZN => n2874);
   U1391 : NOR2_X1 port map( A1 => n2724, A2 => n2563, ZN => n2868);
   U1392 : AND2_X1 port map( A1 => n6777, A2 => n6714, ZN => n2709);
   U1393 : BUF_X1 port map( A => n2767, Z => n14314);
   U1394 : BUF_X1 port map( A => n3993, Z => n14018);
   U1395 : BUF_X1 port map( A => n4019, Z => n13964);
   U1396 : BUF_X1 port map( A => n4030, Z => n13937);
   U1397 : BUF_X1 port map( A => n4025, Z => n13949);
   U1398 : BUF_X1 port map( A => n4054, Z => n13895);
   U1399 : BUF_X1 port map( A => n4060, Z => n13880);
   U1400 : BUF_X1 port map( A => n2814, Z => n14215);
   U1401 : BUF_X1 port map( A => n4034, Z => n13928);
   U1402 : BUF_X1 port map( A => n4023, Z => n13955);
   U1403 : BUF_X1 port map( A => n3997, Z => n14009);
   U1404 : BUF_X1 port map( A => n4058, Z => n13886);
   U1405 : BUF_X1 port map( A => n3995, Z => n14015);
   U1406 : BUF_X1 port map( A => n4032, Z => n13934);
   U1407 : BUF_X1 port map( A => n4056, Z => n13892);
   U1408 : BUF_X1 port map( A => n4021, Z => n13961);
   U1409 : BUF_X1 port map( A => n2852, Z => n14136);
   U1410 : BUF_X1 port map( A => n14966, Z => n14965);
   U1411 : INV_X1 port map( A => n3312, ZN => n2566);
   U1412 : INV_X1 port map( A => n4037, ZN => n2542);
   U1413 : NAND2_X1 port map( A1 => n2710, A2 => n2693, ZN => n2768);
   U1414 : NAND2_X1 port map( A1 => n2710, A2 => n2678, ZN => n2756);
   U1415 : NAND2_X1 port map( A1 => n2710, A2 => n2673, ZN => n2752);
   U1416 : NAND2_X1 port map( A1 => n2710, A2 => n2662, ZN => n2743);
   U1417 : NAND2_X1 port map( A1 => n2710, A2 => n2740, ZN => n2738);
   U1418 : NAND2_X1 port map( A1 => n2710, A2 => n2703, ZN => n2776);
   U1419 : NAND2_X1 port map( A1 => n2710, A2 => n2698, ZN => n2772);
   U1420 : NAND2_X1 port map( A1 => n2710, A2 => n2688, ZN => n2764);
   U1421 : NAND2_X1 port map( A1 => n2710, A2 => n2683, ZN => n2760);
   U1422 : NAND2_X1 port map( A1 => n2710, A2 => n2668, ZN => n2747);
   U1423 : INV_X1 port map( A => n3313, ZN => n2565);
   U1424 : INV_X1 port map( A => n4036, ZN => n2541);
   U1425 : BUF_X1 port map( A => n14966, Z => n14962);
   U1426 : NAND2_X1 port map( A1 => n14081, A2 => n14085, ZN => n3956);
   U1427 : NAND2_X1 port map( A1 => n13861, A2 => n13865, ZN => n5277);
   U1428 : BUF_X1 port map( A => n14966, Z => n14963);
   U1429 : BUF_X1 port map( A => n14966, Z => n14964);
   U1430 : NAND2_X1 port map( A1 => n2730, A2 => n2710, ZN => n2728);
   U1431 : NAND2_X1 port map( A1 => n2709, A2 => n2710, ZN => n2706);
   U1432 : NAND2_X1 port map( A1 => n2735, A2 => n2710, ZN => n2733);
   U1433 : NAND2_X1 port map( A1 => n2725, A2 => n2710, ZN => n2723);
   U1434 : NAND2_X1 port map( A1 => n2720, A2 => n2710, ZN => n2718);
   U1435 : NAND2_X1 port map( A1 => n2715, A2 => n2710, ZN => n2713);
   U1436 : AND2_X1 port map( A1 => n5226, A2 => n5189, ZN => n4049);
   U1437 : AND2_X1 port map( A1 => n6547, A2 => n6510, ZN => n5372);
   U1438 : INV_X1 port map( A => n2761, ZN => n2556);
   U1439 : INV_X1 port map( A => n2757, ZN => n2555);
   U1440 : BUF_X1 port map( A => n14948, Z => n14952);
   U1441 : BUF_X1 port map( A => n14966, Z => n14961);
   U1442 : BUF_X1 port map( A => n14966, Z => n14960);
   U1443 : BUF_X1 port map( A => n14966, Z => n14959);
   U1444 : BUF_X1 port map( A => n14947, Z => n14958);
   U1445 : BUF_X1 port map( A => n14951, Z => n14957);
   U1446 : BUF_X1 port map( A => n14961, Z => n14956);
   U1447 : BUF_X1 port map( A => n14948, Z => n14955);
   U1448 : BUF_X1 port map( A => n14960, Z => n14954);
   U1449 : BUF_X1 port map( A => n14947, Z => n14953);
   U1450 : BUF_X1 port map( A => n14961, Z => n14948);
   U1451 : BUF_X1 port map( A => n14960, Z => n14947);
   U1452 : BUF_X1 port map( A => n14959, Z => n14951);
   U1453 : BUF_X1 port map( A => n14952, Z => n14950);
   U1454 : BUF_X1 port map( A => n14958, Z => n14949);
   U1455 : BUF_X1 port map( A => n14275, Z => n14286);
   U1456 : INV_X1 port map( A => n2765, ZN => n2559);
   U1457 : INV_X1 port map( A => n2753, ZN => n2558);
   U1458 : BUF_X1 port map( A => n14273, Z => n14278);
   U1459 : BUF_X1 port map( A => n14273, Z => n14279);
   U1460 : BUF_X1 port map( A => n14273, Z => n14280);
   U1461 : BUF_X1 port map( A => n14274, Z => n14281);
   U1462 : BUF_X1 port map( A => n14274, Z => n14282);
   U1463 : BUF_X1 port map( A => n14274, Z => n14283);
   U1464 : BUF_X1 port map( A => n14275, Z => n14284);
   U1465 : BUF_X1 port map( A => n14275, Z => n14285);
   U1466 : OAI222_X1 port map( A1 => n14239, A2 => n55, B1 => n14236, B2 => n39
                           , C1 => n14233, C2 => n47, ZN => n2800);
   U1467 : OAI222_X1 port map( A1 => n14185, A2 => n162, B1 => n14182, B2 => 
                           n178, C1 => n14179, C2 => n170, ZN => n2826);
   U1468 : OAI222_X1 port map( A1 => n14239, A2 => n54, B1 => n14236, B2 => n38
                           , C1 => n14233, C2 => n46, ZN => n2889);
   U1469 : OAI222_X1 port map( A1 => n14185, A2 => n161, B1 => n14182, B2 => 
                           n177, C1 => n14179, C2 => n169, ZN => n2897);
   U1470 : OAI222_X1 port map( A1 => n14239, A2 => n53, B1 => n14236, B2 => n37
                           , C1 => n14233, C2 => n45, ZN => n2926);
   U1471 : OAI222_X1 port map( A1 => n14185, A2 => n160, B1 => n14182, B2 => 
                           n176, C1 => n14179, C2 => n168, ZN => n2934);
   U1472 : OAI222_X1 port map( A1 => n14239, A2 => n52, B1 => n14236, B2 => n36
                           , C1 => n14233, C2 => n44, ZN => n2963);
   U1473 : OAI222_X1 port map( A1 => n14185, A2 => n159, B1 => n14182, B2 => 
                           n175, C1 => n14179, C2 => n167, ZN => n2971);
   U1474 : OAI222_X1 port map( A1 => n14239, A2 => n51, B1 => n14236, B2 => n35
                           , C1 => n14233, C2 => n43, ZN => n3000);
   U1475 : OAI222_X1 port map( A1 => n14185, A2 => n158, B1 => n14182, B2 => 
                           n174, C1 => n14179, C2 => n166, ZN => n3008);
   U1476 : OAI222_X1 port map( A1 => n14239, A2 => n50, B1 => n14236, B2 => n34
                           , C1 => n14233, C2 => n42, ZN => n3037);
   U1477 : OAI222_X1 port map( A1 => n14185, A2 => n157, B1 => n14182, B2 => 
                           n173, C1 => n14179, C2 => n165, ZN => n3045);
   U1478 : OAI222_X1 port map( A1 => n14239, A2 => n49, B1 => n14236, B2 => n33
                           , C1 => n14233, C2 => n41, ZN => n3074);
   U1479 : OAI222_X1 port map( A1 => n14185, A2 => n156, B1 => n14182, B2 => 
                           n172, C1 => n14179, C2 => n164, ZN => n3082);
   U1480 : OAI222_X1 port map( A1 => n14239, A2 => n1129, B1 => n14236, B2 => 
                           n738, C1 => n14233, C2 => n771, ZN => n3111);
   U1481 : OAI222_X1 port map( A1 => n14185, A2 => n1375, B1 => n14182, B2 => 
                           n1423, C1 => n14179, C2 => n1399, ZN => n3119);
   U1482 : OAI222_X1 port map( A1 => n310, A2 => n14042, B1 => n326, B2 => 
                           n14039, C1 => n318, C2 => n14036, ZN => n4262);
   U1483 : OAI222_X1 port map( A1 => n315, A2 => n13822, B1 => n331, B2 => 
                           n13819, C1 => n323, C2 => n13816, ZN => n5398);
   U1484 : OAI222_X1 port map( A1 => n313, A2 => n13822, B1 => n329, B2 => 
                           n13819, C1 => n321, C2 => n13816, ZN => n5472);
   U1485 : OAI222_X1 port map( A1 => n312, A2 => n13822, B1 => n328, B2 => 
                           n13819, C1 => n320, C2 => n13816, ZN => n5509);
   U1486 : OAI222_X1 port map( A1 => n311, A2 => n13822, B1 => n327, B2 => 
                           n13819, C1 => n319, C2 => n13816, ZN => n5546);
   U1487 : OAI222_X1 port map( A1 => n310, A2 => n13822, B1 => n326, B2 => 
                           n13819, C1 => n318, C2 => n13816, ZN => n5583);
   U1488 : OAI222_X1 port map( A1 => n315, A2 => n14042, B1 => n331, B2 => 
                           n14039, C1 => n323, C2 => n14036, ZN => n4075);
   U1489 : OAI222_X1 port map( A1 => n314, A2 => n14042, B1 => n330, B2 => 
                           n14039, C1 => n322, C2 => n14036, ZN => n4114);
   U1490 : OAI222_X1 port map( A1 => n314, A2 => n13822, B1 => n330, B2 => 
                           n13819, C1 => n322, C2 => n13816, ZN => n5435);
   U1491 : OAI222_X1 port map( A1 => n313, A2 => n14042, B1 => n329, B2 => 
                           n14039, C1 => n321, C2 => n14036, ZN => n4151);
   U1492 : OAI222_X1 port map( A1 => n312, A2 => n14042, B1 => n328, B2 => 
                           n14039, C1 => n320, C2 => n14036, ZN => n4188);
   U1493 : OAI222_X1 port map( A1 => n311, A2 => n14042, B1 => n327, B2 => 
                           n14039, C1 => n319, C2 => n14036, ZN => n4225);
   U1494 : OAI222_X1 port map( A1 => n309, A2 => n14042, B1 => n325, B2 => 
                           n14039, C1 => n317, C2 => n14036, ZN => n4299);
   U1495 : OAI222_X1 port map( A1 => n309, A2 => n13822, B1 => n325, B2 => 
                           n13819, C1 => n317, C2 => n13816, ZN => n5620);
   U1496 : OAI222_X1 port map( A1 => n2497, A2 => n13986, B1 => n1997, B2 => 
                           n13983, C1 => n2431, C2 => n13980, ZN => n4788);
   U1497 : OAI222_X1 port map( A1 => n2497, A2 => n13766, B1 => n1997, B2 => 
                           n13763, C1 => n2431, C2 => n13760, ZN => n6109);
   U1498 : OAI222_X1 port map( A1 => n2519, A2 => n13987, B1 => n1998, B2 => 
                           n13984, C1 => n2432, C2 => n13981, ZN => n4751);
   U1499 : OAI222_X1 port map( A1 => n2519, A2 => n13767, B1 => n1998, B2 => 
                           n13764, C1 => n2432, C2 => n13761, ZN => n6072);
   U1500 : OAI222_X1 port map( A1 => n964, A2 => n14041, B1 => n1012, B2 => 
                           n14038, C1 => n531, C2 => n14035, ZN => n4336);
   U1501 : OAI222_X1 port map( A1 => n964, A2 => n13821, B1 => n1012, B2 => 
                           n13818, C1 => n531, C2 => n13815, ZN => n5657);
   U1502 : OAI222_X1 port map( A1 => n960, A2 => n14041, B1 => n1011, B2 => 
                           n14038, C1 => n530, C2 => n14035, ZN => n4373);
   U1503 : OAI222_X1 port map( A1 => n960, A2 => n13821, B1 => n1011, B2 => 
                           n13818, C1 => n530, C2 => n13815, ZN => n5694);
   U1504 : OAI222_X1 port map( A1 => n958, A2 => n14041, B1 => n1010, B2 => 
                           n14038, C1 => n529, C2 => n14035, ZN => n4410);
   U1505 : OAI222_X1 port map( A1 => n958, A2 => n13821, B1 => n1010, B2 => 
                           n13818, C1 => n529, C2 => n13815, ZN => n5731);
   U1506 : OAI222_X1 port map( A1 => n954, A2 => n14041, B1 => n1009, B2 => 
                           n14038, C1 => n528, C2 => n14035, ZN => n4447);
   U1507 : OAI222_X1 port map( A1 => n954, A2 => n13821, B1 => n1009, B2 => 
                           n13818, C1 => n528, C2 => n13815, ZN => n5768);
   U1508 : OAI222_X1 port map( A1 => n952, A2 => n14041, B1 => n1008, B2 => 
                           n14038, C1 => n527, C2 => n14035, ZN => n4484);
   U1509 : OAI222_X1 port map( A1 => n952, A2 => n13821, B1 => n1008, B2 => 
                           n13818, C1 => n527, C2 => n13815, ZN => n5805);
   U1510 : OAI222_X1 port map( A1 => n948, A2 => n14041, B1 => n1007, B2 => 
                           n14038, C1 => n526, C2 => n14035, ZN => n4521);
   U1511 : OAI222_X1 port map( A1 => n948, A2 => n13821, B1 => n1007, B2 => 
                           n13818, C1 => n526, C2 => n13815, ZN => n5842);
   U1512 : OAI222_X1 port map( A1 => n946, A2 => n14041, B1 => n1006, B2 => 
                           n14038, C1 => n525, C2 => n14035, ZN => n4558);
   U1513 : OAI222_X1 port map( A1 => n946, A2 => n13821, B1 => n1006, B2 => 
                           n13818, C1 => n525, C2 => n13815, ZN => n5879);
   U1514 : OAI222_X1 port map( A1 => n942, A2 => n14041, B1 => n1005, B2 => 
                           n14038, C1 => n524, C2 => n14035, ZN => n4595);
   U1515 : OAI222_X1 port map( A1 => n942, A2 => n13821, B1 => n1005, B2 => 
                           n13818, C1 => n524, C2 => n13815, ZN => n5916);
   U1516 : OAI222_X1 port map( A1 => n940, A2 => n14041, B1 => n1004, B2 => 
                           n14038, C1 => n523, C2 => n14035, ZN => n4632);
   U1517 : OAI222_X1 port map( A1 => n940, A2 => n13821, B1 => n1004, B2 => 
                           n13818, C1 => n523, C2 => n13815, ZN => n5953);
   U1518 : OAI222_X1 port map( A1 => n936, A2 => n14041, B1 => n1003, B2 => 
                           n14038, C1 => n522, C2 => n14035, ZN => n4669);
   U1519 : OAI222_X1 port map( A1 => n936, A2 => n13821, B1 => n1003, B2 => 
                           n13818, C1 => n522, C2 => n13815, ZN => n5990);
   U1520 : AOI221_X1 port map( B1 => n13854, B2 => n424, C1 => n13851, C2 => 
                           n448, A => n6062, ZN => n6061);
   U1521 : OAI222_X1 port map( A1 => n2481, A2 => n13848, B1 => n2419, B2 => 
                           n13845, C1 => n2483, C2 => n13842, ZN => n6062);
   U1522 : OAI222_X1 port map( A1 => n14237, A2 => n56, B1 => n14234, B2 => n40
                           , C1 => n14231, C2 => n48, ZN => n6571);
   U1523 : OAI222_X1 port map( A1 => n14183, A2 => n163, B1 => n14180, B2 => 
                           n179, C1 => n14177, C2 => n171, ZN => n6584);
   U1524 : OAI222_X1 port map( A1 => n14238, A2 => n1128, B1 => n14235, B2 => 
                           n737, C1 => n14232, C2 => n769, ZN => n3148);
   U1525 : OAI222_X1 port map( A1 => n14184, A2 => n1374, B1 => n14181, B2 => 
                           n1422, C1 => n14178, C2 => n1398, ZN => n3156);
   U1526 : OAI222_X1 port map( A1 => n14238, A2 => n1127, B1 => n14235, B2 => 
                           n733, C1 => n14232, C2 => n768, ZN => n3185);
   U1527 : OAI222_X1 port map( A1 => n14184, A2 => n1373, B1 => n14181, B2 => 
                           n1421, C1 => n14178, C2 => n1397, ZN => n3193);
   U1528 : OAI222_X1 port map( A1 => n14238, A2 => n1126, B1 => n14235, B2 => 
                           n732, C1 => n14232, C2 => n767, ZN => n3222);
   U1529 : OAI222_X1 port map( A1 => n14184, A2 => n1372, B1 => n14181, B2 => 
                           n1420, C1 => n14178, C2 => n1396, ZN => n3230);
   U1530 : OAI222_X1 port map( A1 => n14238, A2 => n1125, B1 => n14235, B2 => 
                           n730, C1 => n14232, C2 => n766, ZN => n3259);
   U1531 : OAI222_X1 port map( A1 => n14184, A2 => n1371, B1 => n14181, B2 => 
                           n1419, C1 => n14178, C2 => n1395, ZN => n3267);
   U1532 : OAI222_X1 port map( A1 => n14238, A2 => n1124, B1 => n14235, B2 => 
                           n729, C1 => n14232, C2 => n765, ZN => n3296);
   U1533 : OAI222_X1 port map( A1 => n14184, A2 => n1370, B1 => n14181, B2 => 
                           n1418, C1 => n14178, C2 => n1394, ZN => n3304);
   U1534 : OAI222_X1 port map( A1 => n14238, A2 => n1123, B1 => n14235, B2 => 
                           n728, C1 => n14232, C2 => n764, ZN => n3335);
   U1535 : OAI222_X1 port map( A1 => n14184, A2 => n1369, B1 => n14181, B2 => 
                           n1417, C1 => n14178, C2 => n1393, ZN => n3343);
   U1536 : OAI222_X1 port map( A1 => n14238, A2 => n1122, B1 => n14235, B2 => 
                           n726, C1 => n14232, C2 => n760, ZN => n3372);
   U1537 : OAI222_X1 port map( A1 => n14184, A2 => n1368, B1 => n14181, B2 => 
                           n1416, C1 => n14178, C2 => n1392, ZN => n3380);
   U1538 : OAI222_X1 port map( A1 => n14238, A2 => n1121, B1 => n14235, B2 => 
                           n725, C1 => n14232, C2 => n759, ZN => n3409);
   U1539 : OAI222_X1 port map( A1 => n14184, A2 => n1367, B1 => n14181, B2 => 
                           n1415, C1 => n14178, C2 => n1391, ZN => n3417);
   U1540 : OAI222_X1 port map( A1 => n14238, A2 => n1120, B1 => n14235, B2 => 
                           n724, C1 => n14232, C2 => n758, ZN => n3446);
   U1541 : OAI222_X1 port map( A1 => n14184, A2 => n1366, B1 => n14181, B2 => 
                           n1414, C1 => n14178, C2 => n1390, ZN => n3454);
   U1542 : OAI222_X1 port map( A1 => n14238, A2 => n1119, B1 => n14235, B2 => 
                           n723, C1 => n14232, C2 => n757, ZN => n3483);
   U1543 : OAI222_X1 port map( A1 => n14184, A2 => n1365, B1 => n14181, B2 => 
                           n1413, C1 => n14178, C2 => n1389, ZN => n3491);
   U1544 : OAI222_X1 port map( A1 => n14238, A2 => n1118, B1 => n14235, B2 => 
                           n722, C1 => n14232, C2 => n755, ZN => n3520);
   U1545 : OAI222_X1 port map( A1 => n14184, A2 => n1364, B1 => n14181, B2 => 
                           n1412, C1 => n14178, C2 => n1388, ZN => n3528);
   U1546 : OAI222_X1 port map( A1 => n14238, A2 => n1117, B1 => n14235, B2 => 
                           n721, C1 => n14232, C2 => n751, ZN => n3557);
   U1547 : OAI222_X1 port map( A1 => n14184, A2 => n1363, B1 => n14181, B2 => 
                           n1411, C1 => n14178, C2 => n1387, ZN => n3565);
   U1548 : OAI222_X1 port map( A1 => n14237, A2 => n1116, B1 => n14234, B2 => 
                           n720, C1 => n14231, C2 => n750, ZN => n3594);
   U1549 : OAI222_X1 port map( A1 => n14183, A2 => n1362, B1 => n14180, B2 => 
                           n1410, C1 => n14177, C2 => n1386, ZN => n3602);
   U1550 : OAI222_X1 port map( A1 => n14237, A2 => n1115, B1 => n14234, B2 => 
                           n719, C1 => n14231, C2 => n749, ZN => n3631);
   U1551 : OAI222_X1 port map( A1 => n14183, A2 => n1361, B1 => n14180, B2 => 
                           n1409, C1 => n14177, C2 => n1385, ZN => n3639);
   U1552 : OAI222_X1 port map( A1 => n14237, A2 => n1114, B1 => n14234, B2 => 
                           n718, C1 => n14231, C2 => n748, ZN => n3668);
   U1553 : OAI222_X1 port map( A1 => n14183, A2 => n1360, B1 => n14180, B2 => 
                           n1408, C1 => n14177, C2 => n1384, ZN => n3676);
   U1554 : OAI222_X1 port map( A1 => n14237, A2 => n1113, B1 => n14234, B2 => 
                           n717, C1 => n14231, C2 => n747, ZN => n3705);
   U1555 : OAI222_X1 port map( A1 => n14183, A2 => n1359, B1 => n14180, B2 => 
                           n1407, C1 => n14177, C2 => n1383, ZN => n3713);
   U1556 : OAI222_X1 port map( A1 => n14237, A2 => n1112, B1 => n14234, B2 => 
                           n716, C1 => n14231, C2 => n746, ZN => n3742);
   U1557 : OAI222_X1 port map( A1 => n14183, A2 => n1358, B1 => n14180, B2 => 
                           n1406, C1 => n14177, C2 => n1382, ZN => n3750);
   U1558 : OAI222_X1 port map( A1 => n14237, A2 => n1111, B1 => n14234, B2 => 
                           n715, C1 => n14231, C2 => n745, ZN => n3779);
   U1559 : OAI222_X1 port map( A1 => n14183, A2 => n1357, B1 => n14180, B2 => 
                           n1405, C1 => n14177, C2 => n1381, ZN => n3787);
   U1560 : OAI222_X1 port map( A1 => n14237, A2 => n1110, B1 => n14234, B2 => 
                           n714, C1 => n14231, C2 => n744, ZN => n3816);
   U1561 : OAI222_X1 port map( A1 => n14183, A2 => n1356, B1 => n14180, B2 => 
                           n1404, C1 => n14177, C2 => n1380, ZN => n3824);
   U1562 : OAI222_X1 port map( A1 => n14237, A2 => n1109, B1 => n14234, B2 => 
                           n713, C1 => n14231, C2 => n742, ZN => n3853);
   U1563 : OAI222_X1 port map( A1 => n14183, A2 => n1355, B1 => n14180, B2 => 
                           n1403, C1 => n14177, C2 => n1379, ZN => n3861);
   U1564 : OAI222_X1 port map( A1 => n14237, A2 => n1108, B1 => n14234, B2 => 
                           n712, C1 => n14231, C2 => n741, ZN => n3890);
   U1565 : OAI222_X1 port map( A1 => n14183, A2 => n1354, B1 => n14180, B2 => 
                           n1402, C1 => n14177, C2 => n1378, ZN => n3898);
   U1566 : OAI222_X1 port map( A1 => n14237, A2 => n1107, B1 => n14234, B2 => 
                           n711, C1 => n14231, C2 => n740, ZN => n3927);
   U1567 : OAI222_X1 port map( A1 => n14183, A2 => n1353, B1 => n14180, B2 => 
                           n1401, C1 => n14177, C2 => n1377, ZN => n3935);
   U1568 : OAI222_X1 port map( A1 => n14237, A2 => n1106, B1 => n14234, B2 => 
                           n710, C1 => n14231, C2 => n739, ZN => n5249);
   U1569 : OAI222_X1 port map( A1 => n14183, A2 => n1352, B1 => n14180, B2 => 
                           n1400, C1 => n14177, C2 => n1376, ZN => n5257);
   U1570 : AOI221_X1 port map( B1 => n14074, B2 => n424, C1 => n14071, C2 => 
                           n448, A => n4741, ZN => n4740);
   U1571 : OAI222_X1 port map( A1 => n2481, A2 => n14068, B1 => n2419, B2 => 
                           n14065, C1 => n2483, C2 => n14062, ZN => n4741);
   U1572 : OAI222_X1 port map( A1 => n14716, A2 => n2432, B1 => n14708, B2 => 
                           n14568, C1 => n14821, C2 => n14705, ZN => n10009);
   U1573 : OAI222_X1 port map( A1 => n14716, A2 => n2431, B1 => n14708, B2 => 
                           n14562, C1 => n14815, C2 => n14705, ZN => n10008);
   U1574 : OAI222_X1 port map( A1 => n14891, A2 => n13395, B1 => n2137, B2 => 
                           n13392, C1 => n14633, C2 => n13390, ZN => n10628);
   U1575 : OAI222_X1 port map( A1 => n14889, A2 => n13557, B1 => n2028, B2 => 
                           n13554, C1 => n14631, C2 => n13552, ZN => n11204);
   U1576 : OAI222_X1 port map( A1 => n14940, A2 => n13306, B1 => n1783, B2 => 
                           n13303, C1 => n14681, C2 => n13300, ZN => n10316);
   U1577 : OAI222_X1 port map( A1 => n14940, A2 => n13315, B1 => n1782, B2 => 
                           n13312, C1 => n14682, C2 => n13309, ZN => n10348);
   U1578 : OAI222_X1 port map( A1 => n14939, A2 => n13387, B1 => n1758, B2 => 
                           n13384, C1 => n14681, C2 => n13381, ZN => n10604);
   U1579 : OAI222_X1 port map( A1 => n14939, A2 => n13396, B1 => n1757, B2 => 
                           n13393, C1 => n14681, C2 => n13390, ZN => n10636);
   U1580 : OAI222_X1 port map( A1 => n14933, A2 => n13396, B1 => n1756, B2 => 
                           n13393, C1 => n14675, C2 => n13390, ZN => n10635);
   U1581 : OAI222_X1 port map( A1 => n14921, A2 => n13396, B1 => n1755, B2 => 
                           n13393, C1 => n14663, C2 => n13390, ZN => n10633);
   U1582 : OAI222_X1 port map( A1 => n14915, A2 => n13396, B1 => n1754, B2 => 
                           n13393, C1 => n14657, C2 => n13390, ZN => n10632);
   U1583 : OAI222_X1 port map( A1 => n14909, A2 => n13396, B1 => n1753, B2 => 
                           n13393, C1 => n14651, C2 => n13390, ZN => n10631);
   U1584 : OAI222_X1 port map( A1 => n14903, A2 => n13396, B1 => n1752, B2 => 
                           n13393, C1 => n14645, C2 => n13390, ZN => n10630);
   U1585 : OAI222_X1 port map( A1 => n14897, A2 => n13396, B1 => n1751, B2 => 
                           n13393, C1 => n14639, C2 => n13390, ZN => n10629);
   U1586 : OAI222_X1 port map( A1 => n14938, A2 => n13468, B1 => n1742, B2 => 
                           n13465, C1 => n14680, C2 => n13462, ZN => n10892);
   U1587 : OAI222_X1 port map( A1 => n14938, A2 => n13477, B1 => n1741, B2 => 
                           n13474, C1 => n14680, C2 => n13471, ZN => n10924);
   U1588 : OAI222_X1 port map( A1 => n14938, A2 => n13549, B1 => n1732, B2 => 
                           n13546, C1 => n14679, C2 => n13543, ZN => n11180);
   U1589 : OAI222_X1 port map( A1 => n14937, A2 => n13558, B1 => n1731, B2 => 
                           n13555, C1 => n14679, C2 => n13552, ZN => n11212);
   U1590 : OAI222_X1 port map( A1 => n14931, A2 => n13558, B1 => n1730, B2 => 
                           n13555, C1 => n14673, C2 => n13552, ZN => n11211);
   U1591 : OAI222_X1 port map( A1 => n14919, A2 => n13558, B1 => n1729, B2 => 
                           n13555, C1 => n14661, C2 => n13552, ZN => n11209);
   U1592 : OAI222_X1 port map( A1 => n14913, A2 => n13558, B1 => n1728, B2 => 
                           n13555, C1 => n14655, C2 => n13552, ZN => n11208);
   U1593 : OAI222_X1 port map( A1 => n14907, A2 => n13558, B1 => n1727, B2 => 
                           n13555, C1 => n14649, C2 => n13552, ZN => n11207);
   U1594 : OAI222_X1 port map( A1 => n14901, A2 => n13558, B1 => n1726, B2 => 
                           n13555, C1 => n14643, C2 => n13552, ZN => n11206);
   U1595 : OAI222_X1 port map( A1 => n14895, A2 => n13558, B1 => n1725, B2 => 
                           n13555, C1 => n14637, C2 => n13552, ZN => n11205);
   U1596 : OAI222_X1 port map( A1 => n14887, A2 => n14444, B1 => n14440, B2 => 
                           n1706, C1 => n14629, C2 => n14439, ZN => n9732);
   U1597 : OAI222_X1 port map( A1 => n14887, A2 => n14462, B1 => n14459, B2 => 
                           n1691, C1 => n14629, C2 => n14457, ZN => n9796);
   U1598 : OAI222_X1 port map( A1 => n14887, A2 => n14471, B1 => n14467, B2 => 
                           n1670, C1 => n14629, C2 => n14466, ZN => n9828);
   U1599 : OAI222_X1 port map( A1 => n14892, A2 => n13305, B1 => n1574, B2 => 
                           n13302, C1 => n14633, C2 => n13300, ZN => n10308);
   U1600 : OAI222_X1 port map( A1 => n14892, A2 => n13323, B1 => n1559, B2 => 
                           n13320, C1 => n14634, C2 => n13318, ZN => n10372);
   U1601 : OAI222_X1 port map( A1 => n14892, A2 => n13332, B1 => n1535, B2 => 
                           n13329, C1 => n14633, C2 => n13327, ZN => n10404);
   U1602 : OAI222_X1 port map( A1 => n14891, A2 => n13386, B1 => n1462, B2 => 
                           n13383, C1 => n14633, C2 => n13381, ZN => n10596);
   U1603 : OAI222_X1 port map( A1 => n14891, A2 => n13413, B1 => n1423, B2 => 
                           n13410, C1 => n14633, C2 => n13408, ZN => n10692);
   U1604 : OAI222_X1 port map( A1 => n14891, A2 => n13422, B1 => n1399, B2 => 
                           n13419, C1 => n14633, C2 => n13417, ZN => n10724);
   U1605 : OAI222_X1 port map( A1 => n14890, A2 => n13467, B1 => n1303, B2 => 
                           n13464, C1 => n14632, C2 => n13462, ZN => n10884);
   U1606 : OAI222_X1 port map( A1 => n14890, A2 => n13485, B1 => n1288, B2 => 
                           n13482, C1 => n14632, C2 => n13480, ZN => n10948);
   U1607 : OAI222_X1 port map( A1 => n14890, A2 => n13494, B1 => n1264, B2 => 
                           n13491, C1 => n14632, C2 => n13489, ZN => n10980);
   U1608 : OAI222_X1 port map( A1 => n14890, A2 => n13503, B1 => n1240, B2 => 
                           n13500, C1 => n14632, C2 => n13498, ZN => n11012);
   U1609 : OAI222_X1 port map( A1 => n14890, A2 => n13512, B1 => n1216, B2 => 
                           n13509, C1 => n14632, C2 => n13507, ZN => n11044);
   U1610 : OAI222_X1 port map( A1 => n14890, A2 => n13548, B1 => n1144, B2 => 
                           n13545, C1 => n14631, C2 => n13543, ZN => n11172);
   U1611 : OAI222_X1 port map( A1 => n14889, A2 => n13566, B1 => n1129, B2 => 
                           n13563, C1 => n14631, C2 => n13561, ZN => n11236);
   U1612 : OAI222_X1 port map( A1 => n14888, A2 => n14352, B1 => n14348, B2 => 
                           n1012, C1 => n14631, C2 => n14347, ZN => n9412);
   U1613 : OAI222_X1 port map( A1 => n14888, A2 => n14381, B1 => n14377, B2 => 
                           n813, C1 => n14630, C2 => n14376, ZN => n9508);
   U1614 : OAI222_X1 port map( A1 => n14889, A2 => n13584, B1 => n738, B2 => 
                           n13581, C1 => n14631, C2 => n13579, ZN => n11300);
   U1615 : OAI222_X1 port map( A1 => n14889, A2 => n13593, B1 => n709, B2 => 
                           n13590, C1 => n14631, C2 => n13588, ZN => n11332);
   U1616 : OAI222_X1 port map( A1 => n14889, A2 => n13602, B1 => n685, B2 => 
                           n13599, C1 => n14631, C2 => n13597, ZN => n11364);
   U1617 : OAI222_X1 port map( A1 => n14889, A2 => n13611, B1 => n661, B2 => 
                           n13608, C1 => n14631, C2 => n13606, ZN => n11396);
   U1618 : OAI222_X1 port map( A1 => n14889, A2 => n13629, B1 => n637, B2 => 
                           n13626, C1 => n14631, C2 => n13624, ZN => n11460);
   U1619 : OAI222_X1 port map( A1 => n14889, A2 => n14294, B1 => n14290, B2 => 
                           n627, C1 => n14630, C2 => n14289, ZN => n9213);
   U1620 : OAI222_X1 port map( A1 => n14889, A2 => n14305, B1 => n14301, B2 => 
                           n603, C1 => n14630, C2 => n14300, ZN => n9252);
   U1621 : OAI222_X1 port map( A1 => n14888, A2 => n14325, B1 => n14322, B2 => 
                           n579, C1 => n14630, C2 => n14320, ZN => n9316);
   U1622 : OAI222_X1 port map( A1 => n14888, A2 => n14363, B1 => n14360, B2 => 
                           n531, C1 => n14630, C2 => n14358, ZN => n9444);
   U1623 : OAI222_X1 port map( A1 => n14888, A2 => n14390, B1 => n14386, B2 => 
                           n507, C1 => n14630, C2 => n14385, ZN => n9540);
   U1624 : OAI222_X1 port map( A1 => n14888, A2 => n14408, B1 => n14405, B2 => 
                           n483, C1 => n14629, C2 => n14403, ZN => n9604);
   U1625 : OAI222_X1 port map( A1 => n14929, A2 => n14445, B1 => n14440, B2 => 
                           n411, C1 => n14671, C2 => n14439, ZN => n9739);
   U1626 : OAI222_X1 port map( A1 => n14923, A2 => n14445, B1 => n14440, B2 => 
                           n410, C1 => n14665, C2 => n14439, ZN => n9738);
   U1627 : OAI222_X1 port map( A1 => n14917, A2 => n14445, B1 => n14440, B2 => 
                           n409, C1 => n14659, C2 => n14439, ZN => n9737);
   U1628 : OAI222_X1 port map( A1 => n14911, A2 => n14445, B1 => n14440, B2 => 
                           n408, C1 => n14653, C2 => n14439, ZN => n9736);
   U1629 : OAI222_X1 port map( A1 => n14905, A2 => n14445, B1 => n14440, B2 => 
                           n407, C1 => n14647, C2 => n14439, ZN => n9735);
   U1630 : OAI222_X1 port map( A1 => n14899, A2 => n14445, B1 => n14440, B2 => 
                           n406, C1 => n14641, C2 => n14439, ZN => n9734);
   U1631 : OAI222_X1 port map( A1 => n14893, A2 => n14445, B1 => n14440, B2 => 
                           n405, C1 => n14635, C2 => n14439, ZN => n9733);
   U1632 : OAI222_X1 port map( A1 => n14935, A2 => n14463, B1 => n14460, B2 => 
                           n404, C1 => n14677, C2 => n14457, ZN => n9804);
   U1633 : OAI222_X1 port map( A1 => n14929, A2 => n14463, B1 => n14460, B2 => 
                           n403, C1 => n14671, C2 => n14457, ZN => n9803);
   U1634 : OAI222_X1 port map( A1 => n14923, A2 => n14463, B1 => n14460, B2 => 
                           n402, C1 => n14665, C2 => n14457, ZN => n9802);
   U1635 : OAI222_X1 port map( A1 => n14917, A2 => n14463, B1 => n14460, B2 => 
                           n401, C1 => n14659, C2 => n14457, ZN => n9801);
   U1636 : OAI222_X1 port map( A1 => n14911, A2 => n14463, B1 => n14460, B2 => 
                           n400, C1 => n14653, C2 => n14457, ZN => n9800);
   U1637 : OAI222_X1 port map( A1 => n14905, A2 => n14463, B1 => n14460, B2 => 
                           n399, C1 => n14647, C2 => n14457, ZN => n9799);
   U1638 : OAI222_X1 port map( A1 => n14899, A2 => n14463, B1 => n14460, B2 => 
                           n398, C1 => n14641, C2 => n14457, ZN => n9798);
   U1639 : OAI222_X1 port map( A1 => n14893, A2 => n14463, B1 => n14460, B2 => 
                           n397, C1 => n14635, C2 => n14457, ZN => n9797);
   U1640 : OAI222_X1 port map( A1 => n14935, A2 => n14472, B1 => n14468, B2 => 
                           n396, C1 => n14677, C2 => n14466, ZN => n9836);
   U1641 : OAI222_X1 port map( A1 => n14929, A2 => n14472, B1 => n14467, B2 => 
                           n395, C1 => n14671, C2 => n14466, ZN => n9835);
   U1642 : OAI222_X1 port map( A1 => n14923, A2 => n14472, B1 => n14467, B2 => 
                           n394, C1 => n14665, C2 => n14466, ZN => n9834);
   U1643 : OAI222_X1 port map( A1 => n14917, A2 => n14472, B1 => n14467, B2 => 
                           n393, C1 => n14659, C2 => n14466, ZN => n9833);
   U1644 : OAI222_X1 port map( A1 => n14911, A2 => n14472, B1 => n14467, B2 => 
                           n392, C1 => n14653, C2 => n14466, ZN => n9832);
   U1645 : OAI222_X1 port map( A1 => n14905, A2 => n14472, B1 => n14467, B2 => 
                           n391, C1 => n14647, C2 => n14466, ZN => n9831);
   U1646 : OAI222_X1 port map( A1 => n14899, A2 => n14472, B1 => n14467, B2 => 
                           n390, C1 => n14641, C2 => n14466, ZN => n9830);
   U1647 : OAI222_X1 port map( A1 => n14893, A2 => n14472, B1 => n14467, B2 => 
                           n389, C1 => n14635, C2 => n14466, ZN => n9829);
   U1648 : OAI222_X1 port map( A1 => n14937, A2 => n14295, B1 => n14291, B2 => 
                           n372, C1 => n14678, C2 => n14289, ZN => n9228);
   U1649 : OAI222_X1 port map( A1 => n14931, A2 => n14295, B1 => n14290, B2 => 
                           n371, C1 => n14672, C2 => n14289, ZN => n9227);
   U1650 : OAI222_X1 port map( A1 => n14925, A2 => n14295, B1 => n14290, B2 => 
                           n370, C1 => n14666, C2 => n14289, ZN => n9225);
   U1651 : OAI222_X1 port map( A1 => n14919, A2 => n14295, B1 => n14290, B2 => 
                           n369, C1 => n14660, C2 => n14289, ZN => n9223);
   U1652 : OAI222_X1 port map( A1 => n14913, A2 => n14295, B1 => n14290, B2 => 
                           n368, C1 => n14654, C2 => n14289, ZN => n9221);
   U1653 : OAI222_X1 port map( A1 => n14907, A2 => n14295, B1 => n14290, B2 => 
                           n367, C1 => n14648, C2 => n14289, ZN => n9219);
   U1654 : OAI222_X1 port map( A1 => n14901, A2 => n14295, B1 => n14290, B2 => 
                           n366, C1 => n14642, C2 => n14289, ZN => n9217);
   U1655 : OAI222_X1 port map( A1 => n14895, A2 => n14295, B1 => n14290, B2 => 
                           n365, C1 => n14636, C2 => n14289, ZN => n9215);
   U1656 : OAI222_X1 port map( A1 => n14937, A2 => n14306, B1 => n14302, B2 => 
                           n364, C1 => n14678, C2 => n14300, ZN => n9260);
   U1657 : OAI222_X1 port map( A1 => n14931, A2 => n14306, B1 => n14301, B2 => 
                           n363, C1 => n14672, C2 => n14300, ZN => n9259);
   U1658 : OAI222_X1 port map( A1 => n14925, A2 => n14306, B1 => n14301, B2 => 
                           n362, C1 => n14666, C2 => n14300, ZN => n9258);
   U1659 : OAI222_X1 port map( A1 => n14919, A2 => n14306, B1 => n14301, B2 => 
                           n361, C1 => n14660, C2 => n14300, ZN => n9257);
   U1660 : OAI222_X1 port map( A1 => n14913, A2 => n14306, B1 => n14301, B2 => 
                           n360, C1 => n14654, C2 => n14300, ZN => n9256);
   U1661 : OAI222_X1 port map( A1 => n14907, A2 => n14306, B1 => n14301, B2 => 
                           n359, C1 => n14648, C2 => n14300, ZN => n9255);
   U1662 : OAI222_X1 port map( A1 => n14901, A2 => n14306, B1 => n14301, B2 => 
                           n358, C1 => n14642, C2 => n14300, ZN => n9254);
   U1663 : OAI222_X1 port map( A1 => n14895, A2 => n14306, B1 => n14301, B2 => 
                           n357, C1 => n14636, C2 => n14300, ZN => n9253);
   U1664 : OAI222_X1 port map( A1 => n14936, A2 => n14326, B1 => n14323, B2 => 
                           n356, C1 => n14678, C2 => n14320, ZN => n9324);
   U1665 : OAI222_X1 port map( A1 => n14930, A2 => n14326, B1 => n14323, B2 => 
                           n355, C1 => n14672, C2 => n14320, ZN => n9323);
   U1666 : OAI222_X1 port map( A1 => n14924, A2 => n14326, B1 => n14323, B2 => 
                           n354, C1 => n14666, C2 => n14320, ZN => n9322);
   U1667 : OAI222_X1 port map( A1 => n14918, A2 => n14326, B1 => n14323, B2 => 
                           n353, C1 => n14660, C2 => n14320, ZN => n9321);
   U1668 : OAI222_X1 port map( A1 => n14912, A2 => n14326, B1 => n14323, B2 => 
                           n352, C1 => n14654, C2 => n14320, ZN => n9320);
   U1669 : OAI222_X1 port map( A1 => n14906, A2 => n14326, B1 => n14323, B2 => 
                           n351, C1 => n14648, C2 => n14320, ZN => n9319);
   U1670 : OAI222_X1 port map( A1 => n14900, A2 => n14326, B1 => n14323, B2 => 
                           n350, C1 => n14642, C2 => n14320, ZN => n9318);
   U1671 : OAI222_X1 port map( A1 => n14894, A2 => n14326, B1 => n14323, B2 => 
                           n349, C1 => n14636, C2 => n14320, ZN => n9317);
   U1672 : OAI222_X1 port map( A1 => n14936, A2 => n14353, B1 => n14349, B2 => 
                           n332, C1 => n14679, C2 => n14347, ZN => n9420);
   U1673 : OAI222_X1 port map( A1 => n14930, A2 => n14353, B1 => n14348, B2 => 
                           n331, C1 => n14673, C2 => n14347, ZN => n9419);
   U1674 : OAI222_X1 port map( A1 => n14924, A2 => n14353, B1 => n14348, B2 => 
                           n330, C1 => n14667, C2 => n14347, ZN => n9418);
   U1675 : OAI222_X1 port map( A1 => n14918, A2 => n14353, B1 => n14348, B2 => 
                           n329, C1 => n14661, C2 => n14347, ZN => n9417);
   U1676 : OAI222_X1 port map( A1 => n14912, A2 => n14353, B1 => n14348, B2 => 
                           n328, C1 => n14655, C2 => n14347, ZN => n9416);
   U1677 : OAI222_X1 port map( A1 => n14906, A2 => n14353, B1 => n14348, B2 => 
                           n327, C1 => n14649, C2 => n14347, ZN => n9415);
   U1678 : OAI222_X1 port map( A1 => n14900, A2 => n14353, B1 => n14348, B2 => 
                           n326, C1 => n14643, C2 => n14347, ZN => n9414);
   U1679 : OAI222_X1 port map( A1 => n14894, A2 => n14353, B1 => n14348, B2 => 
                           n325, C1 => n14637, C2 => n14347, ZN => n9413);
   U1680 : OAI222_X1 port map( A1 => n14936, A2 => n14364, B1 => n14361, B2 => 
                           n324, C1 => n14678, C2 => n14358, ZN => n9452);
   U1681 : OAI222_X1 port map( A1 => n14930, A2 => n14364, B1 => n14361, B2 => 
                           n323, C1 => n14672, C2 => n14358, ZN => n9451);
   U1682 : OAI222_X1 port map( A1 => n14924, A2 => n14364, B1 => n14361, B2 => 
                           n322, C1 => n14666, C2 => n14358, ZN => n9450);
   U1683 : OAI222_X1 port map( A1 => n14918, A2 => n14364, B1 => n14361, B2 => 
                           n321, C1 => n14660, C2 => n14358, ZN => n9449);
   U1684 : OAI222_X1 port map( A1 => n14912, A2 => n14364, B1 => n14361, B2 => 
                           n320, C1 => n14654, C2 => n14358, ZN => n9448);
   U1685 : OAI222_X1 port map( A1 => n14906, A2 => n14364, B1 => n14361, B2 => 
                           n319, C1 => n14648, C2 => n14358, ZN => n9447);
   U1686 : OAI222_X1 port map( A1 => n14900, A2 => n14364, B1 => n14361, B2 => 
                           n318, C1 => n14642, C2 => n14358, ZN => n9446);
   U1687 : OAI222_X1 port map( A1 => n14894, A2 => n14364, B1 => n14361, B2 => 
                           n317, C1 => n14636, C2 => n14358, ZN => n9445);
   U1688 : OAI222_X1 port map( A1 => n14936, A2 => n14382, B1 => n14378, B2 => 
                           n308, C1 => n14678, C2 => n14376, ZN => n9516);
   U1689 : OAI222_X1 port map( A1 => n14930, A2 => n14382, B1 => n14377, B2 => 
                           n307, C1 => n14672, C2 => n14376, ZN => n9515);
   U1690 : OAI222_X1 port map( A1 => n14924, A2 => n14382, B1 => n14377, B2 => 
                           n306, C1 => n14666, C2 => n14376, ZN => n9514);
   U1691 : OAI222_X1 port map( A1 => n14918, A2 => n14382, B1 => n14377, B2 => 
                           n305, C1 => n14660, C2 => n14376, ZN => n9513);
   U1692 : OAI222_X1 port map( A1 => n14912, A2 => n14382, B1 => n14377, B2 => 
                           n304, C1 => n14654, C2 => n14376, ZN => n9512);
   U1693 : OAI222_X1 port map( A1 => n14906, A2 => n14382, B1 => n14377, B2 => 
                           n303, C1 => n14648, C2 => n14376, ZN => n9511);
   U1694 : OAI222_X1 port map( A1 => n14900, A2 => n14382, B1 => n14377, B2 => 
                           n302, C1 => n14642, C2 => n14376, ZN => n9510);
   U1695 : OAI222_X1 port map( A1 => n14894, A2 => n14382, B1 => n14377, B2 => 
                           n301, C1 => n14636, C2 => n14376, ZN => n9509);
   U1696 : OAI222_X1 port map( A1 => n14936, A2 => n14391, B1 => n14387, B2 => 
                           n300, C1 => n14678, C2 => n14385, ZN => n9548);
   U1697 : OAI222_X1 port map( A1 => n14930, A2 => n14391, B1 => n14386, B2 => 
                           n299, C1 => n14672, C2 => n14385, ZN => n9547);
   U1698 : OAI222_X1 port map( A1 => n14924, A2 => n14391, B1 => n14386, B2 => 
                           n298, C1 => n14666, C2 => n14385, ZN => n9546);
   U1699 : OAI222_X1 port map( A1 => n14918, A2 => n14391, B1 => n14386, B2 => 
                           n297, C1 => n14660, C2 => n14385, ZN => n9545);
   U1700 : OAI222_X1 port map( A1 => n14912, A2 => n14391, B1 => n14386, B2 => 
                           n296, C1 => n14654, C2 => n14385, ZN => n9544);
   U1701 : OAI222_X1 port map( A1 => n14906, A2 => n14391, B1 => n14386, B2 => 
                           n295, C1 => n14648, C2 => n14385, ZN => n9543);
   U1702 : OAI222_X1 port map( A1 => n14900, A2 => n14391, B1 => n14386, B2 => 
                           n294, C1 => n14642, C2 => n14385, ZN => n9542);
   U1703 : OAI222_X1 port map( A1 => n14894, A2 => n14391, B1 => n14386, B2 => 
                           n293, C1 => n14636, C2 => n14385, ZN => n9541);
   U1704 : OAI222_X1 port map( A1 => n14936, A2 => n14409, B1 => n14406, B2 => 
                           n292, C1 => n14677, C2 => n14403, ZN => n9612);
   U1705 : OAI222_X1 port map( A1 => n14930, A2 => n14409, B1 => n14406, B2 => 
                           n291, C1 => n14671, C2 => n14403, ZN => n9611);
   U1706 : OAI222_X1 port map( A1 => n14924, A2 => n14409, B1 => n14406, B2 => 
                           n290, C1 => n14665, C2 => n14403, ZN => n9610);
   U1707 : OAI222_X1 port map( A1 => n14918, A2 => n14409, B1 => n14406, B2 => 
                           n289, C1 => n14659, C2 => n14403, ZN => n9609);
   U1708 : OAI222_X1 port map( A1 => n14912, A2 => n14409, B1 => n14406, B2 => 
                           n288, C1 => n14653, C2 => n14403, ZN => n9608);
   U1709 : OAI222_X1 port map( A1 => n14906, A2 => n14409, B1 => n14406, B2 => 
                           n287, C1 => n14647, C2 => n14403, ZN => n9607);
   U1710 : OAI222_X1 port map( A1 => n14900, A2 => n14409, B1 => n14406, B2 => 
                           n286, C1 => n14641, C2 => n14403, ZN => n9606);
   U1711 : OAI222_X1 port map( A1 => n14894, A2 => n14409, B1 => n14406, B2 => 
                           n285, C1 => n14635, C2 => n14403, ZN => n9605);
   U1712 : OAI222_X1 port map( A1 => n14934, A2 => n13306, B1 => n235, B2 => 
                           n13303, C1 => n14675, C2 => n13300, ZN => n10315);
   U1713 : OAI222_X1 port map( A1 => n14928, A2 => n13306, B1 => n234, B2 => 
                           n13303, C1 => n14669, C2 => n13300, ZN => n10314);
   U1714 : OAI222_X1 port map( A1 => n14922, A2 => n13306, B1 => n233, B2 => 
                           n13303, C1 => n14663, C2 => n13300, ZN => n10313);
   U1715 : OAI222_X1 port map( A1 => n14916, A2 => n13306, B1 => n232, B2 => 
                           n13303, C1 => n14657, C2 => n13300, ZN => n10312);
   U1716 : OAI222_X1 port map( A1 => n14910, A2 => n13306, B1 => n231, B2 => 
                           n13303, C1 => n14651, C2 => n13300, ZN => n10311);
   U1717 : OAI222_X1 port map( A1 => n14904, A2 => n13306, B1 => n230, B2 => 
                           n13303, C1 => n14645, C2 => n13300, ZN => n10310);
   U1718 : OAI222_X1 port map( A1 => n14898, A2 => n13306, B1 => n229, B2 => 
                           n13303, C1 => n14639, C2 => n13300, ZN => n10309);
   U1719 : OAI222_X1 port map( A1 => n14940, A2 => n13324, B1 => n228, B2 => 
                           n13321, C1 => n14682, C2 => n13318, ZN => n10380);
   U1720 : OAI222_X1 port map( A1 => n14934, A2 => n13324, B1 => n227, B2 => 
                           n13321, C1 => n14676, C2 => n13318, ZN => n10379);
   U1721 : OAI222_X1 port map( A1 => n14928, A2 => n13324, B1 => n226, B2 => 
                           n13321, C1 => n14670, C2 => n13318, ZN => n10378);
   U1722 : OAI222_X1 port map( A1 => n14922, A2 => n13324, B1 => n225, B2 => 
                           n13321, C1 => n14664, C2 => n13318, ZN => n10377);
   U1723 : OAI222_X1 port map( A1 => n14916, A2 => n13324, B1 => n224, B2 => 
                           n13321, C1 => n14658, C2 => n13318, ZN => n10376);
   U1724 : OAI222_X1 port map( A1 => n14910, A2 => n13324, B1 => n223, B2 => 
                           n13321, C1 => n14652, C2 => n13318, ZN => n10375);
   U1725 : OAI222_X1 port map( A1 => n14904, A2 => n13324, B1 => n222, B2 => 
                           n13321, C1 => n14646, C2 => n13318, ZN => n10374);
   U1726 : OAI222_X1 port map( A1 => n14898, A2 => n13324, B1 => n221, B2 => 
                           n13321, C1 => n14640, C2 => n13318, ZN => n10373);
   U1727 : OAI222_X1 port map( A1 => n14940, A2 => n13333, B1 => n220, B2 => 
                           n13330, C1 => n14681, C2 => n13327, ZN => n10412);
   U1728 : OAI222_X1 port map( A1 => n14934, A2 => n13333, B1 => n219, B2 => 
                           n13330, C1 => n14675, C2 => n13327, ZN => n10411);
   U1729 : OAI222_X1 port map( A1 => n14928, A2 => n13333, B1 => n218, B2 => 
                           n13330, C1 => n14669, C2 => n13327, ZN => n10410);
   U1730 : OAI222_X1 port map( A1 => n14922, A2 => n13333, B1 => n217, B2 => 
                           n13330, C1 => n14663, C2 => n13327, ZN => n10409);
   U1731 : OAI222_X1 port map( A1 => n14916, A2 => n13333, B1 => n216, B2 => 
                           n13330, C1 => n14657, C2 => n13327, ZN => n10408);
   U1732 : OAI222_X1 port map( A1 => n14910, A2 => n13333, B1 => n215, B2 => 
                           n13330, C1 => n14651, C2 => n13327, ZN => n10407);
   U1733 : OAI222_X1 port map( A1 => n14904, A2 => n13333, B1 => n214, B2 => 
                           n13330, C1 => n14645, C2 => n13327, ZN => n10406);
   U1734 : OAI222_X1 port map( A1 => n14898, A2 => n13333, B1 => n213, B2 => 
                           n13330, C1 => n14639, C2 => n13327, ZN => n10405);
   U1735 : OAI222_X1 port map( A1 => n14939, A2 => n13351, B1 => n212, B2 => 
                           n13348, C1 => n14681, C2 => n13345, ZN => n10476);
   U1736 : OAI222_X1 port map( A1 => n14933, A2 => n13387, B1 => n195, B2 => 
                           n13384, C1 => n14675, C2 => n13381, ZN => n10603);
   U1737 : OAI222_X1 port map( A1 => n14927, A2 => n13387, B1 => n194, B2 => 
                           n13384, C1 => n14669, C2 => n13381, ZN => n10602);
   U1738 : OAI222_X1 port map( A1 => n14921, A2 => n13387, B1 => n193, B2 => 
                           n13384, C1 => n14663, C2 => n13381, ZN => n10601);
   U1739 : OAI222_X1 port map( A1 => n14915, A2 => n13387, B1 => n192, B2 => 
                           n13384, C1 => n14657, C2 => n13381, ZN => n10600);
   U1740 : OAI222_X1 port map( A1 => n14909, A2 => n13387, B1 => n191, B2 => 
                           n13384, C1 => n14651, C2 => n13381, ZN => n10599);
   U1741 : OAI222_X1 port map( A1 => n14903, A2 => n13387, B1 => n190, B2 => 
                           n13384, C1 => n14645, C2 => n13381, ZN => n10598);
   U1742 : OAI222_X1 port map( A1 => n14897, A2 => n13387, B1 => n189, B2 => 
                           n13384, C1 => n14639, C2 => n13381, ZN => n10597);
   U1743 : OAI222_X1 port map( A1 => n14927, A2 => n13396, B1 => n188, B2 => 
                           n13393, C1 => n14669, C2 => n13390, ZN => n10634);
   U1744 : OAI222_X1 port map( A1 => n14939, A2 => n13414, B1 => n179, B2 => 
                           n13411, C1 => n14681, C2 => n13408, ZN => n10700);
   U1745 : OAI222_X1 port map( A1 => n14933, A2 => n13414, B1 => n178, B2 => 
                           n13411, C1 => n14675, C2 => n13408, ZN => n10699);
   U1746 : OAI222_X1 port map( A1 => n14927, A2 => n13414, B1 => n177, B2 => 
                           n13411, C1 => n14669, C2 => n13408, ZN => n10698);
   U1747 : OAI222_X1 port map( A1 => n14921, A2 => n13414, B1 => n176, B2 => 
                           n13411, C1 => n14663, C2 => n13408, ZN => n10697);
   U1748 : OAI222_X1 port map( A1 => n14915, A2 => n13414, B1 => n175, B2 => 
                           n13411, C1 => n14657, C2 => n13408, ZN => n10696);
   U1749 : OAI222_X1 port map( A1 => n14909, A2 => n13414, B1 => n174, B2 => 
                           n13411, C1 => n14651, C2 => n13408, ZN => n10695);
   U1750 : OAI222_X1 port map( A1 => n14903, A2 => n13414, B1 => n173, B2 => 
                           n13411, C1 => n14645, C2 => n13408, ZN => n10694);
   U1751 : OAI222_X1 port map( A1 => n14897, A2 => n13414, B1 => n172, B2 => 
                           n13411, C1 => n14639, C2 => n13408, ZN => n10693);
   U1752 : OAI222_X1 port map( A1 => n14939, A2 => n13423, B1 => n171, B2 => 
                           n13420, C1 => n14681, C2 => n13417, ZN => n10732);
   U1753 : OAI222_X1 port map( A1 => n14933, A2 => n13423, B1 => n170, B2 => 
                           n13420, C1 => n14675, C2 => n13417, ZN => n10731);
   U1754 : OAI222_X1 port map( A1 => n14927, A2 => n13423, B1 => n169, B2 => 
                           n13420, C1 => n14669, C2 => n13417, ZN => n10730);
   U1755 : OAI222_X1 port map( A1 => n14921, A2 => n13423, B1 => n168, B2 => 
                           n13420, C1 => n14663, C2 => n13417, ZN => n10729);
   U1756 : OAI222_X1 port map( A1 => n14915, A2 => n13423, B1 => n167, B2 => 
                           n13420, C1 => n14657, C2 => n13417, ZN => n10728);
   U1757 : OAI222_X1 port map( A1 => n14909, A2 => n13423, B1 => n166, B2 => 
                           n13420, C1 => n14651, C2 => n13417, ZN => n10727);
   U1758 : OAI222_X1 port map( A1 => n14903, A2 => n13423, B1 => n165, B2 => 
                           n13420, C1 => n14645, C2 => n13417, ZN => n10726);
   U1759 : OAI222_X1 port map( A1 => n14897, A2 => n13423, B1 => n164, B2 => 
                           n13420, C1 => n14639, C2 => n13417, ZN => n10725);
   U1760 : OAI222_X1 port map( A1 => n14932, A2 => n13468, B1 => n139, B2 => 
                           n13465, C1 => n14674, C2 => n13462, ZN => n10891);
   U1761 : OAI222_X1 port map( A1 => n14926, A2 => n13468, B1 => n138, B2 => 
                           n13465, C1 => n14668, C2 => n13462, ZN => n10890);
   U1762 : OAI222_X1 port map( A1 => n14920, A2 => n13468, B1 => n137, B2 => 
                           n13465, C1 => n14662, C2 => n13462, ZN => n10889);
   U1763 : OAI222_X1 port map( A1 => n14914, A2 => n13468, B1 => n136, B2 => 
                           n13465, C1 => n14656, C2 => n13462, ZN => n10888);
   U1764 : OAI222_X1 port map( A1 => n14908, A2 => n13468, B1 => n135, B2 => 
                           n13465, C1 => n14650, C2 => n13462, ZN => n10887);
   U1765 : OAI222_X1 port map( A1 => n14902, A2 => n13468, B1 => n134, B2 => 
                           n13465, C1 => n14644, C2 => n13462, ZN => n10886);
   U1766 : OAI222_X1 port map( A1 => n14896, A2 => n13468, B1 => n133, B2 => 
                           n13465, C1 => n14638, C2 => n13462, ZN => n10885);
   U1767 : OAI222_X1 port map( A1 => n14926, A2 => n13477, B1 => n132, B2 => 
                           n13474, C1 => n14668, C2 => n13471, ZN => n10922);
   U1768 : OAI222_X1 port map( A1 => n14938, A2 => n13486, B1 => n131, B2 => 
                           n13483, C1 => n14680, C2 => n13480, ZN => n10956);
   U1769 : OAI222_X1 port map( A1 => n14932, A2 => n13486, B1 => n130, B2 => 
                           n13483, C1 => n14674, C2 => n13480, ZN => n10955);
   U1770 : OAI222_X1 port map( A1 => n14926, A2 => n13486, B1 => n129, B2 => 
                           n13483, C1 => n14668, C2 => n13480, ZN => n10954);
   U1771 : OAI222_X1 port map( A1 => n14920, A2 => n13486, B1 => n128, B2 => 
                           n13483, C1 => n14662, C2 => n13480, ZN => n10953);
   U1772 : OAI222_X1 port map( A1 => n14914, A2 => n13486, B1 => n127, B2 => 
                           n13483, C1 => n14656, C2 => n13480, ZN => n10952);
   U1773 : OAI222_X1 port map( A1 => n14908, A2 => n13486, B1 => n126, B2 => 
                           n13483, C1 => n14650, C2 => n13480, ZN => n10951);
   U1774 : OAI222_X1 port map( A1 => n14902, A2 => n13486, B1 => n125, B2 => 
                           n13483, C1 => n14644, C2 => n13480, ZN => n10950);
   U1775 : OAI222_X1 port map( A1 => n14896, A2 => n13486, B1 => n124, B2 => 
                           n13483, C1 => n14638, C2 => n13480, ZN => n10949);
   U1776 : OAI222_X1 port map( A1 => n14938, A2 => n13495, B1 => n123, B2 => 
                           n13492, C1 => n14680, C2 => n13489, ZN => n10988);
   U1777 : OAI222_X1 port map( A1 => n14932, A2 => n13495, B1 => n122, B2 => 
                           n13492, C1 => n14674, C2 => n13489, ZN => n10987);
   U1778 : OAI222_X1 port map( A1 => n14926, A2 => n13495, B1 => n121, B2 => 
                           n13492, C1 => n14668, C2 => n13489, ZN => n10986);
   U1779 : OAI222_X1 port map( A1 => n14920, A2 => n13495, B1 => n120, B2 => 
                           n13492, C1 => n14662, C2 => n13489, ZN => n10985);
   U1780 : OAI222_X1 port map( A1 => n14914, A2 => n13495, B1 => n119, B2 => 
                           n13492, C1 => n14656, C2 => n13489, ZN => n10984);
   U1781 : OAI222_X1 port map( A1 => n14908, A2 => n13495, B1 => n118, B2 => 
                           n13492, C1 => n14650, C2 => n13489, ZN => n10983);
   U1782 : OAI222_X1 port map( A1 => n14902, A2 => n13495, B1 => n117, B2 => 
                           n13492, C1 => n14644, C2 => n13489, ZN => n10982);
   U1783 : OAI222_X1 port map( A1 => n14896, A2 => n13495, B1 => n116, B2 => 
                           n13492, C1 => n14638, C2 => n13489, ZN => n10981);
   U1784 : OAI222_X1 port map( A1 => n14938, A2 => n13504, B1 => n115, B2 => 
                           n13501, C1 => n14680, C2 => n13498, ZN => n11020);
   U1785 : OAI222_X1 port map( A1 => n14932, A2 => n13504, B1 => n114, B2 => 
                           n13501, C1 => n14674, C2 => n13498, ZN => n11019);
   U1786 : OAI222_X1 port map( A1 => n14926, A2 => n13504, B1 => n113, B2 => 
                           n13501, C1 => n14668, C2 => n13498, ZN => n11018);
   U1787 : OAI222_X1 port map( A1 => n14920, A2 => n13504, B1 => n112, B2 => 
                           n13501, C1 => n14662, C2 => n13498, ZN => n11017);
   U1788 : OAI222_X1 port map( A1 => n14914, A2 => n13504, B1 => n111, B2 => 
                           n13501, C1 => n14656, C2 => n13498, ZN => n11016);
   U1789 : OAI222_X1 port map( A1 => n14908, A2 => n13504, B1 => n110, B2 => 
                           n13501, C1 => n14650, C2 => n13498, ZN => n11015);
   U1790 : OAI222_X1 port map( A1 => n14902, A2 => n13504, B1 => n109, B2 => 
                           n13501, C1 => n14644, C2 => n13498, ZN => n11014);
   U1791 : OAI222_X1 port map( A1 => n14896, A2 => n13504, B1 => n108, B2 => 
                           n13501, C1 => n14638, C2 => n13498, ZN => n11013);
   U1792 : OAI222_X1 port map( A1 => n14938, A2 => n13513, B1 => n107, B2 => 
                           n13510, C1 => n14680, C2 => n13507, ZN => n11052);
   U1793 : OAI222_X1 port map( A1 => n14932, A2 => n13513, B1 => n106, B2 => 
                           n13510, C1 => n14674, C2 => n13507, ZN => n11051);
   U1794 : OAI222_X1 port map( A1 => n14926, A2 => n13513, B1 => n105, B2 => 
                           n13510, C1 => n14668, C2 => n13507, ZN => n11050);
   U1795 : OAI222_X1 port map( A1 => n14920, A2 => n13513, B1 => n104, B2 => 
                           n13510, C1 => n14662, C2 => n13507, ZN => n11049);
   U1796 : OAI222_X1 port map( A1 => n14914, A2 => n13513, B1 => n103, B2 => 
                           n13510, C1 => n14656, C2 => n13507, ZN => n11048);
   U1797 : OAI222_X1 port map( A1 => n14908, A2 => n13513, B1 => n102, B2 => 
                           n13510, C1 => n14650, C2 => n13507, ZN => n11047);
   U1798 : OAI222_X1 port map( A1 => n14902, A2 => n13513, B1 => n101, B2 => 
                           n13510, C1 => n14644, C2 => n13507, ZN => n11046);
   U1799 : OAI222_X1 port map( A1 => n14896, A2 => n13513, B1 => n100, B2 => 
                           n13510, C1 => n14638, C2 => n13507, ZN => n11045);
   U1800 : OAI222_X1 port map( A1 => n14932, A2 => n13549, B1 => n64, B2 => 
                           n13546, C1 => n14673, C2 => n13543, ZN => n11179);
   U1801 : OAI222_X1 port map( A1 => n14926, A2 => n13549, B1 => n63, B2 => 
                           n13546, C1 => n14667, C2 => n13543, ZN => n11178);
   U1802 : OAI222_X1 port map( A1 => n14920, A2 => n13549, B1 => n62, B2 => 
                           n13546, C1 => n14661, C2 => n13543, ZN => n11177);
   U1803 : OAI222_X1 port map( A1 => n14914, A2 => n13549, B1 => n61, B2 => 
                           n13546, C1 => n14655, C2 => n13543, ZN => n11176);
   U1804 : OAI222_X1 port map( A1 => n14908, A2 => n13549, B1 => n60, B2 => 
                           n13546, C1 => n14649, C2 => n13543, ZN => n11175);
   U1805 : OAI222_X1 port map( A1 => n14902, A2 => n13549, B1 => n59, B2 => 
                           n13546, C1 => n14643, C2 => n13543, ZN => n11174);
   U1806 : OAI222_X1 port map( A1 => n14896, A2 => n13549, B1 => n58, B2 => 
                           n13546, C1 => n14637, C2 => n13543, ZN => n11173);
   U1807 : OAI222_X1 port map( A1 => n14925, A2 => n13558, B1 => n57, B2 => 
                           n13555, C1 => n14667, C2 => n13552, ZN => n11210);
   U1808 : OAI222_X1 port map( A1 => n14937, A2 => n13567, B1 => n56, B2 => 
                           n13564, C1 => n14679, C2 => n13561, ZN => n11244);
   U1809 : OAI222_X1 port map( A1 => n14931, A2 => n13567, B1 => n55, B2 => 
                           n13564, C1 => n14673, C2 => n13561, ZN => n11243);
   U1810 : OAI222_X1 port map( A1 => n14925, A2 => n13567, B1 => n54, B2 => 
                           n13564, C1 => n14667, C2 => n13561, ZN => n11242);
   U1811 : OAI222_X1 port map( A1 => n14919, A2 => n13567, B1 => n53, B2 => 
                           n13564, C1 => n14661, C2 => n13561, ZN => n11241);
   U1812 : OAI222_X1 port map( A1 => n14913, A2 => n13567, B1 => n52, B2 => 
                           n13564, C1 => n14655, C2 => n13561, ZN => n11240);
   U1813 : OAI222_X1 port map( A1 => n14907, A2 => n13567, B1 => n51, B2 => 
                           n13564, C1 => n14649, C2 => n13561, ZN => n11239);
   U1814 : OAI222_X1 port map( A1 => n14901, A2 => n13567, B1 => n50, B2 => 
                           n13564, C1 => n14643, C2 => n13561, ZN => n11238);
   U1815 : OAI222_X1 port map( A1 => n14895, A2 => n13567, B1 => n49, B2 => 
                           n13564, C1 => n14637, C2 => n13561, ZN => n11237);
   U1816 : OAI222_X1 port map( A1 => n14937, A2 => n13585, B1 => n40, B2 => 
                           n13582, C1 => n14679, C2 => n13579, ZN => n11308);
   U1817 : OAI222_X1 port map( A1 => n14931, A2 => n13585, B1 => n39, B2 => 
                           n13582, C1 => n14673, C2 => n13579, ZN => n11307);
   U1818 : OAI222_X1 port map( A1 => n14925, A2 => n13585, B1 => n38, B2 => 
                           n13582, C1 => n14667, C2 => n13579, ZN => n11306);
   U1819 : OAI222_X1 port map( A1 => n14919, A2 => n13585, B1 => n37, B2 => 
                           n13582, C1 => n14661, C2 => n13579, ZN => n11305);
   U1820 : OAI222_X1 port map( A1 => n14913, A2 => n13585, B1 => n36, B2 => 
                           n13582, C1 => n14655, C2 => n13579, ZN => n11304);
   U1821 : OAI222_X1 port map( A1 => n14907, A2 => n13585, B1 => n35, B2 => 
                           n13582, C1 => n14649, C2 => n13579, ZN => n11303);
   U1822 : OAI222_X1 port map( A1 => n14901, A2 => n13585, B1 => n34, B2 => 
                           n13582, C1 => n14643, C2 => n13579, ZN => n11302);
   U1823 : OAI222_X1 port map( A1 => n14895, A2 => n13585, B1 => n33, B2 => 
                           n13582, C1 => n14637, C2 => n13579, ZN => n11301);
   U1824 : OAI222_X1 port map( A1 => n14937, A2 => n13594, B1 => n32, B2 => 
                           n13591, C1 => n14679, C2 => n13588, ZN => n11340);
   U1825 : OAI222_X1 port map( A1 => n14931, A2 => n13594, B1 => n31, B2 => 
                           n13591, C1 => n14673, C2 => n13588, ZN => n11339);
   U1826 : OAI222_X1 port map( A1 => n14925, A2 => n13594, B1 => n30, B2 => 
                           n13591, C1 => n14667, C2 => n13588, ZN => n11338);
   U1827 : OAI222_X1 port map( A1 => n14919, A2 => n13594, B1 => n29, B2 => 
                           n13591, C1 => n14661, C2 => n13588, ZN => n11337);
   U1828 : OAI222_X1 port map( A1 => n14913, A2 => n13594, B1 => n28, B2 => 
                           n13591, C1 => n14655, C2 => n13588, ZN => n11336);
   U1829 : OAI222_X1 port map( A1 => n14907, A2 => n13594, B1 => n27, B2 => 
                           n13591, C1 => n14649, C2 => n13588, ZN => n11335);
   U1830 : OAI222_X1 port map( A1 => n14901, A2 => n13594, B1 => n26, B2 => 
                           n13591, C1 => n14643, C2 => n13588, ZN => n11334);
   U1831 : OAI222_X1 port map( A1 => n14895, A2 => n13594, B1 => n25, B2 => 
                           n13591, C1 => n14637, C2 => n13588, ZN => n11333);
   U1832 : OAI222_X1 port map( A1 => n14937, A2 => n13603, B1 => n24, B2 => 
                           n13600, C1 => n14679, C2 => n13597, ZN => n11372);
   U1833 : OAI222_X1 port map( A1 => n14931, A2 => n13603, B1 => n23, B2 => 
                           n13600, C1 => n14673, C2 => n13597, ZN => n11371);
   U1834 : OAI222_X1 port map( A1 => n14925, A2 => n13603, B1 => n22, B2 => 
                           n13600, C1 => n14667, C2 => n13597, ZN => n11370);
   U1835 : OAI222_X1 port map( A1 => n14919, A2 => n13603, B1 => n21, B2 => 
                           n13600, C1 => n14661, C2 => n13597, ZN => n11369);
   U1836 : OAI222_X1 port map( A1 => n14913, A2 => n13603, B1 => n20, B2 => 
                           n13600, C1 => n14655, C2 => n13597, ZN => n11368);
   U1837 : OAI222_X1 port map( A1 => n14907, A2 => n13603, B1 => n19, B2 => 
                           n13600, C1 => n14649, C2 => n13597, ZN => n11367);
   U1838 : OAI222_X1 port map( A1 => n14901, A2 => n13603, B1 => n18, B2 => 
                           n13600, C1 => n14643, C2 => n13597, ZN => n11366);
   U1839 : OAI222_X1 port map( A1 => n14895, A2 => n13603, B1 => n17, B2 => 
                           n13600, C1 => n14637, C2 => n13597, ZN => n11365);
   U1840 : OAI222_X1 port map( A1 => n14937, A2 => n13612, B1 => n16, B2 => 
                           n13609, C1 => n14679, C2 => n13606, ZN => n11404);
   U1841 : OAI222_X1 port map( A1 => n14931, A2 => n13612, B1 => n15, B2 => 
                           n13609, C1 => n14673, C2 => n13606, ZN => n11403);
   U1842 : OAI222_X1 port map( A1 => n14925, A2 => n13612, B1 => n14, B2 => 
                           n13609, C1 => n14667, C2 => n13606, ZN => n11402);
   U1843 : OAI222_X1 port map( A1 => n14919, A2 => n13612, B1 => n13, B2 => 
                           n13609, C1 => n14661, C2 => n13606, ZN => n11401);
   U1844 : OAI222_X1 port map( A1 => n14913, A2 => n13612, B1 => n12, B2 => 
                           n13609, C1 => n14655, C2 => n13606, ZN => n11400);
   U1845 : OAI222_X1 port map( A1 => n14907, A2 => n13612, B1 => n11, B2 => 
                           n13609, C1 => n14649, C2 => n13606, ZN => n11399);
   U1846 : OAI222_X1 port map( A1 => n14901, A2 => n13612, B1 => n10, B2 => 
                           n13609, C1 => n14643, C2 => n13606, ZN => n11398);
   U1847 : OAI222_X1 port map( A1 => n14895, A2 => n13612, B1 => n8, B2 => 
                           n13609, C1 => n14637, C2 => n13606, ZN => n11397);
   U1848 : OAI222_X1 port map( A1 => n14931, A2 => n13630, B1 => n7, B2 => 
                           n13627, C1 => n14673, C2 => n13624, ZN => n11467);
   U1849 : OAI222_X1 port map( A1 => n14925, A2 => n13630, B1 => n6, B2 => 
                           n13627, C1 => n14667, C2 => n13624, ZN => n11466);
   U1850 : OAI222_X1 port map( A1 => n14919, A2 => n13630, B1 => n5, B2 => 
                           n13627, C1 => n14661, C2 => n13624, ZN => n11465);
   U1851 : OAI222_X1 port map( A1 => n14913, A2 => n13630, B1 => n4, B2 => 
                           n13627, C1 => n14655, C2 => n13624, ZN => n11464);
   U1852 : OAI222_X1 port map( A1 => n14907, A2 => n13630, B1 => n3, B2 => 
                           n13627, C1 => n14649, C2 => n13624, ZN => n11463);
   U1853 : OAI222_X1 port map( A1 => n14901, A2 => n13630, B1 => n2, B2 => 
                           n13627, C1 => n14643, C2 => n13624, ZN => n11462);
   U1854 : OAI222_X1 port map( A1 => n14895, A2 => n13630, B1 => n1, B2 => 
                           n13627, C1 => n14637, C2 => n13624, ZN => n11461);
   U1855 : OAI222_X1 port map( A1 => n14936, A2 => n14373, B1 => n14370, B2 => 
                           n316, C1 => n14678, C2 => n14367, ZN => n9484);
   U1856 : OAI222_X1 port map( A1 => n14930, A2 => n14373, B1 => n14370, B2 => 
                           n315, C1 => n14672, C2 => n14367, ZN => n9483);
   U1857 : OAI222_X1 port map( A1 => n14924, A2 => n14373, B1 => n14370, B2 => 
                           n314, C1 => n14666, C2 => n14367, ZN => n9482);
   U1858 : OAI222_X1 port map( A1 => n14918, A2 => n14373, B1 => n14370, B2 => 
                           n313, C1 => n14660, C2 => n14367, ZN => n9481);
   U1859 : OAI222_X1 port map( A1 => n14912, A2 => n14373, B1 => n14370, B2 => 
                           n312, C1 => n14654, C2 => n14367, ZN => n9480);
   U1860 : OAI222_X1 port map( A1 => n14906, A2 => n14373, B1 => n14370, B2 => 
                           n311, C1 => n14648, C2 => n14367, ZN => n9479);
   U1861 : OAI222_X1 port map( A1 => n14900, A2 => n14373, B1 => n14370, B2 => 
                           n310, C1 => n14642, C2 => n14367, ZN => n9478);
   U1862 : OAI222_X1 port map( A1 => n14894, A2 => n14373, B1 => n14370, B2 => 
                           n309, C1 => n14636, C2 => n14367, ZN => n9477);
   U1863 : OAI222_X1 port map( A1 => n14940, A2 => n13243, B1 => n268, B2 => 
                           n13240, C1 => n14682, C2 => n13237, ZN => n10092);
   U1864 : OAI222_X1 port map( A1 => n14934, A2 => n13243, B1 => n267, B2 => 
                           n13240, C1 => n14676, C2 => n13237, ZN => n10091);
   U1865 : OAI222_X1 port map( A1 => n14928, A2 => n13243, B1 => n266, B2 => 
                           n13240, C1 => n14670, C2 => n13237, ZN => n10090);
   U1866 : OAI222_X1 port map( A1 => n14922, A2 => n13243, B1 => n265, B2 => 
                           n13240, C1 => n14664, C2 => n13237, ZN => n10089);
   U1867 : OAI222_X1 port map( A1 => n14916, A2 => n13243, B1 => n264, B2 => 
                           n13240, C1 => n14658, C2 => n13237, ZN => n10088);
   U1868 : OAI222_X1 port map( A1 => n14910, A2 => n13243, B1 => n263, B2 => 
                           n13240, C1 => n14652, C2 => n13237, ZN => n10087);
   U1869 : OAI222_X1 port map( A1 => n14904, A2 => n13243, B1 => n262, B2 => 
                           n13240, C1 => n14646, C2 => n13237, ZN => n10086);
   U1870 : OAI222_X1 port map( A1 => n14898, A2 => n13243, B1 => n261, B2 => 
                           n13240, C1 => n14640, C2 => n13237, ZN => n10085);
   U1871 : OAI222_X1 port map( A1 => n14940, A2 => n13252, B1 => n260, B2 => 
                           n13249, C1 => n14682, C2 => n13246, ZN => n10124);
   U1872 : OAI222_X1 port map( A1 => n14934, A2 => n13252, B1 => n259, B2 => 
                           n13249, C1 => n14676, C2 => n13246, ZN => n10123);
   U1873 : OAI222_X1 port map( A1 => n14928, A2 => n13252, B1 => n258, B2 => 
                           n13249, C1 => n14670, C2 => n13246, ZN => n10122);
   U1874 : OAI222_X1 port map( A1 => n14922, A2 => n13252, B1 => n257, B2 => 
                           n13249, C1 => n14664, C2 => n13246, ZN => n10121);
   U1875 : OAI222_X1 port map( A1 => n14916, A2 => n13252, B1 => n256, B2 => 
                           n13249, C1 => n14658, C2 => n13246, ZN => n10120);
   U1876 : OAI222_X1 port map( A1 => n14910, A2 => n13252, B1 => n255, B2 => 
                           n13249, C1 => n14652, C2 => n13246, ZN => n10119);
   U1877 : OAI222_X1 port map( A1 => n14904, A2 => n13252, B1 => n254, B2 => 
                           n13249, C1 => n14646, C2 => n13246, ZN => n10118);
   U1878 : OAI222_X1 port map( A1 => n14898, A2 => n13252, B1 => n253, B2 => 
                           n13249, C1 => n14640, C2 => n13246, ZN => n10117);
   U1879 : OAI222_X1 port map( A1 => n14940, A2 => n13270, B1 => n252, B2 => 
                           n13267, C1 => n14682, C2 => n13264, ZN => n10188);
   U1880 : OAI222_X1 port map( A1 => n14939, A2 => n13432, B1 => n163, B2 => 
                           n13429, C1 => n14680, C2 => n13426, ZN => n10764);
   U1881 : OAI222_X1 port map( A1 => n14933, A2 => n13432, B1 => n162, B2 => 
                           n13429, C1 => n14674, C2 => n13426, ZN => n10763);
   U1882 : OAI222_X1 port map( A1 => n14927, A2 => n13432, B1 => n161, B2 => 
                           n13429, C1 => n14668, C2 => n13426, ZN => n10762);
   U1883 : OAI222_X1 port map( A1 => n14921, A2 => n13432, B1 => n160, B2 => 
                           n13429, C1 => n14662, C2 => n13426, ZN => n10761);
   U1884 : OAI222_X1 port map( A1 => n14915, A2 => n13432, B1 => n159, B2 => 
                           n13429, C1 => n14656, C2 => n13426, ZN => n10760);
   U1885 : OAI222_X1 port map( A1 => n14909, A2 => n13432, B1 => n158, B2 => 
                           n13429, C1 => n14650, C2 => n13426, ZN => n10759);
   U1886 : OAI222_X1 port map( A1 => n14903, A2 => n13432, B1 => n157, B2 => 
                           n13429, C1 => n14644, C2 => n13426, ZN => n10758);
   U1887 : OAI222_X1 port map( A1 => n14897, A2 => n13432, B1 => n156, B2 => 
                           n13429, C1 => n14638, C2 => n13426, ZN => n10757);
   U1888 : OAI222_X1 port map( A1 => n14937, A2 => n13576, B1 => n48, B2 => 
                           n13573, C1 => n14679, C2 => n13570, ZN => n11276);
   U1889 : OAI222_X1 port map( A1 => n14931, A2 => n13576, B1 => n47, B2 => 
                           n13573, C1 => n14673, C2 => n13570, ZN => n11275);
   U1890 : OAI222_X1 port map( A1 => n14925, A2 => n13576, B1 => n46, B2 => 
                           n13573, C1 => n14667, C2 => n13570, ZN => n11274);
   U1891 : OAI222_X1 port map( A1 => n14919, A2 => n13576, B1 => n45, B2 => 
                           n13573, C1 => n14661, C2 => n13570, ZN => n11273);
   U1892 : OAI222_X1 port map( A1 => n14913, A2 => n13576, B1 => n44, B2 => 
                           n13573, C1 => n14655, C2 => n13570, ZN => n11272);
   U1893 : OAI222_X1 port map( A1 => n14907, A2 => n13576, B1 => n43, B2 => 
                           n13573, C1 => n14649, C2 => n13570, ZN => n11271);
   U1894 : OAI222_X1 port map( A1 => n14901, A2 => n13576, B1 => n42, B2 => 
                           n13573, C1 => n14643, C2 => n13570, ZN => n11270);
   U1895 : OAI222_X1 port map( A1 => n14895, A2 => n13576, B1 => n41, B2 => 
                           n13573, C1 => n14637, C2 => n13570, ZN => n11269);
   U1896 : OAI222_X1 port map( A1 => n14821, A2 => n13233, B1 => n2519, B2 => 
                           n13230, C1 => n14568, C2 => n13227, ZN => n10041);
   U1897 : OAI222_X1 port map( A1 => n2506, A2 => n13637, B1 => n14815, B2 => 
                           n13634, C1 => n14558, C2 => n13632, ZN => n11480);
   U1898 : OAI222_X1 port map( A1 => n2505, A2 => n13637, B1 => n14809, B2 => 
                           n13634, C1 => n14552, C2 => n13631, ZN => n11479);
   U1899 : OAI222_X1 port map( A1 => n14815, A2 => n13233, B1 => n2497, B2 => 
                           n13230, C1 => n14562, C2 => n13227, ZN => n10040);
   U1900 : OAI222_X1 port map( A1 => n14821, A2 => n14444, B1 => n14441, B2 => 
                           n2483, C1 => n14563, C2 => n14438, ZN => n9721);
   U1901 : OAI222_X1 port map( A1 => n14815, A2 => n14443, B1 => n14441, B2 => 
                           n2482, C1 => n14557, C2 => n14438, ZN => n9720);
   U1902 : OAI222_X1 port map( A1 => n14821, A2 => n14453, B1 => n14449, B2 => 
                           n2481, C1 => n14563, C2 => n14447, ZN => n9753);
   U1903 : OAI222_X1 port map( A1 => n14815, A2 => n14452, B1 => n14449, B2 => 
                           n2480, C1 => n14557, C2 => n14447, ZN => n9752);
   U1904 : OAI222_X1 port map( A1 => n14821, A2 => n14480, B1 => n14476, B2 => 
                           n2468, C1 => n14563, C2 => n14474, ZN => n9849);
   U1905 : OAI222_X1 port map( A1 => n14821, A2 => n14489, B1 => n14485, B2 => 
                           n2447, C1 => n14563, C2 => n14483, ZN => n9881);
   U1906 : OAI222_X1 port map( A1 => n14821, A2 => n14435, B1 => n14431, B2 => 
                           n2419, C1 => n14563, C2 => n14429, ZN => n9689);
   U1907 : OAI222_X1 port map( A1 => n14815, A2 => n14434, B1 => n14431, B2 => 
                           n2418, C1 => n14557, C2 => n14429, ZN => n9688);
   U1908 : OAI222_X1 port map( A1 => n14820, A2 => n13295, B1 => n2390, B2 => 
                           n13292, C1 => n14562, C2 => n13290, ZN => n10264);
   U1909 : OAI222_X1 port map( A1 => n14832, A2 => n13305, B1 => n2378, B2 => 
                           n13302, C1 => n14573, C2 => n13299, ZN => n10298);
   U1910 : OAI222_X1 port map( A1 => n14826, A2 => n13305, B1 => n2377, B2 => 
                           n13302, C1 => n14567, C2 => n13299, ZN => n10297);
   U1911 : OAI222_X1 port map( A1 => n14820, A2 => n13304, B1 => n2376, B2 => 
                           n13301, C1 => n14561, C2 => n13299, ZN => n10296);
   U1912 : OAI222_X1 port map( A1 => n14814, A2 => n13304, B1 => n2375, B2 => 
                           n13301, C1 => n14555, C2 => n13298, ZN => n10295);
   U1913 : OAI222_X1 port map( A1 => n14808, A2 => n13304, B1 => n2374, B2 => 
                           n13301, C1 => n14549, C2 => n13298, ZN => n10294);
   U1914 : OAI222_X1 port map( A1 => n14802, A2 => n13304, B1 => n2373, B2 => 
                           n13301, C1 => n14543, C2 => n13298, ZN => n10293);
   U1915 : OAI222_X1 port map( A1 => n14796, A2 => n13304, B1 => n2372, B2 => 
                           n13301, C1 => n14537, C2 => n13298, ZN => n10292);
   U1916 : OAI222_X1 port map( A1 => n14790, A2 => n13304, B1 => n2371, B2 => 
                           n13301, C1 => n14531, C2 => n13298, ZN => n10291);
   U1917 : OAI222_X1 port map( A1 => n14784, A2 => n13304, B1 => n2370, B2 => 
                           n13301, C1 => n14525, C2 => n13298, ZN => n10290);
   U1918 : OAI222_X1 port map( A1 => n14778, A2 => n13304, B1 => n2369, B2 => 
                           n13301, C1 => n14519, C2 => n13298, ZN => n10289);
   U1919 : OAI222_X1 port map( A1 => n14772, A2 => n13304, B1 => n2368, B2 => 
                           n13301, C1 => n14513, C2 => n13298, ZN => n10288);
   U1920 : OAI222_X1 port map( A1 => n14766, A2 => n13304, B1 => n2367, B2 => 
                           n13301, C1 => n14715, C2 => n13298, ZN => n10287);
   U1921 : OAI222_X1 port map( A1 => n14760, A2 => n13304, B1 => n2366, B2 => 
                           n13301, C1 => n14703, C2 => n13298, ZN => n10286);
   U1922 : OAI222_X1 port map( A1 => n14754, A2 => n13304, B1 => n2365, B2 => 
                           n13301, C1 => n14692, C2 => n13298, ZN => n10285);
   U1923 : OAI222_X1 port map( A1 => n14832, A2 => n13314, B1 => n2364, B2 => 
                           n13311, C1 => n14574, C2 => n13308, ZN => n10330);
   U1924 : OAI222_X1 port map( A1 => n14826, A2 => n13314, B1 => n2363, B2 => 
                           n13311, C1 => n14568, C2 => n13308, ZN => n10329);
   U1925 : OAI222_X1 port map( A1 => n14820, A2 => n13313, B1 => n2362, B2 => 
                           n13310, C1 => n14562, C2 => n13308, ZN => n10328);
   U1926 : OAI222_X1 port map( A1 => n14814, A2 => n13313, B1 => n2361, B2 => 
                           n13310, C1 => n14556, C2 => n13307, ZN => n10327);
   U1927 : OAI222_X1 port map( A1 => n14808, A2 => n13313, B1 => n2360, B2 => 
                           n13310, C1 => n14550, C2 => n13307, ZN => n10326);
   U1928 : OAI222_X1 port map( A1 => n14802, A2 => n13313, B1 => n2359, B2 => 
                           n13310, C1 => n14544, C2 => n13307, ZN => n10325);
   U1929 : OAI222_X1 port map( A1 => n14796, A2 => n13313, B1 => n2358, B2 => 
                           n13310, C1 => n14538, C2 => n13307, ZN => n10324);
   U1930 : OAI222_X1 port map( A1 => n14790, A2 => n13313, B1 => n2357, B2 => 
                           n13310, C1 => n14532, C2 => n13307, ZN => n10323);
   U1931 : OAI222_X1 port map( A1 => n14784, A2 => n13313, B1 => n2356, B2 => 
                           n13310, C1 => n14526, C2 => n13307, ZN => n10322);
   U1932 : OAI222_X1 port map( A1 => n14778, A2 => n13313, B1 => n2355, B2 => 
                           n13310, C1 => n14520, C2 => n13307, ZN => n10321);
   U1933 : OAI222_X1 port map( A1 => n14772, A2 => n13313, B1 => n2354, B2 => 
                           n13310, C1 => n14514, C2 => n13307, ZN => n10320);
   U1934 : OAI222_X1 port map( A1 => n14766, A2 => n13313, B1 => n2353, B2 => 
                           n13310, C1 => n14714, C2 => n13307, ZN => n10319);
   U1935 : OAI222_X1 port map( A1 => n14760, A2 => n13313, B1 => n2352, B2 => 
                           n13310, C1 => n14702, C2 => n13307, ZN => n10318);
   U1936 : OAI222_X1 port map( A1 => n14754, A2 => n13313, B1 => n2351, B2 => 
                           n13310, C1 => n14692, C2 => n13307, ZN => n10317);
   U1937 : OAI222_X1 port map( A1 => n14819, A2 => n13376, B1 => n2291, B2 => 
                           n13373, C1 => n14561, C2 => n13371, ZN => n10552);
   U1938 : OAI222_X1 port map( A1 => n14831, A2 => n13386, B1 => n2279, B2 => 
                           n13383, C1 => n14573, C2 => n13380, ZN => n10586);
   U1939 : OAI222_X1 port map( A1 => n14825, A2 => n13386, B1 => n2278, B2 => 
                           n13383, C1 => n14567, C2 => n13380, ZN => n10585);
   U1940 : OAI222_X1 port map( A1 => n14819, A2 => n13385, B1 => n2149, B2 => 
                           n13382, C1 => n14561, C2 => n13380, ZN => n10584);
   U1941 : OAI222_X1 port map( A1 => n14813, A2 => n13385, B1 => n2148, B2 => 
                           n13382, C1 => n14555, C2 => n13379, ZN => n10583);
   U1942 : OAI222_X1 port map( A1 => n14807, A2 => n13385, B1 => n2147, B2 => 
                           n13382, C1 => n14549, C2 => n13379, ZN => n10582);
   U1943 : OAI222_X1 port map( A1 => n14801, A2 => n13385, B1 => n2146, B2 => 
                           n13382, C1 => n14543, C2 => n13379, ZN => n10581);
   U1944 : OAI222_X1 port map( A1 => n14795, A2 => n13385, B1 => n2145, B2 => 
                           n13382, C1 => n14537, C2 => n13379, ZN => n10580);
   U1945 : OAI222_X1 port map( A1 => n14789, A2 => n13385, B1 => n2144, B2 => 
                           n13382, C1 => n14531, C2 => n13379, ZN => n10579);
   U1946 : OAI222_X1 port map( A1 => n14783, A2 => n13385, B1 => n2143, B2 => 
                           n13382, C1 => n14525, C2 => n13379, ZN => n10578);
   U1947 : OAI222_X1 port map( A1 => n14777, A2 => n13385, B1 => n2142, B2 => 
                           n13382, C1 => n14519, C2 => n13379, ZN => n10577);
   U1948 : OAI222_X1 port map( A1 => n14771, A2 => n13385, B1 => n2141, B2 => 
                           n13382, C1 => n14513, C2 => n13379, ZN => n10576);
   U1949 : OAI222_X1 port map( A1 => n14765, A2 => n13385, B1 => n2140, B2 => 
                           n13382, C1 => n14714, C2 => n13379, ZN => n10575);
   U1950 : OAI222_X1 port map( A1 => n14759, A2 => n13385, B1 => n2139, B2 => 
                           n13382, C1 => n14702, C2 => n13379, ZN => n10574);
   U1951 : OAI222_X1 port map( A1 => n14753, A2 => n13385, B1 => n2138, B2 => 
                           n13382, C1 => n14693, C2 => n13379, ZN => n10573);
   U1952 : OAI222_X1 port map( A1 => n14885, A2 => n13395, B1 => n2136, B2 => 
                           n13392, C1 => n14627, C2 => n13389, ZN => n10627);
   U1953 : OAI222_X1 port map( A1 => n14879, A2 => n13395, B1 => n2135, B2 => 
                           n13392, C1 => n14621, C2 => n13389, ZN => n10626);
   U1954 : OAI222_X1 port map( A1 => n14873, A2 => n13395, B1 => n2134, B2 => 
                           n13392, C1 => n14615, C2 => n13389, ZN => n10625);
   U1955 : OAI222_X1 port map( A1 => n14867, A2 => n13395, B1 => n2133, B2 => 
                           n13392, C1 => n14609, C2 => n13389, ZN => n10624);
   U1956 : OAI222_X1 port map( A1 => n14831, A2 => n13395, B1 => n2132, B2 => 
                           n13392, C1 => n14573, C2 => n13389, ZN => n10618);
   U1957 : OAI222_X1 port map( A1 => n14825, A2 => n13395, B1 => n2131, B2 => 
                           n13392, C1 => n14567, C2 => n13389, ZN => n10617);
   U1958 : OAI222_X1 port map( A1 => n14819, A2 => n13394, B1 => n2130, B2 => 
                           n13391, C1 => n14561, C2 => n13389, ZN => n10616);
   U1959 : OAI222_X1 port map( A1 => n14813, A2 => n13394, B1 => n2129, B2 => 
                           n13391, C1 => n14555, C2 => n13388, ZN => n10615);
   U1960 : OAI222_X1 port map( A1 => n14807, A2 => n13394, B1 => n2128, B2 => 
                           n13391, C1 => n14549, C2 => n13388, ZN => n10614);
   U1961 : OAI222_X1 port map( A1 => n14801, A2 => n13394, B1 => n2127, B2 => 
                           n13391, C1 => n14543, C2 => n13388, ZN => n10613);
   U1962 : OAI222_X1 port map( A1 => n14795, A2 => n13394, B1 => n2126, B2 => 
                           n13391, C1 => n14537, C2 => n13388, ZN => n10612);
   U1963 : OAI222_X1 port map( A1 => n14789, A2 => n13394, B1 => n2125, B2 => 
                           n13391, C1 => n14531, C2 => n13388, ZN => n10611);
   U1964 : OAI222_X1 port map( A1 => n14783, A2 => n13394, B1 => n2124, B2 => 
                           n13391, C1 => n14525, C2 => n13388, ZN => n10610);
   U1965 : OAI222_X1 port map( A1 => n14777, A2 => n13394, B1 => n2123, B2 => 
                           n13391, C1 => n14519, C2 => n13388, ZN => n10609);
   U1966 : OAI222_X1 port map( A1 => n14771, A2 => n13394, B1 => n2122, B2 => 
                           n13391, C1 => n14513, C2 => n13388, ZN => n10608);
   U1967 : OAI222_X1 port map( A1 => n14765, A2 => n13394, B1 => n2121, B2 => 
                           n13391, C1 => n14714, C2 => n13388, ZN => n10607);
   U1968 : OAI222_X1 port map( A1 => n14759, A2 => n13394, B1 => n2120, B2 => 
                           n13391, C1 => n14702, C2 => n13388, ZN => n10606);
   U1969 : OAI222_X1 port map( A1 => n14753, A2 => n13394, B1 => n2119, B2 => 
                           n13391, C1 => n14693, C2 => n13388, ZN => n10605);
   U1970 : OAI222_X1 port map( A1 => n14818, A2 => n13457, B1 => n2106, B2 => 
                           n13454, C1 => n14560, C2 => n13452, ZN => n10840);
   U1971 : OAI222_X1 port map( A1 => n14830, A2 => n13467, B1 => n2094, B2 => 
                           n13464, C1 => n14572, C2 => n13461, ZN => n10874);
   U1972 : OAI222_X1 port map( A1 => n14824, A2 => n13467, B1 => n2093, B2 => 
                           n13464, C1 => n14566, C2 => n13461, ZN => n10873);
   U1973 : OAI222_X1 port map( A1 => n14818, A2 => n13466, B1 => n2092, B2 => 
                           n13463, C1 => n14560, C2 => n13461, ZN => n10872);
   U1974 : OAI222_X1 port map( A1 => n14812, A2 => n13466, B1 => n2091, B2 => 
                           n13463, C1 => n14554, C2 => n13460, ZN => n10871);
   U1975 : OAI222_X1 port map( A1 => n14806, A2 => n13466, B1 => n2090, B2 => 
                           n13463, C1 => n14548, C2 => n13460, ZN => n10870);
   U1976 : OAI222_X1 port map( A1 => n14800, A2 => n13466, B1 => n2089, B2 => 
                           n13463, C1 => n14542, C2 => n13460, ZN => n10869);
   U1977 : OAI222_X1 port map( A1 => n14794, A2 => n13466, B1 => n2088, B2 => 
                           n13463, C1 => n14536, C2 => n13460, ZN => n10868);
   U1978 : OAI222_X1 port map( A1 => n14788, A2 => n13466, B1 => n2087, B2 => 
                           n13463, C1 => n14530, C2 => n13460, ZN => n10867);
   U1979 : OAI222_X1 port map( A1 => n14782, A2 => n13466, B1 => n2086, B2 => 
                           n13463, C1 => n14524, C2 => n13460, ZN => n10866);
   U1980 : OAI222_X1 port map( A1 => n14776, A2 => n13466, B1 => n2085, B2 => 
                           n13463, C1 => n14518, C2 => n13460, ZN => n10865);
   U1981 : OAI222_X1 port map( A1 => n14770, A2 => n13466, B1 => n2084, B2 => 
                           n13463, C1 => n14512, C2 => n13460, ZN => n10864);
   U1982 : OAI222_X1 port map( A1 => n14764, A2 => n13466, B1 => n2083, B2 => 
                           n13463, C1 => n14713, C2 => n13460, ZN => n10863);
   U1983 : OAI222_X1 port map( A1 => n14758, A2 => n13466, B1 => n2082, B2 => 
                           n13463, C1 => n14701, C2 => n13460, ZN => n10862);
   U1984 : OAI222_X1 port map( A1 => n14752, A2 => n13466, B1 => n2081, B2 => 
                           n13463, C1 => n14694, C2 => n13460, ZN => n10861);
   U1985 : OAI222_X1 port map( A1 => n14830, A2 => n13476, B1 => n2080, B2 => 
                           n13473, C1 => n14572, C2 => n13470, ZN => n10906);
   U1986 : OAI222_X1 port map( A1 => n14824, A2 => n13476, B1 => n2079, B2 => 
                           n13473, C1 => n14566, C2 => n13470, ZN => n10905);
   U1987 : OAI222_X1 port map( A1 => n14818, A2 => n13475, B1 => n2078, B2 => 
                           n13472, C1 => n14560, C2 => n13470, ZN => n10904);
   U1988 : OAI222_X1 port map( A1 => n14812, A2 => n13475, B1 => n2077, B2 => 
                           n13472, C1 => n14554, C2 => n13469, ZN => n10903);
   U1989 : OAI222_X1 port map( A1 => n14806, A2 => n13475, B1 => n2076, B2 => 
                           n13472, C1 => n14548, C2 => n13469, ZN => n10902);
   U1990 : OAI222_X1 port map( A1 => n14800, A2 => n13475, B1 => n2075, B2 => 
                           n13472, C1 => n14542, C2 => n13469, ZN => n10901);
   U1991 : OAI222_X1 port map( A1 => n14794, A2 => n13475, B1 => n2074, B2 => 
                           n13472, C1 => n14536, C2 => n13469, ZN => n10900);
   U1992 : OAI222_X1 port map( A1 => n14788, A2 => n13475, B1 => n2073, B2 => 
                           n13472, C1 => n14530, C2 => n13469, ZN => n10899);
   U1993 : OAI222_X1 port map( A1 => n14782, A2 => n13475, B1 => n2072, B2 => 
                           n13472, C1 => n14524, C2 => n13469, ZN => n10898);
   U1994 : OAI222_X1 port map( A1 => n14776, A2 => n13475, B1 => n2071, B2 => 
                           n13472, C1 => n14518, C2 => n13469, ZN => n10897);
   U1995 : OAI222_X1 port map( A1 => n14770, A2 => n13475, B1 => n2070, B2 => 
                           n13472, C1 => n14512, C2 => n13469, ZN => n10896);
   U1996 : OAI222_X1 port map( A1 => n14764, A2 => n13475, B1 => n2069, B2 => 
                           n13472, C1 => n14713, C2 => n13469, ZN => n10895);
   U1997 : OAI222_X1 port map( A1 => n14758, A2 => n13475, B1 => n2068, B2 => 
                           n13472, C1 => n14701, C2 => n13469, ZN => n10894);
   U1998 : OAI222_X1 port map( A1 => n14752, A2 => n13475, B1 => n2067, B2 => 
                           n13472, C1 => n14694, C2 => n13469, ZN => n10893);
   U1999 : OAI222_X1 port map( A1 => n14818, A2 => n13538, B1 => n2054, B2 => 
                           n13535, C1 => n14559, C2 => n13533, ZN => n11128);
   U2000 : OAI222_X1 port map( A1 => n14812, A2 => n13538, B1 => n2053, B2 => 
                           n13535, C1 => n14553, C2 => n13532, ZN => n11127);
   U2001 : OAI222_X1 port map( A1 => n14830, A2 => n13548, B1 => n2042, B2 => 
                           n13545, C1 => n14571, C2 => n13542, ZN => n11162);
   U2002 : OAI222_X1 port map( A1 => n14824, A2 => n13548, B1 => n2041, B2 => 
                           n13545, C1 => n14565, C2 => n13542, ZN => n11161);
   U2003 : OAI222_X1 port map( A1 => n14818, A2 => n13547, B1 => n2040, B2 => 
                           n13544, C1 => n14559, C2 => n13542, ZN => n11160);
   U2004 : OAI222_X1 port map( A1 => n14812, A2 => n13547, B1 => n2039, B2 => 
                           n13544, C1 => n14553, C2 => n13541, ZN => n11159);
   U2005 : OAI222_X1 port map( A1 => n14806, A2 => n13547, B1 => n2038, B2 => 
                           n13544, C1 => n14547, C2 => n13541, ZN => n11158);
   U2006 : OAI222_X1 port map( A1 => n14800, A2 => n13547, B1 => n2037, B2 => 
                           n13544, C1 => n14541, C2 => n13541, ZN => n11157);
   U2007 : OAI222_X1 port map( A1 => n14794, A2 => n13547, B1 => n2036, B2 => 
                           n13544, C1 => n14535, C2 => n13541, ZN => n11156);
   U2008 : OAI222_X1 port map( A1 => n14788, A2 => n13547, B1 => n2035, B2 => 
                           n13544, C1 => n14529, C2 => n13541, ZN => n11155);
   U2009 : OAI222_X1 port map( A1 => n14782, A2 => n13547, B1 => n2034, B2 => 
                           n13544, C1 => n14523, C2 => n13541, ZN => n11154);
   U2010 : OAI222_X1 port map( A1 => n14776, A2 => n13547, B1 => n2033, B2 => 
                           n13544, C1 => n14517, C2 => n13541, ZN => n11153);
   U2011 : OAI222_X1 port map( A1 => n14769, A2 => n13547, B1 => n2032, B2 => 
                           n13544, C1 => n14511, C2 => n13541, ZN => n11152);
   U2012 : OAI222_X1 port map( A1 => n14764, A2 => n13547, B1 => n2031, B2 => 
                           n13544, C1 => n14712, C2 => n13541, ZN => n11151);
   U2013 : OAI222_X1 port map( A1 => n14758, A2 => n13547, B1 => n2030, B2 => 
                           n13544, C1 => n14700, C2 => n13541, ZN => n11150);
   U2014 : OAI222_X1 port map( A1 => n14752, A2 => n13547, B1 => n2029, B2 => 
                           n13544, C1 => n14694, C2 => n13541, ZN => n11149);
   U2015 : OAI222_X1 port map( A1 => n14883, A2 => n13557, B1 => n2027, B2 => 
                           n13554, C1 => n14625, C2 => n13551, ZN => n11203);
   U2016 : OAI222_X1 port map( A1 => n14877, A2 => n13557, B1 => n2026, B2 => 
                           n13554, C1 => n14619, C2 => n13551, ZN => n11202);
   U2017 : OAI222_X1 port map( A1 => n14871, A2 => n13557, B1 => n2025, B2 => 
                           n13554, C1 => n14613, C2 => n13551, ZN => n11201);
   U2018 : OAI222_X1 port map( A1 => n14865, A2 => n13557, B1 => n2024, B2 => 
                           n13554, C1 => n14607, C2 => n13551, ZN => n11200);
   U2019 : OAI222_X1 port map( A1 => n14829, A2 => n13557, B1 => n2023, B2 => 
                           n13554, C1 => n14571, C2 => n13551, ZN => n11194);
   U2020 : OAI222_X1 port map( A1 => n14823, A2 => n13557, B1 => n2022, B2 => 
                           n13554, C1 => n14565, C2 => n13551, ZN => n11193);
   U2021 : OAI222_X1 port map( A1 => n14817, A2 => n13556, B1 => n2021, B2 => 
                           n13553, C1 => n14559, C2 => n13551, ZN => n11192);
   U2022 : OAI222_X1 port map( A1 => n14811, A2 => n13556, B1 => n2020, B2 => 
                           n13553, C1 => n14553, C2 => n13550, ZN => n11191);
   U2023 : OAI222_X1 port map( A1 => n14805, A2 => n13556, B1 => n2019, B2 => 
                           n13553, C1 => n14547, C2 => n13550, ZN => n11190);
   U2024 : OAI222_X1 port map( A1 => n14799, A2 => n13556, B1 => n2018, B2 => 
                           n13553, C1 => n14541, C2 => n13550, ZN => n11189);
   U2025 : OAI222_X1 port map( A1 => n14793, A2 => n13556, B1 => n2017, B2 => 
                           n13553, C1 => n14535, C2 => n13550, ZN => n11188);
   U2026 : OAI222_X1 port map( A1 => n14787, A2 => n13556, B1 => n2016, B2 => 
                           n13553, C1 => n14529, C2 => n13550, ZN => n11187);
   U2027 : OAI222_X1 port map( A1 => n14781, A2 => n13556, B1 => n2015, B2 => 
                           n13553, C1 => n14523, C2 => n13550, ZN => n11186);
   U2028 : OAI222_X1 port map( A1 => n14775, A2 => n13556, B1 => n2014, B2 => 
                           n13553, C1 => n14517, C2 => n13550, ZN => n11185);
   U2029 : OAI222_X1 port map( A1 => n14769, A2 => n13556, B1 => n2013, B2 => 
                           n13553, C1 => n14511, C2 => n13550, ZN => n11184);
   U2030 : OAI222_X1 port map( A1 => n14764, A2 => n13556, B1 => n2012, B2 => 
                           n13553, C1 => n14712, C2 => n13550, ZN => n11183);
   U2031 : OAI222_X1 port map( A1 => n14758, A2 => n13556, B1 => n2011, B2 => 
                           n13553, C1 => n14700, C2 => n13550, ZN => n11182);
   U2032 : OAI222_X1 port map( A1 => n14751, A2 => n13556, B1 => n2010, B2 => 
                           n13553, C1 => n14695, C2 => n13550, ZN => n11181);
   U2033 : OAI222_X1 port map( A1 => n14824, A2 => n14690, B1 => n14686, B2 => 
                           n1998, C1 => n14684, C2 => n14568, ZN => n9977);
   U2034 : OAI222_X1 port map( A1 => n14818, A2 => n14689, B1 => n14686, B2 => 
                           n1997, C1 => n14684, C2 => n14562, ZN => n9976);
   U2035 : OAI222_X1 port map( A1 => n14817, A2 => n13619, B1 => n1929, B2 => 
                           n13616, C1 => n14559, C2 => n13614, ZN => n11416);
   U2036 : OAI222_X1 port map( A1 => n14811, A2 => n13619, B1 => n1928, B2 => 
                           n13616, C1 => n14553, C2 => n13613, ZN => n11415);
   U2037 : OAI222_X1 port map( A1 => n14817, A2 => n13628, B1 => n1915, B2 => 
                           n13625, C1 => n14559, C2 => n13623, ZN => n11448);
   U2038 : OAI222_X1 port map( A1 => n14811, A2 => n13628, B1 => n1914, B2 => 
                           n13625, C1 => n14553, C2 => n13622, ZN => n11447);
   U2039 : OAI222_X1 port map( A1 => n14823, A2 => n14316, B1 => n14312, B2 => 
                           n1892, C1 => n14564, C2 => n14310, ZN => n9273);
   U2040 : OAI222_X1 port map( A1 => n14822, A2 => n14399, B1 => n14395, B2 => 
                           n1868, C1 => n14564, C2 => n14393, ZN => n9561);
   U2041 : OAI222_X1 port map( A1 => n14857, A2 => n13233, B1 => n1715, B2 => 
                           n13230, C1 => n14604, C2 => n13227, ZN => n10047);
   U2042 : OAI222_X1 port map( A1 => n14851, A2 => n13233, B1 => n1714, B2 => 
                           n13230, C1 => n14598, C2 => n13227, ZN => n10046);
   U2043 : OAI222_X1 port map( A1 => n14845, A2 => n13233, B1 => n1713, B2 => 
                           n13230, C1 => n14592, C2 => n13227, ZN => n10045);
   U2044 : OAI222_X1 port map( A1 => n14839, A2 => n13233, B1 => n1712, B2 => 
                           n13230, C1 => n14586, C2 => n13227, ZN => n10044);
   U2045 : OAI222_X1 port map( A1 => n14767, A2 => n14461, B1 => n14458, B2 => 
                           n1711, C1 => n14509, C2 => n14455, ZN => n9776);
   U2046 : OAI222_X1 port map( A1 => n14767, A2 => n14470, B1 => n14469, B2 => 
                           n1710, C1 => n14509, C2 => n14464, ZN => n9808);
   U2047 : OAI222_X1 port map( A1 => n14772, A2 => n13241, B1 => n1707, B2 => 
                           n13238, C1 => n14514, C2 => n13235, ZN => n10064);
   U2048 : OAI222_X1 port map( A1 => n14881, A2 => n14444, B1 => n14440, B2 => 
                           n1705, C1 => n14623, C2 => n14438, ZN => n9731);
   U2049 : OAI222_X1 port map( A1 => n14875, A2 => n14444, B1 => n14440, B2 => 
                           n1704, C1 => n14617, C2 => n14438, ZN => n9730);
   U2050 : OAI222_X1 port map( A1 => n14869, A2 => n14444, B1 => n14440, B2 => 
                           n1703, C1 => n14611, C2 => n14438, ZN => n9729);
   U2051 : OAI222_X1 port map( A1 => n14863, A2 => n14444, B1 => n14440, B2 => 
                           n1702, C1 => n14605, C2 => n14438, ZN => n9728);
   U2052 : OAI222_X1 port map( A1 => n14857, A2 => n14444, B1 => n14441, B2 => 
                           n1701, C1 => n14599, C2 => n14438, ZN => n9727);
   U2053 : OAI222_X1 port map( A1 => n14851, A2 => n14444, B1 => n14441, B2 => 
                           n1700, C1 => n14593, C2 => n14438, ZN => n9726);
   U2054 : OAI222_X1 port map( A1 => n14845, A2 => n14444, B1 => n14441, B2 => 
                           n1699, C1 => n14587, C2 => n14438, ZN => n9725);
   U2055 : OAI222_X1 port map( A1 => n14839, A2 => n14444, B1 => n14441, B2 => 
                           n1698, C1 => n14581, C2 => n14438, ZN => n9724);
   U2056 : OAI222_X1 port map( A1 => n14833, A2 => n14444, B1 => n14441, B2 => 
                           n1697, C1 => n14575, C2 => n14438, ZN => n9723);
   U2057 : OAI222_X1 port map( A1 => n14863, A2 => n14453, B1 => n14449, B2 => 
                           n1696, C1 => n14605, C2 => n14447, ZN => n9760);
   U2058 : OAI222_X1 port map( A1 => n14857, A2 => n14453, B1 => n14449, B2 => 
                           n1695, C1 => n14599, C2 => n14447, ZN => n9759);
   U2059 : OAI222_X1 port map( A1 => n14851, A2 => n14453, B1 => n14449, B2 => 
                           n1694, C1 => n14593, C2 => n14447, ZN => n9758);
   U2060 : OAI222_X1 port map( A1 => n14845, A2 => n14453, B1 => n14449, B2 => 
                           n1693, C1 => n14587, C2 => n14447, ZN => n9757);
   U2061 : OAI222_X1 port map( A1 => n14839, A2 => n14453, B1 => n14449, B2 => 
                           n1692, C1 => n14581, C2 => n14447, ZN => n9756);
   U2062 : OAI222_X1 port map( A1 => n14881, A2 => n14462, B1 => n14459, B2 => 
                           n1690, C1 => n14623, C2 => n14456, ZN => n9795);
   U2063 : OAI222_X1 port map( A1 => n14875, A2 => n14462, B1 => n14459, B2 => 
                           n1689, C1 => n14617, C2 => n14456, ZN => n9794);
   U2064 : OAI222_X1 port map( A1 => n14869, A2 => n14462, B1 => n14459, B2 => 
                           n1688, C1 => n14611, C2 => n14456, ZN => n9793);
   U2065 : OAI222_X1 port map( A1 => n14863, A2 => n14462, B1 => n14459, B2 => 
                           n1687, C1 => n14605, C2 => n14456, ZN => n9792);
   U2066 : OAI222_X1 port map( A1 => n14857, A2 => n14462, B1 => n14459, B2 => 
                           n1686, C1 => n14599, C2 => n14456, ZN => n9791);
   U2067 : OAI222_X1 port map( A1 => n14851, A2 => n14462, B1 => n14459, B2 => 
                           n1685, C1 => n14593, C2 => n14456, ZN => n9790);
   U2068 : OAI222_X1 port map( A1 => n14845, A2 => n14462, B1 => n14459, B2 => 
                           n1684, C1 => n14587, C2 => n14456, ZN => n9789);
   U2069 : OAI222_X1 port map( A1 => n14839, A2 => n14462, B1 => n14459, B2 => 
                           n1683, C1 => n14581, C2 => n14456, ZN => n9788);
   U2070 : OAI222_X1 port map( A1 => n14833, A2 => n14462, B1 => n14459, B2 => 
                           n1682, C1 => n14575, C2 => n14456, ZN => n9787);
   U2071 : OAI222_X1 port map( A1 => n14827, A2 => n14462, B1 => n14459, B2 => 
                           n1681, C1 => n14569, C2 => n14456, ZN => n9786);
   U2072 : OAI222_X1 port map( A1 => n14821, A2 => n14462, B1 => n14459, B2 => 
                           n1680, C1 => n14563, C2 => n14456, ZN => n9785);
   U2073 : OAI222_X1 port map( A1 => n14815, A2 => n14461, B1 => n14458, B2 => 
                           n1679, C1 => n14557, C2 => n14456, ZN => n9784);
   U2074 : OAI222_X1 port map( A1 => n14809, A2 => n14461, B1 => n14458, B2 => 
                           n1678, C1 => n14551, C2 => n14455, ZN => n9783);
   U2075 : OAI222_X1 port map( A1 => n14803, A2 => n14461, B1 => n14458, B2 => 
                           n1677, C1 => n14545, C2 => n14455, ZN => n9782);
   U2076 : OAI222_X1 port map( A1 => n14797, A2 => n14461, B1 => n14458, B2 => 
                           n1676, C1 => n14539, C2 => n14455, ZN => n9781);
   U2077 : OAI222_X1 port map( A1 => n14791, A2 => n14461, B1 => n14458, B2 => 
                           n1675, C1 => n14533, C2 => n14455, ZN => n9780);
   U2078 : OAI222_X1 port map( A1 => n14785, A2 => n14461, B1 => n14458, B2 => 
                           n1674, C1 => n14527, C2 => n14455, ZN => n9779);
   U2079 : OAI222_X1 port map( A1 => n14779, A2 => n14461, B1 => n14458, B2 => 
                           n1673, C1 => n14521, C2 => n14455, ZN => n9778);
   U2080 : OAI222_X1 port map( A1 => n14773, A2 => n14461, B1 => n14458, B2 => 
                           n1672, C1 => n14515, C2 => n14455, ZN => n9777);
   U2081 : OAI222_X1 port map( A1 => n14749, A2 => n14461, B1 => n14458, B2 => 
                           n1671, C1 => n14697, C2 => n14455, ZN => n9773);
   U2082 : OAI222_X1 port map( A1 => n14881, A2 => n14471, B1 => n14467, B2 => 
                           n1669, C1 => n14623, C2 => n14465, ZN => n9827);
   U2083 : OAI222_X1 port map( A1 => n14875, A2 => n14471, B1 => n14467, B2 => 
                           n1668, C1 => n14617, C2 => n14465, ZN => n9826);
   U2084 : OAI222_X1 port map( A1 => n14869, A2 => n14471, B1 => n14467, B2 => 
                           n1667, C1 => n14611, C2 => n14465, ZN => n9825);
   U2085 : OAI222_X1 port map( A1 => n14863, A2 => n14471, B1 => n14468, B2 => 
                           n1666, C1 => n14605, C2 => n14465, ZN => n9824);
   U2086 : OAI222_X1 port map( A1 => n14857, A2 => n14471, B1 => n14468, B2 => 
                           n1665, C1 => n14599, C2 => n14465, ZN => n9823);
   U2087 : OAI222_X1 port map( A1 => n14851, A2 => n14471, B1 => n14468, B2 => 
                           n1664, C1 => n14593, C2 => n14465, ZN => n9822);
   U2088 : OAI222_X1 port map( A1 => n14845, A2 => n14471, B1 => n14468, B2 => 
                           n1663, C1 => n14587, C2 => n14465, ZN => n9821);
   U2089 : OAI222_X1 port map( A1 => n14839, A2 => n14471, B1 => n14468, B2 => 
                           n1662, C1 => n14581, C2 => n14465, ZN => n9820);
   U2090 : OAI222_X1 port map( A1 => n14833, A2 => n14471, B1 => n14468, B2 => 
                           n1661, C1 => n14575, C2 => n14465, ZN => n9819);
   U2091 : OAI222_X1 port map( A1 => n14827, A2 => n14471, B1 => n14468, B2 => 
                           n1660, C1 => n14569, C2 => n14465, ZN => n9818);
   U2092 : OAI222_X1 port map( A1 => n14809, A2 => n14470, B1 => n14468, B2 => 
                           n1657, C1 => n14551, C2 => n14464, ZN => n9815);
   U2093 : OAI222_X1 port map( A1 => n14803, A2 => n14470, B1 => n14468, B2 => 
                           n1656, C1 => n14545, C2 => n14464, ZN => n9814);
   U2094 : OAI222_X1 port map( A1 => n14797, A2 => n14470, B1 => n14468, B2 => 
                           n1655, C1 => n14539, C2 => n14464, ZN => n9813);
   U2095 : OAI222_X1 port map( A1 => n14791, A2 => n14470, B1 => n14468, B2 => 
                           n1654, C1 => n14533, C2 => n14464, ZN => n9812);
   U2096 : OAI222_X1 port map( A1 => n14785, A2 => n14470, B1 => n14469, B2 => 
                           n1653, C1 => n14527, C2 => n14464, ZN => n9811);
   U2097 : OAI222_X1 port map( A1 => n14779, A2 => n14470, B1 => n14469, B2 => 
                           n1652, C1 => n14521, C2 => n14464, ZN => n9810);
   U2098 : OAI222_X1 port map( A1 => n14773, A2 => n14470, B1 => n14469, B2 => 
                           n1651, C1 => n14515, C2 => n14464, ZN => n9809);
   U2099 : OAI222_X1 port map( A1 => n14749, A2 => n14470, B1 => n14467, B2 => 
                           n1650, C1 => n14697, C2 => n14464, ZN => n9805);
   U2100 : OAI222_X1 port map( A1 => n14857, A2 => n14498, B1 => n14495, B2 => 
                           n1644, C1 => n14599, C2 => n14492, ZN => n9919);
   U2101 : OAI222_X1 port map( A1 => n14851, A2 => n14498, B1 => n14495, B2 => 
                           n1643, C1 => n14593, C2 => n14492, ZN => n9918);
   U2102 : OAI222_X1 port map( A1 => n14845, A2 => n14498, B1 => n14495, B2 => 
                           n1642, C1 => n14587, C2 => n14492, ZN => n9917);
   U2103 : OAI222_X1 port map( A1 => n14839, A2 => n14498, B1 => n14495, B2 => 
                           n1641, C1 => n14581, C2 => n14492, ZN => n9916);
   U2104 : OAI222_X1 port map( A1 => n14815, A2 => n14497, B1 => n14495, B2 => 
                           n1637, C1 => n14557, C2 => n14492, ZN => n9912);
   U2105 : OAI222_X1 port map( A1 => n14857, A2 => n14507, B1 => n14504, B2 => 
                           n1623, C1 => n14599, C2 => n14501, ZN => n9951);
   U2106 : OAI222_X1 port map( A1 => n14851, A2 => n14507, B1 => n14504, B2 => 
                           n1622, C1 => n14593, C2 => n14501, ZN => n9950);
   U2107 : OAI222_X1 port map( A1 => n14845, A2 => n14507, B1 => n14504, B2 => 
                           n1621, C1 => n14587, C2 => n14501, ZN => n9949);
   U2108 : OAI222_X1 port map( A1 => n14839, A2 => n14507, B1 => n14504, B2 => 
                           n1620, C1 => n14581, C2 => n14501, ZN => n9948);
   U2109 : OAI222_X1 port map( A1 => n14815, A2 => n14506, B1 => n14504, B2 => 
                           n1616, C1 => n14557, C2 => n14501, ZN => n9944);
   U2110 : OAI222_X1 port map( A1 => n14754, A2 => n13241, B1 => n1607, B2 => 
                           n13238, C1 => n14692, C2 => n13235, ZN => n10061);
   U2111 : OAI222_X1 port map( A1 => n14761, A2 => n14461, B1 => n14458, B2 => 
                           n1606, C1 => n14710, C2 => n14455, ZN => n9775);
   U2112 : OAI222_X1 port map( A1 => n14755, A2 => n14461, B1 => n14458, B2 => 
                           n1605, C1 => n14698, C2 => n14455, ZN => n9774);
   U2113 : OAI222_X1 port map( A1 => n14761, A2 => n14470, B1 => n14469, B2 => 
                           n1604, C1 => n14710, C2 => n14464, ZN => n9807);
   U2114 : OAI222_X1 port map( A1 => n14755, A2 => n14470, B1 => n14469, B2 => 
                           n1603, C1 => n14698, C2 => n14464, ZN => n9806);
   U2115 : OAI222_X1 port map( A1 => n14886, A2 => n13305, B1 => n1573, B2 => 
                           n13302, C1 => n14627, C2 => n13299, ZN => n10307);
   U2116 : OAI222_X1 port map( A1 => n14880, A2 => n13305, B1 => n1572, B2 => 
                           n13302, C1 => n14621, C2 => n13299, ZN => n10306);
   U2117 : OAI222_X1 port map( A1 => n14874, A2 => n13305, B1 => n1571, B2 => 
                           n13302, C1 => n14615, C2 => n13299, ZN => n10305);
   U2118 : OAI222_X1 port map( A1 => n14868, A2 => n13305, B1 => n1570, B2 => 
                           n13302, C1 => n14609, C2 => n13299, ZN => n10304);
   U2119 : OAI222_X1 port map( A1 => n14862, A2 => n13305, B1 => n1569, B2 => 
                           n13302, C1 => n14603, C2 => n13299, ZN => n10303);
   U2120 : OAI222_X1 port map( A1 => n14856, A2 => n13305, B1 => n1568, B2 => 
                           n13302, C1 => n14597, C2 => n13299, ZN => n10302);
   U2121 : OAI222_X1 port map( A1 => n14850, A2 => n13305, B1 => n1567, B2 => 
                           n13302, C1 => n14591, C2 => n13299, ZN => n10301);
   U2122 : OAI222_X1 port map( A1 => n14844, A2 => n13305, B1 => n1566, B2 => 
                           n13302, C1 => n14585, C2 => n13299, ZN => n10300);
   U2123 : OAI222_X1 port map( A1 => n14838, A2 => n13305, B1 => n1565, B2 => 
                           n13302, C1 => n14579, C2 => n13299, ZN => n10299);
   U2124 : OAI222_X1 port map( A1 => n14868, A2 => n13314, B1 => n1564, B2 => 
                           n13311, C1 => n14610, C2 => n13308, ZN => n10336);
   U2125 : OAI222_X1 port map( A1 => n14862, A2 => n13314, B1 => n1563, B2 => 
                           n13311, C1 => n14604, C2 => n13308, ZN => n10335);
   U2126 : OAI222_X1 port map( A1 => n14856, A2 => n13314, B1 => n1562, B2 => 
                           n13311, C1 => n14598, C2 => n13308, ZN => n10334);
   U2127 : OAI222_X1 port map( A1 => n14850, A2 => n13314, B1 => n1561, B2 => 
                           n13311, C1 => n14592, C2 => n13308, ZN => n10333);
   U2128 : OAI222_X1 port map( A1 => n14844, A2 => n13314, B1 => n1560, B2 => 
                           n13311, C1 => n14586, C2 => n13308, ZN => n10332);
   U2129 : OAI222_X1 port map( A1 => n14886, A2 => n13323, B1 => n1558, B2 => 
                           n13320, C1 => n14628, C2 => n13317, ZN => n10371);
   U2130 : OAI222_X1 port map( A1 => n14880, A2 => n13323, B1 => n1557, B2 => 
                           n13320, C1 => n14622, C2 => n13317, ZN => n10370);
   U2131 : OAI222_X1 port map( A1 => n14874, A2 => n13323, B1 => n1556, B2 => 
                           n13320, C1 => n14616, C2 => n13317, ZN => n10369);
   U2132 : OAI222_X1 port map( A1 => n14868, A2 => n13323, B1 => n1555, B2 => 
                           n13320, C1 => n14610, C2 => n13317, ZN => n10368);
   U2133 : OAI222_X1 port map( A1 => n14862, A2 => n13323, B1 => n1554, B2 => 
                           n13320, C1 => n14604, C2 => n13317, ZN => n10367);
   U2134 : OAI222_X1 port map( A1 => n14856, A2 => n13323, B1 => n1553, B2 => 
                           n13320, C1 => n14598, C2 => n13317, ZN => n10366);
   U2135 : OAI222_X1 port map( A1 => n14850, A2 => n13323, B1 => n1552, B2 => 
                           n13320, C1 => n14592, C2 => n13317, ZN => n10365);
   U2136 : OAI222_X1 port map( A1 => n14844, A2 => n13323, B1 => n1551, B2 => 
                           n13320, C1 => n14586, C2 => n13317, ZN => n10364);
   U2137 : OAI222_X1 port map( A1 => n14838, A2 => n13323, B1 => n1550, B2 => 
                           n13320, C1 => n14580, C2 => n13317, ZN => n10363);
   U2138 : OAI222_X1 port map( A1 => n14832, A2 => n13323, B1 => n1549, B2 => 
                           n13320, C1 => n14574, C2 => n13317, ZN => n10362);
   U2139 : OAI222_X1 port map( A1 => n14826, A2 => n13323, B1 => n1548, B2 => 
                           n13320, C1 => n14568, C2 => n13317, ZN => n10361);
   U2140 : OAI222_X1 port map( A1 => n14820, A2 => n13322, B1 => n1547, B2 => 
                           n13319, C1 => n14562, C2 => n13317, ZN => n10360);
   U2141 : OAI222_X1 port map( A1 => n14814, A2 => n13322, B1 => n1546, B2 => 
                           n13319, C1 => n14556, C2 => n13316, ZN => n10359);
   U2142 : OAI222_X1 port map( A1 => n14808, A2 => n13322, B1 => n1545, B2 => 
                           n13319, C1 => n14550, C2 => n13316, ZN => n10358);
   U2143 : OAI222_X1 port map( A1 => n14802, A2 => n13322, B1 => n1544, B2 => 
                           n13319, C1 => n14544, C2 => n13316, ZN => n10357);
   U2144 : OAI222_X1 port map( A1 => n14796, A2 => n13322, B1 => n1543, B2 => 
                           n13319, C1 => n14538, C2 => n13316, ZN => n10356);
   U2145 : OAI222_X1 port map( A1 => n14790, A2 => n13322, B1 => n1542, B2 => 
                           n13319, C1 => n14532, C2 => n13316, ZN => n10355);
   U2146 : OAI222_X1 port map( A1 => n14784, A2 => n13322, B1 => n1541, B2 => 
                           n13319, C1 => n14526, C2 => n13316, ZN => n10354);
   U2147 : OAI222_X1 port map( A1 => n14778, A2 => n13322, B1 => n1540, B2 => 
                           n13319, C1 => n14520, C2 => n13316, ZN => n10353);
   U2148 : OAI222_X1 port map( A1 => n14772, A2 => n13322, B1 => n1539, B2 => 
                           n13319, C1 => n14514, C2 => n13316, ZN => n10352);
   U2149 : OAI222_X1 port map( A1 => n14766, A2 => n13322, B1 => n1538, B2 => 
                           n13319, C1 => n14715, C2 => n13316, ZN => n10351);
   U2150 : OAI222_X1 port map( A1 => n14760, A2 => n13322, B1 => n1537, B2 => 
                           n13319, C1 => n14703, C2 => n13316, ZN => n10350);
   U2151 : OAI222_X1 port map( A1 => n14754, A2 => n13322, B1 => n1536, B2 => 
                           n13319, C1 => n14692, C2 => n13316, ZN => n10349);
   U2152 : OAI222_X1 port map( A1 => n14886, A2 => n13332, B1 => n1534, B2 => 
                           n13329, C1 => n14627, C2 => n13326, ZN => n10403);
   U2153 : OAI222_X1 port map( A1 => n14880, A2 => n13332, B1 => n1533, B2 => 
                           n13329, C1 => n14621, C2 => n13326, ZN => n10402);
   U2154 : OAI222_X1 port map( A1 => n14874, A2 => n13332, B1 => n1532, B2 => 
                           n13329, C1 => n14615, C2 => n13326, ZN => n10401);
   U2155 : OAI222_X1 port map( A1 => n14868, A2 => n13332, B1 => n1531, B2 => 
                           n13329, C1 => n14609, C2 => n13326, ZN => n10400);
   U2156 : OAI222_X1 port map( A1 => n14862, A2 => n13332, B1 => n1530, B2 => 
                           n13329, C1 => n14603, C2 => n13326, ZN => n10399);
   U2157 : OAI222_X1 port map( A1 => n14856, A2 => n13332, B1 => n1529, B2 => 
                           n13329, C1 => n14597, C2 => n13326, ZN => n10398);
   U2158 : OAI222_X1 port map( A1 => n14850, A2 => n13332, B1 => n1528, B2 => 
                           n13329, C1 => n14591, C2 => n13326, ZN => n10397);
   U2159 : OAI222_X1 port map( A1 => n14844, A2 => n13332, B1 => n1527, B2 => 
                           n13329, C1 => n14585, C2 => n13326, ZN => n10396);
   U2160 : OAI222_X1 port map( A1 => n14838, A2 => n13332, B1 => n1526, B2 => 
                           n13329, C1 => n14579, C2 => n13326, ZN => n10395);
   U2161 : OAI222_X1 port map( A1 => n14832, A2 => n13332, B1 => n1525, B2 => 
                           n13329, C1 => n14573, C2 => n13326, ZN => n10394);
   U2162 : OAI222_X1 port map( A1 => n14826, A2 => n13332, B1 => n1524, B2 => 
                           n13329, C1 => n14567, C2 => n13326, ZN => n10393);
   U2163 : OAI222_X1 port map( A1 => n14820, A2 => n13331, B1 => n1523, B2 => 
                           n13328, C1 => n14561, C2 => n13326, ZN => n10392);
   U2164 : OAI222_X1 port map( A1 => n14814, A2 => n13331, B1 => n1522, B2 => 
                           n13328, C1 => n14555, C2 => n13325, ZN => n10391);
   U2165 : OAI222_X1 port map( A1 => n14808, A2 => n13331, B1 => n1521, B2 => 
                           n13328, C1 => n14549, C2 => n13325, ZN => n10390);
   U2166 : OAI222_X1 port map( A1 => n14802, A2 => n13331, B1 => n1520, B2 => 
                           n13328, C1 => n14543, C2 => n13325, ZN => n10389);
   U2167 : OAI222_X1 port map( A1 => n14796, A2 => n13331, B1 => n1519, B2 => 
                           n13328, C1 => n14537, C2 => n13325, ZN => n10388);
   U2168 : OAI222_X1 port map( A1 => n14790, A2 => n13331, B1 => n1518, B2 => 
                           n13328, C1 => n14531, C2 => n13325, ZN => n10387);
   U2169 : OAI222_X1 port map( A1 => n14784, A2 => n13331, B1 => n1517, B2 => 
                           n13328, C1 => n14525, C2 => n13325, ZN => n10386);
   U2170 : OAI222_X1 port map( A1 => n14778, A2 => n13331, B1 => n1516, B2 => 
                           n13328, C1 => n14519, C2 => n13325, ZN => n10385);
   U2171 : OAI222_X1 port map( A1 => n14772, A2 => n13331, B1 => n1515, B2 => 
                           n13328, C1 => n14513, C2 => n13325, ZN => n10384);
   U2172 : OAI222_X1 port map( A1 => n14766, A2 => n13331, B1 => n1514, B2 => 
                           n13328, C1 => n14715, C2 => n13325, ZN => n10383);
   U2173 : OAI222_X1 port map( A1 => n14760, A2 => n13331, B1 => n1513, B2 => 
                           n13328, C1 => n14703, C2 => n13325, ZN => n10382);
   U2174 : OAI222_X1 port map( A1 => n14754, A2 => n13331, B1 => n1512, B2 => 
                           n13328, C1 => n14692, C2 => n13325, ZN => n10381);
   U2175 : OAI222_X1 port map( A1 => n14753, A2 => n13349, B1 => n1511, B2 => 
                           n13346, C1 => n14693, C2 => n13343, ZN => n10445);
   U2176 : OAI222_X1 port map( A1 => n14885, A2 => n13386, B1 => n1461, B2 => 
                           n13383, C1 => n14627, C2 => n13380, ZN => n10595);
   U2177 : OAI222_X1 port map( A1 => n14879, A2 => n13386, B1 => n1460, B2 => 
                           n13383, C1 => n14621, C2 => n13380, ZN => n10594);
   U2178 : OAI222_X1 port map( A1 => n14873, A2 => n13386, B1 => n1459, B2 => 
                           n13383, C1 => n14615, C2 => n13380, ZN => n10593);
   U2179 : OAI222_X1 port map( A1 => n14867, A2 => n13386, B1 => n1458, B2 => 
                           n13383, C1 => n14609, C2 => n13380, ZN => n10592);
   U2180 : OAI222_X1 port map( A1 => n14861, A2 => n13386, B1 => n1457, B2 => 
                           n13383, C1 => n14603, C2 => n13380, ZN => n10591);
   U2181 : OAI222_X1 port map( A1 => n14855, A2 => n13386, B1 => n1456, B2 => 
                           n13383, C1 => n14597, C2 => n13380, ZN => n10590);
   U2182 : OAI222_X1 port map( A1 => n14849, A2 => n13386, B1 => n1455, B2 => 
                           n13383, C1 => n14591, C2 => n13380, ZN => n10589);
   U2183 : OAI222_X1 port map( A1 => n14843, A2 => n13386, B1 => n1454, B2 => 
                           n13383, C1 => n14585, C2 => n13380, ZN => n10588);
   U2184 : OAI222_X1 port map( A1 => n14837, A2 => n13386, B1 => n1453, B2 => 
                           n13383, C1 => n14579, C2 => n13380, ZN => n10587);
   U2185 : OAI222_X1 port map( A1 => n14861, A2 => n13395, B1 => n1452, B2 => 
                           n13392, C1 => n14603, C2 => n13389, ZN => n10623);
   U2186 : OAI222_X1 port map( A1 => n14855, A2 => n13395, B1 => n1451, B2 => 
                           n13392, C1 => n14597, C2 => n13389, ZN => n10622);
   U2187 : OAI222_X1 port map( A1 => n14849, A2 => n13395, B1 => n1450, B2 => 
                           n13392, C1 => n14591, C2 => n13389, ZN => n10621);
   U2188 : OAI222_X1 port map( A1 => n14843, A2 => n13395, B1 => n1449, B2 => 
                           n13392, C1 => n14585, C2 => n13389, ZN => n10620);
   U2189 : OAI222_X1 port map( A1 => n14837, A2 => n13395, B1 => n1448, B2 => 
                           n13392, C1 => n14579, C2 => n13389, ZN => n10619);
   U2190 : OAI222_X1 port map( A1 => n14885, A2 => n13413, B1 => n1422, B2 => 
                           n13410, C1 => n14627, C2 => n13407, ZN => n10691);
   U2191 : OAI222_X1 port map( A1 => n14879, A2 => n13413, B1 => n1421, B2 => 
                           n13410, C1 => n14621, C2 => n13407, ZN => n10690);
   U2192 : OAI222_X1 port map( A1 => n14873, A2 => n13413, B1 => n1420, B2 => 
                           n13410, C1 => n14615, C2 => n13407, ZN => n10689);
   U2193 : OAI222_X1 port map( A1 => n14867, A2 => n13413, B1 => n1419, B2 => 
                           n13410, C1 => n14609, C2 => n13407, ZN => n10688);
   U2194 : OAI222_X1 port map( A1 => n14861, A2 => n13413, B1 => n1418, B2 => 
                           n13410, C1 => n14603, C2 => n13407, ZN => n10687);
   U2195 : OAI222_X1 port map( A1 => n14855, A2 => n13413, B1 => n1417, B2 => 
                           n13410, C1 => n14597, C2 => n13407, ZN => n10686);
   U2196 : OAI222_X1 port map( A1 => n14849, A2 => n13413, B1 => n1416, B2 => 
                           n13410, C1 => n14591, C2 => n13407, ZN => n10685);
   U2197 : OAI222_X1 port map( A1 => n14843, A2 => n13413, B1 => n1415, B2 => 
                           n13410, C1 => n14585, C2 => n13407, ZN => n10684);
   U2198 : OAI222_X1 port map( A1 => n14837, A2 => n13413, B1 => n1414, B2 => 
                           n13410, C1 => n14579, C2 => n13407, ZN => n10683);
   U2199 : OAI222_X1 port map( A1 => n14831, A2 => n13413, B1 => n1413, B2 => 
                           n13410, C1 => n14573, C2 => n13407, ZN => n10682);
   U2200 : OAI222_X1 port map( A1 => n14825, A2 => n13413, B1 => n1412, B2 => 
                           n13410, C1 => n14567, C2 => n13407, ZN => n10681);
   U2201 : OAI222_X1 port map( A1 => n14819, A2 => n13412, B1 => n1411, B2 => 
                           n13409, C1 => n14561, C2 => n13407, ZN => n10680);
   U2202 : OAI222_X1 port map( A1 => n14813, A2 => n13412, B1 => n1410, B2 => 
                           n13409, C1 => n14555, C2 => n13406, ZN => n10679);
   U2203 : OAI222_X1 port map( A1 => n14807, A2 => n13412, B1 => n1409, B2 => 
                           n13409, C1 => n14549, C2 => n13406, ZN => n10678);
   U2204 : OAI222_X1 port map( A1 => n14801, A2 => n13412, B1 => n1408, B2 => 
                           n13409, C1 => n14543, C2 => n13406, ZN => n10677);
   U2205 : OAI222_X1 port map( A1 => n14795, A2 => n13412, B1 => n1407, B2 => 
                           n13409, C1 => n14537, C2 => n13406, ZN => n10676);
   U2206 : OAI222_X1 port map( A1 => n14789, A2 => n13412, B1 => n1406, B2 => 
                           n13409, C1 => n14531, C2 => n13406, ZN => n10675);
   U2207 : OAI222_X1 port map( A1 => n14783, A2 => n13412, B1 => n1405, B2 => 
                           n13409, C1 => n14525, C2 => n13406, ZN => n10674);
   U2208 : OAI222_X1 port map( A1 => n14777, A2 => n13412, B1 => n1404, B2 => 
                           n13409, C1 => n14519, C2 => n13406, ZN => n10673);
   U2209 : OAI222_X1 port map( A1 => n14771, A2 => n13412, B1 => n1403, B2 => 
                           n13409, C1 => n14513, C2 => n13406, ZN => n10672);
   U2210 : OAI222_X1 port map( A1 => n14765, A2 => n13412, B1 => n1402, B2 => 
                           n13409, C1 => n14714, C2 => n13406, ZN => n10671);
   U2211 : OAI222_X1 port map( A1 => n14759, A2 => n13412, B1 => n1401, B2 => 
                           n13409, C1 => n14702, C2 => n13406, ZN => n10670);
   U2212 : OAI222_X1 port map( A1 => n14753, A2 => n13412, B1 => n1400, B2 => 
                           n13409, C1 => n14693, C2 => n13406, ZN => n10669);
   U2213 : OAI222_X1 port map( A1 => n14885, A2 => n13422, B1 => n1398, B2 => 
                           n13419, C1 => n14627, C2 => n13416, ZN => n10723);
   U2214 : OAI222_X1 port map( A1 => n14879, A2 => n13422, B1 => n1397, B2 => 
                           n13419, C1 => n14621, C2 => n13416, ZN => n10722);
   U2215 : OAI222_X1 port map( A1 => n14873, A2 => n13422, B1 => n1396, B2 => 
                           n13419, C1 => n14615, C2 => n13416, ZN => n10721);
   U2216 : OAI222_X1 port map( A1 => n14867, A2 => n13422, B1 => n1395, B2 => 
                           n13419, C1 => n14609, C2 => n13416, ZN => n10720);
   U2217 : OAI222_X1 port map( A1 => n14861, A2 => n13422, B1 => n1394, B2 => 
                           n13419, C1 => n14603, C2 => n13416, ZN => n10719);
   U2218 : OAI222_X1 port map( A1 => n14855, A2 => n13422, B1 => n1393, B2 => 
                           n13419, C1 => n14597, C2 => n13416, ZN => n10718);
   U2219 : OAI222_X1 port map( A1 => n14849, A2 => n13422, B1 => n1392, B2 => 
                           n13419, C1 => n14591, C2 => n13416, ZN => n10717);
   U2220 : OAI222_X1 port map( A1 => n14843, A2 => n13422, B1 => n1391, B2 => 
                           n13419, C1 => n14585, C2 => n13416, ZN => n10716);
   U2221 : OAI222_X1 port map( A1 => n14837, A2 => n13422, B1 => n1390, B2 => 
                           n13419, C1 => n14579, C2 => n13416, ZN => n10715);
   U2222 : OAI222_X1 port map( A1 => n14831, A2 => n13422, B1 => n1389, B2 => 
                           n13419, C1 => n14573, C2 => n13416, ZN => n10714);
   U2223 : OAI222_X1 port map( A1 => n14825, A2 => n13422, B1 => n1388, B2 => 
                           n13419, C1 => n14567, C2 => n13416, ZN => n10713);
   U2224 : OAI222_X1 port map( A1 => n14819, A2 => n13421, B1 => n1387, B2 => 
                           n13418, C1 => n14561, C2 => n13416, ZN => n10712);
   U2225 : OAI222_X1 port map( A1 => n14813, A2 => n13421, B1 => n1386, B2 => 
                           n13418, C1 => n14555, C2 => n13415, ZN => n10711);
   U2226 : OAI222_X1 port map( A1 => n14807, A2 => n13421, B1 => n1385, B2 => 
                           n13418, C1 => n14549, C2 => n13415, ZN => n10710);
   U2227 : OAI222_X1 port map( A1 => n14801, A2 => n13421, B1 => n1384, B2 => 
                           n13418, C1 => n14543, C2 => n13415, ZN => n10709);
   U2228 : OAI222_X1 port map( A1 => n14795, A2 => n13421, B1 => n1383, B2 => 
                           n13418, C1 => n14537, C2 => n13415, ZN => n10708);
   U2229 : OAI222_X1 port map( A1 => n14789, A2 => n13421, B1 => n1382, B2 => 
                           n13418, C1 => n14531, C2 => n13415, ZN => n10707);
   U2230 : OAI222_X1 port map( A1 => n14783, A2 => n13421, B1 => n1381, B2 => 
                           n13418, C1 => n14525, C2 => n13415, ZN => n10706);
   U2231 : OAI222_X1 port map( A1 => n14777, A2 => n13421, B1 => n1380, B2 => 
                           n13418, C1 => n14519, C2 => n13415, ZN => n10705);
   U2232 : OAI222_X1 port map( A1 => n14771, A2 => n13421, B1 => n1379, B2 => 
                           n13418, C1 => n14513, C2 => n13415, ZN => n10704);
   U2233 : OAI222_X1 port map( A1 => n14765, A2 => n13421, B1 => n1378, B2 => 
                           n13418, C1 => n14714, C2 => n13415, ZN => n10703);
   U2234 : OAI222_X1 port map( A1 => n14759, A2 => n13421, B1 => n1377, B2 => 
                           n13418, C1 => n14702, C2 => n13415, ZN => n10702);
   U2235 : OAI222_X1 port map( A1 => n14753, A2 => n13421, B1 => n1376, B2 => 
                           n13418, C1 => n14693, C2 => n13415, ZN => n10701);
   U2236 : OAI222_X1 port map( A1 => n14891, A2 => n13431, B1 => n1375, B2 => 
                           n13428, C1 => n14632, C2 => n13425, ZN => n10756);
   U2237 : OAI222_X1 port map( A1 => n14885, A2 => n13431, B1 => n1374, B2 => 
                           n13428, C1 => n14626, C2 => n13425, ZN => n10755);
   U2238 : OAI222_X1 port map( A1 => n14879, A2 => n13431, B1 => n1373, B2 => 
                           n13428, C1 => n14620, C2 => n13425, ZN => n10754);
   U2239 : OAI222_X1 port map( A1 => n14873, A2 => n13431, B1 => n1372, B2 => 
                           n13428, C1 => n14614, C2 => n13425, ZN => n10753);
   U2240 : OAI222_X1 port map( A1 => n14867, A2 => n13431, B1 => n1371, B2 => 
                           n13428, C1 => n14608, C2 => n13425, ZN => n10752);
   U2241 : OAI222_X1 port map( A1 => n14861, A2 => n13431, B1 => n1370, B2 => 
                           n13428, C1 => n14602, C2 => n13425, ZN => n10751);
   U2242 : OAI222_X1 port map( A1 => n14855, A2 => n13431, B1 => n1369, B2 => 
                           n13428, C1 => n14596, C2 => n13425, ZN => n10750);
   U2243 : OAI222_X1 port map( A1 => n14849, A2 => n13431, B1 => n1368, B2 => 
                           n13428, C1 => n14590, C2 => n13425, ZN => n10749);
   U2244 : OAI222_X1 port map( A1 => n14843, A2 => n13431, B1 => n1367, B2 => 
                           n13428, C1 => n14584, C2 => n13425, ZN => n10748);
   U2245 : OAI222_X1 port map( A1 => n14837, A2 => n13431, B1 => n1366, B2 => 
                           n13428, C1 => n14578, C2 => n13425, ZN => n10747);
   U2246 : OAI222_X1 port map( A1 => n14831, A2 => n13431, B1 => n1365, B2 => 
                           n13428, C1 => n14572, C2 => n13425, ZN => n10746);
   U2247 : OAI222_X1 port map( A1 => n14825, A2 => n13431, B1 => n1364, B2 => 
                           n13428, C1 => n14566, C2 => n13425, ZN => n10745);
   U2248 : OAI222_X1 port map( A1 => n14819, A2 => n13430, B1 => n1363, B2 => 
                           n13427, C1 => n14560, C2 => n13425, ZN => n10744);
   U2249 : OAI222_X1 port map( A1 => n14813, A2 => n13430, B1 => n1362, B2 => 
                           n13427, C1 => n14554, C2 => n13424, ZN => n10743);
   U2250 : OAI222_X1 port map( A1 => n14807, A2 => n13430, B1 => n1361, B2 => 
                           n13427, C1 => n14548, C2 => n13424, ZN => n10742);
   U2251 : OAI222_X1 port map( A1 => n14801, A2 => n13430, B1 => n1360, B2 => 
                           n13427, C1 => n14542, C2 => n13424, ZN => n10741);
   U2252 : OAI222_X1 port map( A1 => n14795, A2 => n13430, B1 => n1359, B2 => 
                           n13427, C1 => n14536, C2 => n13424, ZN => n10740);
   U2253 : OAI222_X1 port map( A1 => n14789, A2 => n13430, B1 => n1358, B2 => 
                           n13427, C1 => n14530, C2 => n13424, ZN => n10739);
   U2254 : OAI222_X1 port map( A1 => n14783, A2 => n13430, B1 => n1357, B2 => 
                           n13427, C1 => n14524, C2 => n13424, ZN => n10738);
   U2255 : OAI222_X1 port map( A1 => n14777, A2 => n13430, B1 => n1356, B2 => 
                           n13427, C1 => n14518, C2 => n13424, ZN => n10737);
   U2256 : OAI222_X1 port map( A1 => n14771, A2 => n13430, B1 => n1355, B2 => 
                           n13427, C1 => n14512, C2 => n13424, ZN => n10736);
   U2257 : OAI222_X1 port map( A1 => n14765, A2 => n13430, B1 => n1354, B2 => 
                           n13427, C1 => n14714, C2 => n13424, ZN => n10735);
   U2258 : OAI222_X1 port map( A1 => n14759, A2 => n13430, B1 => n1353, B2 => 
                           n13427, C1 => n14702, C2 => n13424, ZN => n10734);
   U2259 : OAI222_X1 port map( A1 => n14753, A2 => n13430, B1 => n1352, B2 => 
                           n13427, C1 => n14693, C2 => n13424, ZN => n10733);
   U2260 : OAI222_X1 port map( A1 => n14884, A2 => n13467, B1 => n1302, B2 => 
                           n13464, C1 => n14626, C2 => n13461, ZN => n10883);
   U2261 : OAI222_X1 port map( A1 => n14878, A2 => n13467, B1 => n1301, B2 => 
                           n13464, C1 => n14620, C2 => n13461, ZN => n10882);
   U2262 : OAI222_X1 port map( A1 => n14872, A2 => n13467, B1 => n1300, B2 => 
                           n13464, C1 => n14614, C2 => n13461, ZN => n10881);
   U2263 : OAI222_X1 port map( A1 => n14866, A2 => n13467, B1 => n1299, B2 => 
                           n13464, C1 => n14608, C2 => n13461, ZN => n10880);
   U2264 : OAI222_X1 port map( A1 => n14860, A2 => n13467, B1 => n1298, B2 => 
                           n13464, C1 => n14602, C2 => n13461, ZN => n10879);
   U2265 : OAI222_X1 port map( A1 => n14854, A2 => n13467, B1 => n1297, B2 => 
                           n13464, C1 => n14596, C2 => n13461, ZN => n10878);
   U2266 : OAI222_X1 port map( A1 => n14848, A2 => n13467, B1 => n1296, B2 => 
                           n13464, C1 => n14590, C2 => n13461, ZN => n10877);
   U2267 : OAI222_X1 port map( A1 => n14842, A2 => n13467, B1 => n1295, B2 => 
                           n13464, C1 => n14584, C2 => n13461, ZN => n10876);
   U2268 : OAI222_X1 port map( A1 => n14836, A2 => n13467, B1 => n1294, B2 => 
                           n13464, C1 => n14578, C2 => n13461, ZN => n10875);
   U2269 : OAI222_X1 port map( A1 => n14860, A2 => n13476, B1 => n1293, B2 => 
                           n13473, C1 => n14602, C2 => n13470, ZN => n10911);
   U2270 : OAI222_X1 port map( A1 => n14854, A2 => n13476, B1 => n1292, B2 => 
                           n13473, C1 => n14596, C2 => n13470, ZN => n10910);
   U2271 : OAI222_X1 port map( A1 => n14848, A2 => n13476, B1 => n1291, B2 => 
                           n13473, C1 => n14590, C2 => n13470, ZN => n10909);
   U2272 : OAI222_X1 port map( A1 => n14842, A2 => n13476, B1 => n1290, B2 => 
                           n13473, C1 => n14584, C2 => n13470, ZN => n10908);
   U2273 : OAI222_X1 port map( A1 => n14836, A2 => n13476, B1 => n1289, B2 => 
                           n13473, C1 => n14578, C2 => n13470, ZN => n10907);
   U2274 : OAI222_X1 port map( A1 => n14884, A2 => n13485, B1 => n1287, B2 => 
                           n13482, C1 => n14626, C2 => n13479, ZN => n10947);
   U2275 : OAI222_X1 port map( A1 => n14878, A2 => n13485, B1 => n1286, B2 => 
                           n13482, C1 => n14620, C2 => n13479, ZN => n10946);
   U2276 : OAI222_X1 port map( A1 => n14872, A2 => n13485, B1 => n1285, B2 => 
                           n13482, C1 => n14614, C2 => n13479, ZN => n10945);
   U2277 : OAI222_X1 port map( A1 => n14866, A2 => n13485, B1 => n1284, B2 => 
                           n13482, C1 => n14608, C2 => n13479, ZN => n10944);
   U2278 : OAI222_X1 port map( A1 => n14860, A2 => n13485, B1 => n1283, B2 => 
                           n13482, C1 => n14602, C2 => n13479, ZN => n10943);
   U2279 : OAI222_X1 port map( A1 => n14854, A2 => n13485, B1 => n1282, B2 => 
                           n13482, C1 => n14596, C2 => n13479, ZN => n10942);
   U2280 : OAI222_X1 port map( A1 => n14848, A2 => n13485, B1 => n1281, B2 => 
                           n13482, C1 => n14590, C2 => n13479, ZN => n10941);
   U2281 : OAI222_X1 port map( A1 => n14842, A2 => n13485, B1 => n1280, B2 => 
                           n13482, C1 => n14584, C2 => n13479, ZN => n10940);
   U2282 : OAI222_X1 port map( A1 => n14836, A2 => n13485, B1 => n1279, B2 => 
                           n13482, C1 => n14578, C2 => n13479, ZN => n10939);
   U2283 : OAI222_X1 port map( A1 => n14830, A2 => n13485, B1 => n1278, B2 => 
                           n13482, C1 => n14572, C2 => n13479, ZN => n10938);
   U2284 : OAI222_X1 port map( A1 => n14824, A2 => n13485, B1 => n1277, B2 => 
                           n13482, C1 => n14566, C2 => n13479, ZN => n10937);
   U2285 : OAI222_X1 port map( A1 => n14818, A2 => n13484, B1 => n1276, B2 => 
                           n13481, C1 => n14560, C2 => n13479, ZN => n10936);
   U2286 : OAI222_X1 port map( A1 => n14812, A2 => n13484, B1 => n1275, B2 => 
                           n13481, C1 => n14554, C2 => n13478, ZN => n10935);
   U2287 : OAI222_X1 port map( A1 => n14806, A2 => n13484, B1 => n1274, B2 => 
                           n13481, C1 => n14548, C2 => n13478, ZN => n10934);
   U2288 : OAI222_X1 port map( A1 => n14800, A2 => n13484, B1 => n1273, B2 => 
                           n13481, C1 => n14542, C2 => n13478, ZN => n10933);
   U2289 : OAI222_X1 port map( A1 => n14794, A2 => n13484, B1 => n1272, B2 => 
                           n13481, C1 => n14536, C2 => n13478, ZN => n10932);
   U2290 : OAI222_X1 port map( A1 => n14788, A2 => n13484, B1 => n1271, B2 => 
                           n13481, C1 => n14530, C2 => n13478, ZN => n10931);
   U2291 : OAI222_X1 port map( A1 => n14782, A2 => n13484, B1 => n1270, B2 => 
                           n13481, C1 => n14524, C2 => n13478, ZN => n10930);
   U2292 : OAI222_X1 port map( A1 => n14776, A2 => n13484, B1 => n1269, B2 => 
                           n13481, C1 => n14518, C2 => n13478, ZN => n10929);
   U2293 : OAI222_X1 port map( A1 => n14770, A2 => n13484, B1 => n1268, B2 => 
                           n13481, C1 => n14512, C2 => n13478, ZN => n10928);
   U2294 : OAI222_X1 port map( A1 => n14764, A2 => n13484, B1 => n1267, B2 => 
                           n13481, C1 => n14713, C2 => n13478, ZN => n10927);
   U2295 : OAI222_X1 port map( A1 => n14758, A2 => n13484, B1 => n1266, B2 => 
                           n13481, C1 => n14701, C2 => n13478, ZN => n10926);
   U2296 : OAI222_X1 port map( A1 => n14752, A2 => n13484, B1 => n1265, B2 => 
                           n13481, C1 => n14694, C2 => n13478, ZN => n10925);
   U2297 : OAI222_X1 port map( A1 => n14884, A2 => n13494, B1 => n1263, B2 => 
                           n13491, C1 => n14626, C2 => n13488, ZN => n10979);
   U2298 : OAI222_X1 port map( A1 => n14878, A2 => n13494, B1 => n1262, B2 => 
                           n13491, C1 => n14620, C2 => n13488, ZN => n10978);
   U2299 : OAI222_X1 port map( A1 => n14872, A2 => n13494, B1 => n1261, B2 => 
                           n13491, C1 => n14614, C2 => n13488, ZN => n10977);
   U2300 : OAI222_X1 port map( A1 => n14866, A2 => n13494, B1 => n1260, B2 => 
                           n13491, C1 => n14608, C2 => n13488, ZN => n10976);
   U2301 : OAI222_X1 port map( A1 => n14860, A2 => n13494, B1 => n1259, B2 => 
                           n13491, C1 => n14602, C2 => n13488, ZN => n10975);
   U2302 : OAI222_X1 port map( A1 => n14854, A2 => n13494, B1 => n1258, B2 => 
                           n13491, C1 => n14596, C2 => n13488, ZN => n10974);
   U2303 : OAI222_X1 port map( A1 => n14848, A2 => n13494, B1 => n1257, B2 => 
                           n13491, C1 => n14590, C2 => n13488, ZN => n10973);
   U2304 : OAI222_X1 port map( A1 => n14842, A2 => n13494, B1 => n1256, B2 => 
                           n13491, C1 => n14584, C2 => n13488, ZN => n10972);
   U2305 : OAI222_X1 port map( A1 => n14836, A2 => n13494, B1 => n1255, B2 => 
                           n13491, C1 => n14578, C2 => n13488, ZN => n10971);
   U2306 : OAI222_X1 port map( A1 => n14830, A2 => n13494, B1 => n1254, B2 => 
                           n13491, C1 => n14572, C2 => n13488, ZN => n10970);
   U2307 : OAI222_X1 port map( A1 => n14824, A2 => n13494, B1 => n1253, B2 => 
                           n13491, C1 => n14566, C2 => n13488, ZN => n10969);
   U2308 : OAI222_X1 port map( A1 => n14812, A2 => n13493, B1 => n1251, B2 => 
                           n13490, C1 => n14554, C2 => n13487, ZN => n10967);
   U2309 : OAI222_X1 port map( A1 => n14806, A2 => n13493, B1 => n1250, B2 => 
                           n13490, C1 => n14548, C2 => n13487, ZN => n10966);
   U2310 : OAI222_X1 port map( A1 => n14800, A2 => n13493, B1 => n1249, B2 => 
                           n13490, C1 => n14542, C2 => n13487, ZN => n10965);
   U2311 : OAI222_X1 port map( A1 => n14794, A2 => n13493, B1 => n1248, B2 => 
                           n13490, C1 => n14536, C2 => n13487, ZN => n10964);
   U2312 : OAI222_X1 port map( A1 => n14788, A2 => n13493, B1 => n1247, B2 => 
                           n13490, C1 => n14530, C2 => n13487, ZN => n10963);
   U2313 : OAI222_X1 port map( A1 => n14782, A2 => n13493, B1 => n1246, B2 => 
                           n13490, C1 => n14524, C2 => n13487, ZN => n10962);
   U2314 : OAI222_X1 port map( A1 => n14776, A2 => n13493, B1 => n1245, B2 => 
                           n13490, C1 => n14518, C2 => n13487, ZN => n10961);
   U2315 : OAI222_X1 port map( A1 => n14770, A2 => n13493, B1 => n1244, B2 => 
                           n13490, C1 => n14512, C2 => n13487, ZN => n10960);
   U2316 : OAI222_X1 port map( A1 => n14764, A2 => n13493, B1 => n1243, B2 => 
                           n13490, C1 => n14713, C2 => n13487, ZN => n10959);
   U2317 : OAI222_X1 port map( A1 => n14758, A2 => n13493, B1 => n1242, B2 => 
                           n13490, C1 => n14701, C2 => n13487, ZN => n10958);
   U2318 : OAI222_X1 port map( A1 => n14752, A2 => n13493, B1 => n1241, B2 => 
                           n13490, C1 => n14694, C2 => n13487, ZN => n10957);
   U2319 : OAI222_X1 port map( A1 => n14884, A2 => n13503, B1 => n1239, B2 => 
                           n13500, C1 => n14626, C2 => n13497, ZN => n11011);
   U2320 : OAI222_X1 port map( A1 => n14878, A2 => n13503, B1 => n1238, B2 => 
                           n13500, C1 => n14620, C2 => n13497, ZN => n11010);
   U2321 : OAI222_X1 port map( A1 => n14872, A2 => n13503, B1 => n1237, B2 => 
                           n13500, C1 => n14614, C2 => n13497, ZN => n11009);
   U2322 : OAI222_X1 port map( A1 => n14866, A2 => n13503, B1 => n1236, B2 => 
                           n13500, C1 => n14608, C2 => n13497, ZN => n11008);
   U2323 : OAI222_X1 port map( A1 => n14860, A2 => n13503, B1 => n1235, B2 => 
                           n13500, C1 => n14602, C2 => n13497, ZN => n11007);
   U2324 : OAI222_X1 port map( A1 => n14854, A2 => n13503, B1 => n1234, B2 => 
                           n13500, C1 => n14596, C2 => n13497, ZN => n11006);
   U2325 : OAI222_X1 port map( A1 => n14848, A2 => n13503, B1 => n1233, B2 => 
                           n13500, C1 => n14590, C2 => n13497, ZN => n11005);
   U2326 : OAI222_X1 port map( A1 => n14842, A2 => n13503, B1 => n1232, B2 => 
                           n13500, C1 => n14584, C2 => n13497, ZN => n11004);
   U2327 : OAI222_X1 port map( A1 => n14836, A2 => n13503, B1 => n1231, B2 => 
                           n13500, C1 => n14578, C2 => n13497, ZN => n11003);
   U2328 : OAI222_X1 port map( A1 => n14830, A2 => n13503, B1 => n1230, B2 => 
                           n13500, C1 => n14572, C2 => n13497, ZN => n11002);
   U2329 : OAI222_X1 port map( A1 => n14824, A2 => n13503, B1 => n1229, B2 => 
                           n13500, C1 => n14566, C2 => n13497, ZN => n11001);
   U2330 : OAI222_X1 port map( A1 => n14818, A2 => n13502, B1 => n1228, B2 => 
                           n13499, C1 => n14560, C2 => n13497, ZN => n11000);
   U2331 : OAI222_X1 port map( A1 => n14812, A2 => n13502, B1 => n1227, B2 => 
                           n13499, C1 => n14554, C2 => n13496, ZN => n10999);
   U2332 : OAI222_X1 port map( A1 => n14806, A2 => n13502, B1 => n1226, B2 => 
                           n13499, C1 => n14548, C2 => n13496, ZN => n10998);
   U2333 : OAI222_X1 port map( A1 => n14800, A2 => n13502, B1 => n1225, B2 => 
                           n13499, C1 => n14542, C2 => n13496, ZN => n10997);
   U2334 : OAI222_X1 port map( A1 => n14794, A2 => n13502, B1 => n1224, B2 => 
                           n13499, C1 => n14536, C2 => n13496, ZN => n10996);
   U2335 : OAI222_X1 port map( A1 => n14788, A2 => n13502, B1 => n1223, B2 => 
                           n13499, C1 => n14530, C2 => n13496, ZN => n10995);
   U2336 : OAI222_X1 port map( A1 => n14782, A2 => n13502, B1 => n1222, B2 => 
                           n13499, C1 => n14524, C2 => n13496, ZN => n10994);
   U2337 : OAI222_X1 port map( A1 => n14776, A2 => n13502, B1 => n1221, B2 => 
                           n13499, C1 => n14518, C2 => n13496, ZN => n10993);
   U2338 : OAI222_X1 port map( A1 => n14770, A2 => n13502, B1 => n1220, B2 => 
                           n13499, C1 => n14512, C2 => n13496, ZN => n10992);
   U2339 : OAI222_X1 port map( A1 => n14764, A2 => n13502, B1 => n1219, B2 => 
                           n13499, C1 => n14713, C2 => n13496, ZN => n10991);
   U2340 : OAI222_X1 port map( A1 => n14758, A2 => n13502, B1 => n1218, B2 => 
                           n13499, C1 => n14701, C2 => n13496, ZN => n10990);
   U2341 : OAI222_X1 port map( A1 => n14752, A2 => n13502, B1 => n1217, B2 => 
                           n13499, C1 => n14694, C2 => n13496, ZN => n10989);
   U2342 : OAI222_X1 port map( A1 => n14884, A2 => n13512, B1 => n1215, B2 => 
                           n13509, C1 => n14626, C2 => n13506, ZN => n11043);
   U2343 : OAI222_X1 port map( A1 => n14878, A2 => n13512, B1 => n1214, B2 => 
                           n13509, C1 => n14620, C2 => n13506, ZN => n11042);
   U2344 : OAI222_X1 port map( A1 => n14872, A2 => n13512, B1 => n1213, B2 => 
                           n13509, C1 => n14614, C2 => n13506, ZN => n11041);
   U2345 : OAI222_X1 port map( A1 => n14866, A2 => n13512, B1 => n1212, B2 => 
                           n13509, C1 => n14608, C2 => n13506, ZN => n11040);
   U2346 : OAI222_X1 port map( A1 => n14860, A2 => n13512, B1 => n1211, B2 => 
                           n13509, C1 => n14602, C2 => n13506, ZN => n11039);
   U2347 : OAI222_X1 port map( A1 => n14854, A2 => n13512, B1 => n1210, B2 => 
                           n13509, C1 => n14596, C2 => n13506, ZN => n11038);
   U2348 : OAI222_X1 port map( A1 => n14848, A2 => n13512, B1 => n1209, B2 => 
                           n13509, C1 => n14590, C2 => n13506, ZN => n11037);
   U2349 : OAI222_X1 port map( A1 => n14842, A2 => n13512, B1 => n1208, B2 => 
                           n13509, C1 => n14584, C2 => n13506, ZN => n11036);
   U2350 : OAI222_X1 port map( A1 => n14836, A2 => n13512, B1 => n1207, B2 => 
                           n13509, C1 => n14578, C2 => n13506, ZN => n11035);
   U2351 : OAI222_X1 port map( A1 => n14830, A2 => n13512, B1 => n1206, B2 => 
                           n13509, C1 => n14572, C2 => n13506, ZN => n11034);
   U2352 : OAI222_X1 port map( A1 => n14824, A2 => n13512, B1 => n1205, B2 => 
                           n13509, C1 => n14566, C2 => n13506, ZN => n11033);
   U2353 : OAI222_X1 port map( A1 => n14818, A2 => n13511, B1 => n1204, B2 => 
                           n13508, C1 => n14560, C2 => n13506, ZN => n11032);
   U2354 : OAI222_X1 port map( A1 => n14812, A2 => n13511, B1 => n1203, B2 => 
                           n13508, C1 => n14554, C2 => n13505, ZN => n11031);
   U2355 : OAI222_X1 port map( A1 => n14806, A2 => n13511, B1 => n1202, B2 => 
                           n13508, C1 => n14548, C2 => n13505, ZN => n11030);
   U2356 : OAI222_X1 port map( A1 => n14800, A2 => n13511, B1 => n1201, B2 => 
                           n13508, C1 => n14542, C2 => n13505, ZN => n11029);
   U2357 : OAI222_X1 port map( A1 => n14794, A2 => n13511, B1 => n1200, B2 => 
                           n13508, C1 => n14536, C2 => n13505, ZN => n11028);
   U2358 : OAI222_X1 port map( A1 => n14788, A2 => n13511, B1 => n1199, B2 => 
                           n13508, C1 => n14530, C2 => n13505, ZN => n11027);
   U2359 : OAI222_X1 port map( A1 => n14782, A2 => n13511, B1 => n1198, B2 => 
                           n13508, C1 => n14524, C2 => n13505, ZN => n11026);
   U2360 : OAI222_X1 port map( A1 => n14776, A2 => n13511, B1 => n1197, B2 => 
                           n13508, C1 => n14518, C2 => n13505, ZN => n11025);
   U2361 : OAI222_X1 port map( A1 => n14770, A2 => n13511, B1 => n1196, B2 => 
                           n13508, C1 => n14512, C2 => n13505, ZN => n11024);
   U2362 : OAI222_X1 port map( A1 => n14764, A2 => n13511, B1 => n1195, B2 => 
                           n13508, C1 => n14713, C2 => n13505, ZN => n11023);
   U2363 : OAI222_X1 port map( A1 => n14758, A2 => n13511, B1 => n1194, B2 => 
                           n13508, C1 => n14701, C2 => n13505, ZN => n11022);
   U2364 : OAI222_X1 port map( A1 => n14752, A2 => n13511, B1 => n1193, B2 => 
                           n13508, C1 => n14694, C2 => n13505, ZN => n11021);
   U2365 : OAI222_X1 port map( A1 => n14884, A2 => n13548, B1 => n1143, B2 => 
                           n13545, C1 => n14625, C2 => n13542, ZN => n11171);
   U2366 : OAI222_X1 port map( A1 => n14878, A2 => n13548, B1 => n1142, B2 => 
                           n13545, C1 => n14619, C2 => n13542, ZN => n11170);
   U2367 : OAI222_X1 port map( A1 => n14872, A2 => n13548, B1 => n1141, B2 => 
                           n13545, C1 => n14613, C2 => n13542, ZN => n11169);
   U2368 : OAI222_X1 port map( A1 => n14866, A2 => n13548, B1 => n1140, B2 => 
                           n13545, C1 => n14607, C2 => n13542, ZN => n11168);
   U2369 : OAI222_X1 port map( A1 => n14860, A2 => n13548, B1 => n1139, B2 => 
                           n13545, C1 => n14601, C2 => n13542, ZN => n11167);
   U2370 : OAI222_X1 port map( A1 => n14854, A2 => n13548, B1 => n1138, B2 => 
                           n13545, C1 => n14595, C2 => n13542, ZN => n11166);
   U2371 : OAI222_X1 port map( A1 => n14848, A2 => n13548, B1 => n1137, B2 => 
                           n13545, C1 => n14589, C2 => n13542, ZN => n11165);
   U2372 : OAI222_X1 port map( A1 => n14842, A2 => n13548, B1 => n1136, B2 => 
                           n13545, C1 => n14583, C2 => n13542, ZN => n11164);
   U2373 : OAI222_X1 port map( A1 => n14836, A2 => n13548, B1 => n1135, B2 => 
                           n13545, C1 => n14577, C2 => n13542, ZN => n11163);
   U2374 : OAI222_X1 port map( A1 => n14859, A2 => n13557, B1 => n1134, B2 => 
                           n13554, C1 => n14601, C2 => n13551, ZN => n11199);
   U2375 : OAI222_X1 port map( A1 => n14853, A2 => n13557, B1 => n1133, B2 => 
                           n13554, C1 => n14595, C2 => n13551, ZN => n11198);
   U2376 : OAI222_X1 port map( A1 => n14847, A2 => n13557, B1 => n1132, B2 => 
                           n13554, C1 => n14589, C2 => n13551, ZN => n11197);
   U2377 : OAI222_X1 port map( A1 => n14841, A2 => n13557, B1 => n1131, B2 => 
                           n13554, C1 => n14583, C2 => n13551, ZN => n11196);
   U2378 : OAI222_X1 port map( A1 => n14835, A2 => n13557, B1 => n1130, B2 => 
                           n13554, C1 => n14577, C2 => n13551, ZN => n11195);
   U2379 : OAI222_X1 port map( A1 => n14883, A2 => n13566, B1 => n1128, B2 => 
                           n13563, C1 => n14625, C2 => n13560, ZN => n11235);
   U2380 : OAI222_X1 port map( A1 => n14877, A2 => n13566, B1 => n1127, B2 => 
                           n13563, C1 => n14619, C2 => n13560, ZN => n11234);
   U2381 : OAI222_X1 port map( A1 => n14871, A2 => n13566, B1 => n1126, B2 => 
                           n13563, C1 => n14613, C2 => n13560, ZN => n11233);
   U2382 : OAI222_X1 port map( A1 => n14865, A2 => n13566, B1 => n1125, B2 => 
                           n13563, C1 => n14607, C2 => n13560, ZN => n11232);
   U2383 : OAI222_X1 port map( A1 => n14859, A2 => n13566, B1 => n1124, B2 => 
                           n13563, C1 => n14601, C2 => n13560, ZN => n11231);
   U2384 : OAI222_X1 port map( A1 => n14853, A2 => n13566, B1 => n1123, B2 => 
                           n13563, C1 => n14595, C2 => n13560, ZN => n11230);
   U2385 : OAI222_X1 port map( A1 => n14847, A2 => n13566, B1 => n1122, B2 => 
                           n13563, C1 => n14589, C2 => n13560, ZN => n11229);
   U2386 : OAI222_X1 port map( A1 => n14841, A2 => n13566, B1 => n1121, B2 => 
                           n13563, C1 => n14583, C2 => n13560, ZN => n11228);
   U2387 : OAI222_X1 port map( A1 => n14835, A2 => n13566, B1 => n1120, B2 => 
                           n13563, C1 => n14577, C2 => n13560, ZN => n11227);
   U2388 : OAI222_X1 port map( A1 => n14829, A2 => n13566, B1 => n1119, B2 => 
                           n13563, C1 => n14571, C2 => n13560, ZN => n11226);
   U2389 : OAI222_X1 port map( A1 => n14823, A2 => n13566, B1 => n1118, B2 => 
                           n13563, C1 => n14565, C2 => n13560, ZN => n11225);
   U2390 : OAI222_X1 port map( A1 => n14817, A2 => n13565, B1 => n1117, B2 => 
                           n13562, C1 => n14559, C2 => n13560, ZN => n11224);
   U2391 : OAI222_X1 port map( A1 => n14811, A2 => n13565, B1 => n1116, B2 => 
                           n13562, C1 => n14553, C2 => n13559, ZN => n11223);
   U2392 : OAI222_X1 port map( A1 => n14805, A2 => n13565, B1 => n1115, B2 => 
                           n13562, C1 => n14547, C2 => n13559, ZN => n11222);
   U2393 : OAI222_X1 port map( A1 => n14799, A2 => n13565, B1 => n1114, B2 => 
                           n13562, C1 => n14541, C2 => n13559, ZN => n11221);
   U2394 : OAI222_X1 port map( A1 => n14793, A2 => n13565, B1 => n1113, B2 => 
                           n13562, C1 => n14535, C2 => n13559, ZN => n11220);
   U2395 : OAI222_X1 port map( A1 => n14787, A2 => n13565, B1 => n1112, B2 => 
                           n13562, C1 => n14529, C2 => n13559, ZN => n11219);
   U2396 : OAI222_X1 port map( A1 => n14781, A2 => n13565, B1 => n1111, B2 => 
                           n13562, C1 => n14523, C2 => n13559, ZN => n11218);
   U2397 : OAI222_X1 port map( A1 => n14775, A2 => n13565, B1 => n1110, B2 => 
                           n13562, C1 => n14517, C2 => n13559, ZN => n11217);
   U2398 : OAI222_X1 port map( A1 => n14769, A2 => n13565, B1 => n1109, B2 => 
                           n13562, C1 => n14511, C2 => n13559, ZN => n11216);
   U2399 : OAI222_X1 port map( A1 => n14763, A2 => n13565, B1 => n1108, B2 => 
                           n13562, C1 => n14712, C2 => n13559, ZN => n11215);
   U2400 : OAI222_X1 port map( A1 => n14757, A2 => n13565, B1 => n1107, B2 => 
                           n13562, C1 => n14700, C2 => n13559, ZN => n11214);
   U2401 : OAI222_X1 port map( A1 => n14751, A2 => n13565, B1 => n1106, B2 => 
                           n13562, C1 => n14695, C2 => n13559, ZN => n11213);
   U2402 : OAI222_X1 port map( A1 => n14892, A2 => n13242, B1 => n1105, B2 => 
                           n13239, C1 => n14634, C2 => n13236, ZN => n10084);
   U2403 : OAI222_X1 port map( A1 => n14886, A2 => n13242, B1 => n1104, B2 => 
                           n13239, C1 => n14628, C2 => n13236, ZN => n10083);
   U2404 : OAI222_X1 port map( A1 => n14880, A2 => n13242, B1 => n1103, B2 => 
                           n13239, C1 => n14622, C2 => n13236, ZN => n10082);
   U2405 : OAI222_X1 port map( A1 => n14874, A2 => n13242, B1 => n1102, B2 => 
                           n13239, C1 => n14616, C2 => n13236, ZN => n10081);
   U2406 : OAI222_X1 port map( A1 => n14868, A2 => n13242, B1 => n1101, B2 => 
                           n13239, C1 => n14610, C2 => n13236, ZN => n10080);
   U2407 : OAI222_X1 port map( A1 => n14862, A2 => n13242, B1 => n1100, B2 => 
                           n13239, C1 => n14604, C2 => n13236, ZN => n10079);
   U2408 : OAI222_X1 port map( A1 => n14856, A2 => n13242, B1 => n1099, B2 => 
                           n13239, C1 => n14598, C2 => n13236, ZN => n10078);
   U2409 : OAI222_X1 port map( A1 => n14850, A2 => n13242, B1 => n1098, B2 => 
                           n13239, C1 => n14592, C2 => n13236, ZN => n10077);
   U2410 : OAI222_X1 port map( A1 => n14844, A2 => n13242, B1 => n1097, B2 => 
                           n13239, C1 => n14586, C2 => n13236, ZN => n10076);
   U2411 : OAI222_X1 port map( A1 => n14838, A2 => n13242, B1 => n1096, B2 => 
                           n13239, C1 => n14580, C2 => n13236, ZN => n10075);
   U2412 : OAI222_X1 port map( A1 => n14832, A2 => n13242, B1 => n1095, B2 => 
                           n13239, C1 => n14574, C2 => n13236, ZN => n10074);
   U2413 : OAI222_X1 port map( A1 => n14820, A2 => n13241, B1 => n1094, B2 => 
                           n13238, C1 => n14562, C2 => n13236, ZN => n10072);
   U2414 : OAI222_X1 port map( A1 => n14814, A2 => n13241, B1 => n1093, B2 => 
                           n13238, C1 => n14556, C2 => n13235, ZN => n10071);
   U2415 : OAI222_X1 port map( A1 => n14808, A2 => n13241, B1 => n1092, B2 => 
                           n13238, C1 => n14550, C2 => n13235, ZN => n10070);
   U2416 : OAI222_X1 port map( A1 => n14802, A2 => n13241, B1 => n1091, B2 => 
                           n13238, C1 => n14544, C2 => n13235, ZN => n10069);
   U2417 : OAI222_X1 port map( A1 => n14796, A2 => n13241, B1 => n1090, B2 => 
                           n13238, C1 => n14538, C2 => n13235, ZN => n10068);
   U2418 : OAI222_X1 port map( A1 => n14790, A2 => n13241, B1 => n1089, B2 => 
                           n13238, C1 => n14532, C2 => n13235, ZN => n10067);
   U2419 : OAI222_X1 port map( A1 => n14784, A2 => n13241, B1 => n1088, B2 => 
                           n13238, C1 => n14526, C2 => n13235, ZN => n10066);
   U2420 : OAI222_X1 port map( A1 => n14778, A2 => n13241, B1 => n1087, B2 => 
                           n13238, C1 => n14520, C2 => n13235, ZN => n10065);
   U2421 : OAI222_X1 port map( A1 => n14761, A2 => n13241, B1 => n1086, B2 => 
                           n13238, C1 => n14715, C2 => n13235, ZN => n10063);
   U2422 : OAI222_X1 port map( A1 => n14755, A2 => n13241, B1 => n1085, B2 => 
                           n13238, C1 => n14703, C2 => n13235, ZN => n10062);
   U2423 : OAI222_X1 port map( A1 => n14892, A2 => n13251, B1 => n1084, B2 => 
                           n13248, C1 => n14634, C2 => n13245, ZN => n10116);
   U2424 : OAI222_X1 port map( A1 => n14886, A2 => n13251, B1 => n1083, B2 => 
                           n13248, C1 => n14628, C2 => n13245, ZN => n10115);
   U2425 : OAI222_X1 port map( A1 => n14880, A2 => n13251, B1 => n1082, B2 => 
                           n13248, C1 => n14622, C2 => n13245, ZN => n10114);
   U2426 : OAI222_X1 port map( A1 => n14874, A2 => n13251, B1 => n1081, B2 => 
                           n13248, C1 => n14616, C2 => n13245, ZN => n10113);
   U2427 : OAI222_X1 port map( A1 => n14868, A2 => n13251, B1 => n1080, B2 => 
                           n13248, C1 => n14610, C2 => n13245, ZN => n10112);
   U2428 : OAI222_X1 port map( A1 => n14862, A2 => n13251, B1 => n1079, B2 => 
                           n13248, C1 => n14604, C2 => n13245, ZN => n10111);
   U2429 : OAI222_X1 port map( A1 => n14856, A2 => n13251, B1 => n1078, B2 => 
                           n13248, C1 => n14598, C2 => n13245, ZN => n10110);
   U2430 : OAI222_X1 port map( A1 => n14850, A2 => n13251, B1 => n1077, B2 => 
                           n13248, C1 => n14592, C2 => n13245, ZN => n10109);
   U2431 : OAI222_X1 port map( A1 => n14844, A2 => n13251, B1 => n1076, B2 => 
                           n13248, C1 => n14586, C2 => n13245, ZN => n10108);
   U2432 : OAI222_X1 port map( A1 => n14838, A2 => n13251, B1 => n1075, B2 => 
                           n13248, C1 => n14580, C2 => n13245, ZN => n10107);
   U2433 : OAI222_X1 port map( A1 => n14832, A2 => n13251, B1 => n1074, B2 => 
                           n13248, C1 => n14574, C2 => n13245, ZN => n10106);
   U2434 : OAI222_X1 port map( A1 => n14820, A2 => n13250, B1 => n1073, B2 => 
                           n13247, C1 => n14562, C2 => n13245, ZN => n10104);
   U2435 : OAI222_X1 port map( A1 => n14814, A2 => n13250, B1 => n1072, B2 => 
                           n13247, C1 => n14556, C2 => n13244, ZN => n10103);
   U2436 : OAI222_X1 port map( A1 => n14808, A2 => n13250, B1 => n1071, B2 => 
                           n13247, C1 => n14550, C2 => n13244, ZN => n10102);
   U2437 : OAI222_X1 port map( A1 => n14802, A2 => n13250, B1 => n1070, B2 => 
                           n13247, C1 => n14544, C2 => n13244, ZN => n10101);
   U2438 : OAI222_X1 port map( A1 => n14796, A2 => n13250, B1 => n1069, B2 => 
                           n13247, C1 => n14538, C2 => n13244, ZN => n10100);
   U2439 : OAI222_X1 port map( A1 => n14790, A2 => n13250, B1 => n1068, B2 => 
                           n13247, C1 => n14532, C2 => n13244, ZN => n10099);
   U2440 : OAI222_X1 port map( A1 => n14784, A2 => n13250, B1 => n1067, B2 => 
                           n13247, C1 => n14526, C2 => n13244, ZN => n10098);
   U2441 : OAI222_X1 port map( A1 => n14778, A2 => n13250, B1 => n1066, B2 => 
                           n13247, C1 => n14520, C2 => n13244, ZN => n10097);
   U2442 : OAI222_X1 port map( A1 => n14772, A2 => n13250, B1 => n1065, B2 => 
                           n13247, C1 => n14514, C2 => n13244, ZN => n10096);
   U2443 : OAI222_X1 port map( A1 => n14766, A2 => n13250, B1 => n1064, B2 => 
                           n13247, C1 => n14715, C2 => n13244, ZN => n10095);
   U2444 : OAI222_X1 port map( A1 => n14760, A2 => n13250, B1 => n1063, B2 => 
                           n13247, C1 => n14703, C2 => n13244, ZN => n10094);
   U2445 : OAI222_X1 port map( A1 => n14754, A2 => n13250, B1 => n1062, B2 => 
                           n13247, C1 => n14692, C2 => n13244, ZN => n10093);
   U2446 : OAI222_X1 port map( A1 => n14754, A2 => n13268, B1 => n1061, B2 => 
                           n13265, C1 => n14692, C2 => n13262, ZN => n10157);
   U2447 : OAI222_X1 port map( A1 => n14882, A2 => n14352, B1 => n14348, B2 => 
                           n1011, C1 => n14625, C2 => n14346, ZN => n9411);
   U2448 : OAI222_X1 port map( A1 => n14876, A2 => n14352, B1 => n14348, B2 => 
                           n1010, C1 => n14619, C2 => n14346, ZN => n9410);
   U2449 : OAI222_X1 port map( A1 => n14870, A2 => n14352, B1 => n14348, B2 => 
                           n1009, C1 => n14613, C2 => n14346, ZN => n9409);
   U2450 : OAI222_X1 port map( A1 => n14864, A2 => n14352, B1 => n14349, B2 => 
                           n1008, C1 => n14607, C2 => n14346, ZN => n9408);
   U2451 : OAI222_X1 port map( A1 => n14858, A2 => n14352, B1 => n14349, B2 => 
                           n1007, C1 => n14601, C2 => n14346, ZN => n9407);
   U2452 : OAI222_X1 port map( A1 => n14852, A2 => n14352, B1 => n14349, B2 => 
                           n1006, C1 => n14595, C2 => n14346, ZN => n9406);
   U2453 : OAI222_X1 port map( A1 => n14846, A2 => n14352, B1 => n14349, B2 => 
                           n1005, C1 => n14589, C2 => n14346, ZN => n9405);
   U2454 : OAI222_X1 port map( A1 => n14840, A2 => n14352, B1 => n14349, B2 => 
                           n1004, C1 => n14583, C2 => n14346, ZN => n9404);
   U2455 : OAI222_X1 port map( A1 => n14834, A2 => n14352, B1 => n14349, B2 => 
                           n1003, C1 => n14577, C2 => n14346, ZN => n9403);
   U2456 : OAI222_X1 port map( A1 => n14828, A2 => n14352, B1 => n14349, B2 => 
                           n1002, C1 => n14571, C2 => n14346, ZN => n9402);
   U2457 : OAI222_X1 port map( A1 => n14810, A2 => n14351, B1 => n14349, B2 => 
                           n996, C1 => n14553, C2 => n14345, ZN => n9399);
   U2458 : OAI222_X1 port map( A1 => n14804, A2 => n14351, B1 => n14349, B2 => 
                           n994, C1 => n14547, C2 => n14345, ZN => n9398);
   U2459 : OAI222_X1 port map( A1 => n14798, A2 => n14351, B1 => n14349, B2 => 
                           n990, C1 => n14541, C2 => n14345, ZN => n9397);
   U2460 : OAI222_X1 port map( A1 => n14792, A2 => n14351, B1 => n14349, B2 => 
                           n988, C1 => n14535, C2 => n14345, ZN => n9396);
   U2461 : OAI222_X1 port map( A1 => n14786, A2 => n14351, B1 => n14350, B2 => 
                           n984, C1 => n14529, C2 => n14345, ZN => n9395);
   U2462 : OAI222_X1 port map( A1 => n14780, A2 => n14351, B1 => n14350, B2 => 
                           n982, C1 => n14523, C2 => n14345, ZN => n9394);
   U2463 : OAI222_X1 port map( A1 => n14774, A2 => n14351, B1 => n14350, B2 => 
                           n978, C1 => n14517, C2 => n14345, ZN => n9393);
   U2464 : OAI222_X1 port map( A1 => n14768, A2 => n14351, B1 => n14350, B2 => 
                           n976, C1 => n14511, C2 => n14345, ZN => n9392);
   U2465 : OAI222_X1 port map( A1 => n14762, A2 => n14351, B1 => n14350, B2 => 
                           n972, C1 => n14711, C2 => n14345, ZN => n9391);
   U2466 : OAI222_X1 port map( A1 => n14756, A2 => n14351, B1 => n14350, B2 => 
                           n970, C1 => n14699, C2 => n14345, ZN => n9390);
   U2467 : OAI222_X1 port map( A1 => n14750, A2 => n14351, B1 => n14348, B2 => 
                           n966, C1 => n14696, C2 => n14345, ZN => n9389);
   U2468 : OAI222_X1 port map( A1 => n14888, A2 => n14372, B1 => n14369, B2 => 
                           n964, C1 => n14630, C2 => n14366, ZN => n9476);
   U2469 : OAI222_X1 port map( A1 => n14882, A2 => n14372, B1 => n14369, B2 => 
                           n960, C1 => n14624, C2 => n14366, ZN => n9475);
   U2470 : OAI222_X1 port map( A1 => n14876, A2 => n14372, B1 => n14369, B2 => 
                           n958, C1 => n14618, C2 => n14366, ZN => n9474);
   U2471 : OAI222_X1 port map( A1 => n14870, A2 => n14372, B1 => n14369, B2 => 
                           n954, C1 => n14612, C2 => n14366, ZN => n9473);
   U2472 : OAI222_X1 port map( A1 => n14864, A2 => n14372, B1 => n14369, B2 => 
                           n952, C1 => n14606, C2 => n14366, ZN => n9472);
   U2473 : OAI222_X1 port map( A1 => n14858, A2 => n14372, B1 => n14369, B2 => 
                           n948, C1 => n14600, C2 => n14366, ZN => n9471);
   U2474 : OAI222_X1 port map( A1 => n14852, A2 => n14372, B1 => n14369, B2 => 
                           n946, C1 => n14594, C2 => n14366, ZN => n9470);
   U2475 : OAI222_X1 port map( A1 => n14846, A2 => n14372, B1 => n14369, B2 => 
                           n942, C1 => n14588, C2 => n14366, ZN => n9469);
   U2476 : OAI222_X1 port map( A1 => n14840, A2 => n14372, B1 => n14369, B2 => 
                           n940, C1 => n14582, C2 => n14366, ZN => n9468);
   U2477 : OAI222_X1 port map( A1 => n14834, A2 => n14372, B1 => n14369, B2 => 
                           n936, C1 => n14576, C2 => n14366, ZN => n9467);
   U2478 : OAI222_X1 port map( A1 => n14828, A2 => n14372, B1 => n14369, B2 => 
                           n934, C1 => n14570, C2 => n14366, ZN => n9466);
   U2479 : OAI222_X1 port map( A1 => n14822, A2 => n14372, B1 => n14369, B2 => 
                           n930, C1 => n14564, C2 => n14366, ZN => n9465);
   U2480 : OAI222_X1 port map( A1 => n14816, A2 => n14371, B1 => n14368, B2 => 
                           n928, C1 => n14558, C2 => n14366, ZN => n9464);
   U2481 : OAI222_X1 port map( A1 => n14810, A2 => n14371, B1 => n14368, B2 => 
                           n924, C1 => n14552, C2 => n14365, ZN => n9463);
   U2482 : OAI222_X1 port map( A1 => n14804, A2 => n14371, B1 => n14368, B2 => 
                           n922, C1 => n14546, C2 => n14365, ZN => n9462);
   U2483 : OAI222_X1 port map( A1 => n14798, A2 => n14371, B1 => n14368, B2 => 
                           n918, C1 => n14540, C2 => n14365, ZN => n9461);
   U2484 : OAI222_X1 port map( A1 => n14792, A2 => n14371, B1 => n14368, B2 => 
                           n916, C1 => n14534, C2 => n14365, ZN => n9460);
   U2485 : OAI222_X1 port map( A1 => n14786, A2 => n14371, B1 => n14368, B2 => 
                           n912, C1 => n14528, C2 => n14365, ZN => n9459);
   U2486 : OAI222_X1 port map( A1 => n14780, A2 => n14371, B1 => n14368, B2 => 
                           n910, C1 => n14522, C2 => n14365, ZN => n9458);
   U2487 : OAI222_X1 port map( A1 => n14774, A2 => n14371, B1 => n14368, B2 => 
                           n906, C1 => n14516, C2 => n14365, ZN => n9457);
   U2488 : OAI222_X1 port map( A1 => n14768, A2 => n14371, B1 => n14368, B2 => 
                           n904, C1 => n14510, C2 => n14365, ZN => n9456);
   U2489 : OAI222_X1 port map( A1 => n14762, A2 => n14371, B1 => n14368, B2 => 
                           n900, C1 => n14711, C2 => n14365, ZN => n9455);
   U2490 : OAI222_X1 port map( A1 => n14756, A2 => n14371, B1 => n14368, B2 => 
                           n898, C1 => n14699, C2 => n14365, ZN => n9454);
   U2491 : OAI222_X1 port map( A1 => n14750, A2 => n14371, B1 => n14368, B2 => 
                           n819, C1 => n14696, C2 => n14365, ZN => n9453);
   U2492 : OAI222_X1 port map( A1 => n14882, A2 => n14381, B1 => n14377, B2 => 
                           n809, C1 => n14624, C2 => n14375, ZN => n9507);
   U2493 : OAI222_X1 port map( A1 => n14876, A2 => n14381, B1 => n14377, B2 => 
                           n808, C1 => n14618, C2 => n14375, ZN => n9506);
   U2494 : OAI222_X1 port map( A1 => n14870, A2 => n14381, B1 => n14377, B2 => 
                           n804, C1 => n14612, C2 => n14375, ZN => n9505);
   U2495 : OAI222_X1 port map( A1 => n14864, A2 => n14381, B1 => n14378, B2 => 
                           n797, C1 => n14606, C2 => n14375, ZN => n9504);
   U2496 : OAI222_X1 port map( A1 => n14858, A2 => n14381, B1 => n14378, B2 => 
                           n796, C1 => n14600, C2 => n14375, ZN => n9503);
   U2497 : OAI222_X1 port map( A1 => n14852, A2 => n14381, B1 => n14378, B2 => 
                           n794, C1 => n14594, C2 => n14375, ZN => n9502);
   U2498 : OAI222_X1 port map( A1 => n14846, A2 => n14381, B1 => n14378, B2 => 
                           n793, C1 => n14588, C2 => n14375, ZN => n9501);
   U2499 : OAI222_X1 port map( A1 => n14840, A2 => n14381, B1 => n14378, B2 => 
                           n792, C1 => n14582, C2 => n14375, ZN => n9500);
   U2500 : OAI222_X1 port map( A1 => n14834, A2 => n14381, B1 => n14378, B2 => 
                           n790, C1 => n14576, C2 => n14375, ZN => n9499);
   U2501 : OAI222_X1 port map( A1 => n14828, A2 => n14381, B1 => n14378, B2 => 
                           n789, C1 => n14570, C2 => n14375, ZN => n9498);
   U2502 : OAI222_X1 port map( A1 => n14816, A2 => n14380, B1 => n14378, B2 => 
                           n787, C1 => n14558, C2 => n14375, ZN => n9496);
   U2503 : OAI222_X1 port map( A1 => n14810, A2 => n14380, B1 => n14378, B2 => 
                           n785, C1 => n14552, C2 => n14374, ZN => n9495);
   U2504 : OAI222_X1 port map( A1 => n14804, A2 => n14380, B1 => n14378, B2 => 
                           n783, C1 => n14546, C2 => n14374, ZN => n9494);
   U2505 : OAI222_X1 port map( A1 => n14798, A2 => n14380, B1 => n14378, B2 => 
                           n782, C1 => n14540, C2 => n14374, ZN => n9493);
   U2506 : OAI222_X1 port map( A1 => n14792, A2 => n14380, B1 => n14379, B2 => 
                           n781, C1 => n14534, C2 => n14374, ZN => n9492);
   U2507 : OAI222_X1 port map( A1 => n14786, A2 => n14380, B1 => n14379, B2 => 
                           n780, C1 => n14528, C2 => n14374, ZN => n9491);
   U2508 : OAI222_X1 port map( A1 => n14780, A2 => n14380, B1 => n14379, B2 => 
                           n779, C1 => n14522, C2 => n14374, ZN => n9490);
   U2509 : OAI222_X1 port map( A1 => n14774, A2 => n14380, B1 => n14379, B2 => 
                           n778, C1 => n14516, C2 => n14374, ZN => n9489);
   U2510 : OAI222_X1 port map( A1 => n14768, A2 => n14380, B1 => n14379, B2 => 
                           n776, C1 => n14510, C2 => n14374, ZN => n9488);
   U2511 : OAI222_X1 port map( A1 => n14762, A2 => n14380, B1 => n14379, B2 => 
                           n775, C1 => n14711, C2 => n14374, ZN => n9487);
   U2512 : OAI222_X1 port map( A1 => n14756, A2 => n14380, B1 => n14379, B2 => 
                           n773, C1 => n14699, C2 => n14374, ZN => n9486);
   U2513 : OAI222_X1 port map( A1 => n14750, A2 => n14380, B1 => n14377, B2 => 
                           n772, C1 => n14696, C2 => n14374, ZN => n9485);
   U2514 : OAI222_X1 port map( A1 => n14889, A2 => n13575, B1 => n771, B2 => 
                           n13572, C1 => n14631, C2 => n13569, ZN => n11268);
   U2515 : OAI222_X1 port map( A1 => n14883, A2 => n13575, B1 => n769, B2 => 
                           n13572, C1 => n14625, C2 => n13569, ZN => n11267);
   U2516 : OAI222_X1 port map( A1 => n14877, A2 => n13575, B1 => n768, B2 => 
                           n13572, C1 => n14619, C2 => n13569, ZN => n11266);
   U2517 : OAI222_X1 port map( A1 => n14871, A2 => n13575, B1 => n767, B2 => 
                           n13572, C1 => n14613, C2 => n13569, ZN => n11265);
   U2518 : OAI222_X1 port map( A1 => n14865, A2 => n13575, B1 => n766, B2 => 
                           n13572, C1 => n14607, C2 => n13569, ZN => n11264);
   U2519 : OAI222_X1 port map( A1 => n14859, A2 => n13575, B1 => n765, B2 => 
                           n13572, C1 => n14601, C2 => n13569, ZN => n11263);
   U2520 : OAI222_X1 port map( A1 => n14853, A2 => n13575, B1 => n764, B2 => 
                           n13572, C1 => n14595, C2 => n13569, ZN => n11262);
   U2521 : OAI222_X1 port map( A1 => n14847, A2 => n13575, B1 => n760, B2 => 
                           n13572, C1 => n14589, C2 => n13569, ZN => n11261);
   U2522 : OAI222_X1 port map( A1 => n14841, A2 => n13575, B1 => n759, B2 => 
                           n13572, C1 => n14583, C2 => n13569, ZN => n11260);
   U2523 : OAI222_X1 port map( A1 => n14835, A2 => n13575, B1 => n758, B2 => 
                           n13572, C1 => n14577, C2 => n13569, ZN => n11259);
   U2524 : OAI222_X1 port map( A1 => n14829, A2 => n13575, B1 => n757, B2 => 
                           n13572, C1 => n14571, C2 => n13569, ZN => n11258);
   U2525 : OAI222_X1 port map( A1 => n14823, A2 => n13575, B1 => n755, B2 => 
                           n13572, C1 => n14565, C2 => n13569, ZN => n11257);
   U2526 : OAI222_X1 port map( A1 => n14817, A2 => n13574, B1 => n751, B2 => 
                           n13571, C1 => n14559, C2 => n13569, ZN => n11256);
   U2527 : OAI222_X1 port map( A1 => n14811, A2 => n13574, B1 => n750, B2 => 
                           n13571, C1 => n14553, C2 => n13568, ZN => n11255);
   U2528 : OAI222_X1 port map( A1 => n14805, A2 => n13574, B1 => n749, B2 => 
                           n13571, C1 => n14547, C2 => n13568, ZN => n11254);
   U2529 : OAI222_X1 port map( A1 => n14799, A2 => n13574, B1 => n748, B2 => 
                           n13571, C1 => n14541, C2 => n13568, ZN => n11253);
   U2530 : OAI222_X1 port map( A1 => n14793, A2 => n13574, B1 => n747, B2 => 
                           n13571, C1 => n14535, C2 => n13568, ZN => n11252);
   U2531 : OAI222_X1 port map( A1 => n14787, A2 => n13574, B1 => n746, B2 => 
                           n13571, C1 => n14529, C2 => n13568, ZN => n11251);
   U2532 : OAI222_X1 port map( A1 => n14781, A2 => n13574, B1 => n745, B2 => 
                           n13571, C1 => n14523, C2 => n13568, ZN => n11250);
   U2533 : OAI222_X1 port map( A1 => n14775, A2 => n13574, B1 => n744, B2 => 
                           n13571, C1 => n14517, C2 => n13568, ZN => n11249);
   U2534 : OAI222_X1 port map( A1 => n14769, A2 => n13574, B1 => n742, B2 => 
                           n13571, C1 => n14511, C2 => n13568, ZN => n11248);
   U2535 : OAI222_X1 port map( A1 => n14763, A2 => n13574, B1 => n741, B2 => 
                           n13571, C1 => n14712, C2 => n13568, ZN => n11247);
   U2536 : OAI222_X1 port map( A1 => n14757, A2 => n13574, B1 => n740, B2 => 
                           n13571, C1 => n14700, C2 => n13568, ZN => n11246);
   U2537 : OAI222_X1 port map( A1 => n14751, A2 => n13574, B1 => n739, B2 => 
                           n13571, C1 => n14695, C2 => n13568, ZN => n11245);
   U2538 : OAI222_X1 port map( A1 => n14883, A2 => n13584, B1 => n737, B2 => 
                           n13581, C1 => n14625, C2 => n13578, ZN => n11299);
   U2539 : OAI222_X1 port map( A1 => n14877, A2 => n13584, B1 => n733, B2 => 
                           n13581, C1 => n14619, C2 => n13578, ZN => n11298);
   U2540 : OAI222_X1 port map( A1 => n14871, A2 => n13584, B1 => n732, B2 => 
                           n13581, C1 => n14613, C2 => n13578, ZN => n11297);
   U2541 : OAI222_X1 port map( A1 => n14865, A2 => n13584, B1 => n730, B2 => 
                           n13581, C1 => n14607, C2 => n13578, ZN => n11296);
   U2542 : OAI222_X1 port map( A1 => n14859, A2 => n13584, B1 => n729, B2 => 
                           n13581, C1 => n14601, C2 => n13578, ZN => n11295);
   U2543 : OAI222_X1 port map( A1 => n14853, A2 => n13584, B1 => n728, B2 => 
                           n13581, C1 => n14595, C2 => n13578, ZN => n11294);
   U2544 : OAI222_X1 port map( A1 => n14847, A2 => n13584, B1 => n726, B2 => 
                           n13581, C1 => n14589, C2 => n13578, ZN => n11293);
   U2545 : OAI222_X1 port map( A1 => n14841, A2 => n13584, B1 => n725, B2 => 
                           n13581, C1 => n14583, C2 => n13578, ZN => n11292);
   U2546 : OAI222_X1 port map( A1 => n14835, A2 => n13584, B1 => n724, B2 => 
                           n13581, C1 => n14577, C2 => n13578, ZN => n11291);
   U2547 : OAI222_X1 port map( A1 => n14829, A2 => n13584, B1 => n723, B2 => 
                           n13581, C1 => n14571, C2 => n13578, ZN => n11290);
   U2548 : OAI222_X1 port map( A1 => n14823, A2 => n13584, B1 => n722, B2 => 
                           n13581, C1 => n14565, C2 => n13578, ZN => n11289);
   U2549 : OAI222_X1 port map( A1 => n14817, A2 => n13583, B1 => n721, B2 => 
                           n13580, C1 => n14559, C2 => n13578, ZN => n11288);
   U2550 : OAI222_X1 port map( A1 => n14811, A2 => n13583, B1 => n720, B2 => 
                           n13580, C1 => n14553, C2 => n13577, ZN => n11287);
   U2551 : OAI222_X1 port map( A1 => n14805, A2 => n13583, B1 => n719, B2 => 
                           n13580, C1 => n14547, C2 => n13577, ZN => n11286);
   U2552 : OAI222_X1 port map( A1 => n14799, A2 => n13583, B1 => n718, B2 => 
                           n13580, C1 => n14541, C2 => n13577, ZN => n11285);
   U2553 : OAI222_X1 port map( A1 => n14793, A2 => n13583, B1 => n717, B2 => 
                           n13580, C1 => n14535, C2 => n13577, ZN => n11284);
   U2554 : OAI222_X1 port map( A1 => n14787, A2 => n13583, B1 => n716, B2 => 
                           n13580, C1 => n14529, C2 => n13577, ZN => n11283);
   U2555 : OAI222_X1 port map( A1 => n14781, A2 => n13583, B1 => n715, B2 => 
                           n13580, C1 => n14523, C2 => n13577, ZN => n11282);
   U2556 : OAI222_X1 port map( A1 => n14775, A2 => n13583, B1 => n714, B2 => 
                           n13580, C1 => n14517, C2 => n13577, ZN => n11281);
   U2557 : OAI222_X1 port map( A1 => n14769, A2 => n13583, B1 => n713, B2 => 
                           n13580, C1 => n14511, C2 => n13577, ZN => n11280);
   U2558 : OAI222_X1 port map( A1 => n14763, A2 => n13583, B1 => n712, B2 => 
                           n13580, C1 => n14712, C2 => n13577, ZN => n11279);
   U2559 : OAI222_X1 port map( A1 => n14757, A2 => n13583, B1 => n711, B2 => 
                           n13580, C1 => n14700, C2 => n13577, ZN => n11278);
   U2560 : OAI222_X1 port map( A1 => n14751, A2 => n13583, B1 => n710, B2 => 
                           n13580, C1 => n14695, C2 => n13577, ZN => n11277);
   U2561 : OAI222_X1 port map( A1 => n14883, A2 => n13593, B1 => n708, B2 => 
                           n13590, C1 => n14625, C2 => n13587, ZN => n11331);
   U2562 : OAI222_X1 port map( A1 => n14877, A2 => n13593, B1 => n707, B2 => 
                           n13590, C1 => n14619, C2 => n13587, ZN => n11330);
   U2563 : OAI222_X1 port map( A1 => n14871, A2 => n13593, B1 => n706, B2 => 
                           n13590, C1 => n14613, C2 => n13587, ZN => n11329);
   U2564 : OAI222_X1 port map( A1 => n14865, A2 => n13593, B1 => n705, B2 => 
                           n13590, C1 => n14607, C2 => n13587, ZN => n11328);
   U2565 : OAI222_X1 port map( A1 => n14859, A2 => n13593, B1 => n704, B2 => 
                           n13590, C1 => n14601, C2 => n13587, ZN => n11327);
   U2566 : OAI222_X1 port map( A1 => n14853, A2 => n13593, B1 => n703, B2 => 
                           n13590, C1 => n14595, C2 => n13587, ZN => n11326);
   U2567 : OAI222_X1 port map( A1 => n14847, A2 => n13593, B1 => n702, B2 => 
                           n13590, C1 => n14589, C2 => n13587, ZN => n11325);
   U2568 : OAI222_X1 port map( A1 => n14841, A2 => n13593, B1 => n701, B2 => 
                           n13590, C1 => n14583, C2 => n13587, ZN => n11324);
   U2569 : OAI222_X1 port map( A1 => n14835, A2 => n13593, B1 => n700, B2 => 
                           n13590, C1 => n14577, C2 => n13587, ZN => n11323);
   U2570 : OAI222_X1 port map( A1 => n14829, A2 => n13593, B1 => n699, B2 => 
                           n13590, C1 => n14571, C2 => n13587, ZN => n11322);
   U2571 : OAI222_X1 port map( A1 => n14823, A2 => n13593, B1 => n698, B2 => 
                           n13590, C1 => n14565, C2 => n13587, ZN => n11321);
   U2572 : OAI222_X1 port map( A1 => n14805, A2 => n13592, B1 => n695, B2 => 
                           n13589, C1 => n14547, C2 => n13586, ZN => n11318);
   U2573 : OAI222_X1 port map( A1 => n14799, A2 => n13592, B1 => n694, B2 => 
                           n13589, C1 => n14541, C2 => n13586, ZN => n11317);
   U2574 : OAI222_X1 port map( A1 => n14793, A2 => n13592, B1 => n693, B2 => 
                           n13589, C1 => n14535, C2 => n13586, ZN => n11316);
   U2575 : OAI222_X1 port map( A1 => n14787, A2 => n13592, B1 => n692, B2 => 
                           n13589, C1 => n14529, C2 => n13586, ZN => n11315);
   U2576 : OAI222_X1 port map( A1 => n14781, A2 => n13592, B1 => n691, B2 => 
                           n13589, C1 => n14523, C2 => n13586, ZN => n11314);
   U2577 : OAI222_X1 port map( A1 => n14775, A2 => n13592, B1 => n690, B2 => 
                           n13589, C1 => n14517, C2 => n13586, ZN => n11313);
   U2578 : OAI222_X1 port map( A1 => n14769, A2 => n13592, B1 => n689, B2 => 
                           n13589, C1 => n14511, C2 => n13586, ZN => n11312);
   U2579 : OAI222_X1 port map( A1 => n14763, A2 => n13592, B1 => n688, B2 => 
                           n13589, C1 => n14712, C2 => n13586, ZN => n11311);
   U2580 : OAI222_X1 port map( A1 => n14757, A2 => n13592, B1 => n687, B2 => 
                           n13589, C1 => n14700, C2 => n13586, ZN => n11310);
   U2581 : OAI222_X1 port map( A1 => n14751, A2 => n13592, B1 => n686, B2 => 
                           n13589, C1 => n14695, C2 => n13586, ZN => n11309);
   U2582 : OAI222_X1 port map( A1 => n14883, A2 => n13602, B1 => n684, B2 => 
                           n13599, C1 => n14625, C2 => n13596, ZN => n11363);
   U2583 : OAI222_X1 port map( A1 => n14877, A2 => n13602, B1 => n683, B2 => 
                           n13599, C1 => n14619, C2 => n13596, ZN => n11362);
   U2584 : OAI222_X1 port map( A1 => n14871, A2 => n13602, B1 => n682, B2 => 
                           n13599, C1 => n14613, C2 => n13596, ZN => n11361);
   U2585 : OAI222_X1 port map( A1 => n14865, A2 => n13602, B1 => n681, B2 => 
                           n13599, C1 => n14607, C2 => n13596, ZN => n11360);
   U2586 : OAI222_X1 port map( A1 => n14859, A2 => n13602, B1 => n680, B2 => 
                           n13599, C1 => n14601, C2 => n13596, ZN => n11359);
   U2587 : OAI222_X1 port map( A1 => n14853, A2 => n13602, B1 => n679, B2 => 
                           n13599, C1 => n14595, C2 => n13596, ZN => n11358);
   U2588 : OAI222_X1 port map( A1 => n14847, A2 => n13602, B1 => n678, B2 => 
                           n13599, C1 => n14589, C2 => n13596, ZN => n11357);
   U2589 : OAI222_X1 port map( A1 => n14841, A2 => n13602, B1 => n677, B2 => 
                           n13599, C1 => n14583, C2 => n13596, ZN => n11356);
   U2590 : OAI222_X1 port map( A1 => n14835, A2 => n13602, B1 => n676, B2 => 
                           n13599, C1 => n14577, C2 => n13596, ZN => n11355);
   U2591 : OAI222_X1 port map( A1 => n14829, A2 => n13602, B1 => n675, B2 => 
                           n13599, C1 => n14571, C2 => n13596, ZN => n11354);
   U2592 : OAI222_X1 port map( A1 => n14823, A2 => n13602, B1 => n674, B2 => 
                           n13599, C1 => n14565, C2 => n13596, ZN => n11353);
   U2593 : OAI222_X1 port map( A1 => n14817, A2 => n13601, B1 => n673, B2 => 
                           n13598, C1 => n14559, C2 => n13596, ZN => n11352);
   U2594 : OAI222_X1 port map( A1 => n14811, A2 => n13601, B1 => n672, B2 => 
                           n13598, C1 => n14553, C2 => n13595, ZN => n11351);
   U2595 : OAI222_X1 port map( A1 => n14805, A2 => n13601, B1 => n671, B2 => 
                           n13598, C1 => n14547, C2 => n13595, ZN => n11350);
   U2596 : OAI222_X1 port map( A1 => n14799, A2 => n13601, B1 => n670, B2 => 
                           n13598, C1 => n14541, C2 => n13595, ZN => n11349);
   U2597 : OAI222_X1 port map( A1 => n14793, A2 => n13601, B1 => n669, B2 => 
                           n13598, C1 => n14535, C2 => n13595, ZN => n11348);
   U2598 : OAI222_X1 port map( A1 => n14787, A2 => n13601, B1 => n668, B2 => 
                           n13598, C1 => n14529, C2 => n13595, ZN => n11347);
   U2599 : OAI222_X1 port map( A1 => n14781, A2 => n13601, B1 => n667, B2 => 
                           n13598, C1 => n14523, C2 => n13595, ZN => n11346);
   U2600 : OAI222_X1 port map( A1 => n14775, A2 => n13601, B1 => n666, B2 => 
                           n13598, C1 => n14517, C2 => n13595, ZN => n11345);
   U2601 : OAI222_X1 port map( A1 => n14769, A2 => n13601, B1 => n665, B2 => 
                           n13598, C1 => n14511, C2 => n13595, ZN => n11344);
   U2602 : OAI222_X1 port map( A1 => n14763, A2 => n13601, B1 => n664, B2 => 
                           n13598, C1 => n14712, C2 => n13595, ZN => n11343);
   U2603 : OAI222_X1 port map( A1 => n14757, A2 => n13601, B1 => n663, B2 => 
                           n13598, C1 => n14700, C2 => n13595, ZN => n11342);
   U2604 : OAI222_X1 port map( A1 => n14751, A2 => n13601, B1 => n662, B2 => 
                           n13598, C1 => n14695, C2 => n13595, ZN => n11341);
   U2605 : OAI222_X1 port map( A1 => n14883, A2 => n13611, B1 => n660, B2 => 
                           n13608, C1 => n14625, C2 => n13605, ZN => n11395);
   U2606 : OAI222_X1 port map( A1 => n14877, A2 => n13611, B1 => n659, B2 => 
                           n13608, C1 => n14619, C2 => n13605, ZN => n11394);
   U2607 : OAI222_X1 port map( A1 => n14871, A2 => n13611, B1 => n658, B2 => 
                           n13608, C1 => n14613, C2 => n13605, ZN => n11393);
   U2608 : OAI222_X1 port map( A1 => n14865, A2 => n13611, B1 => n657, B2 => 
                           n13608, C1 => n14607, C2 => n13605, ZN => n11392);
   U2609 : OAI222_X1 port map( A1 => n14859, A2 => n13611, B1 => n656, B2 => 
                           n13608, C1 => n14601, C2 => n13605, ZN => n11391);
   U2610 : OAI222_X1 port map( A1 => n14853, A2 => n13611, B1 => n655, B2 => 
                           n13608, C1 => n14595, C2 => n13605, ZN => n11390);
   U2611 : OAI222_X1 port map( A1 => n14847, A2 => n13611, B1 => n654, B2 => 
                           n13608, C1 => n14589, C2 => n13605, ZN => n11389);
   U2612 : OAI222_X1 port map( A1 => n14841, A2 => n13611, B1 => n653, B2 => 
                           n13608, C1 => n14583, C2 => n13605, ZN => n11388);
   U2613 : OAI222_X1 port map( A1 => n14835, A2 => n13611, B1 => n652, B2 => 
                           n13608, C1 => n14577, C2 => n13605, ZN => n11387);
   U2614 : OAI222_X1 port map( A1 => n14829, A2 => n13611, B1 => n651, B2 => 
                           n13608, C1 => n14571, C2 => n13605, ZN => n11386);
   U2615 : OAI222_X1 port map( A1 => n14823, A2 => n13611, B1 => n650, B2 => 
                           n13608, C1 => n14565, C2 => n13605, ZN => n11385);
   U2616 : OAI222_X1 port map( A1 => n14817, A2 => n13610, B1 => n649, B2 => 
                           n13607, C1 => n14559, C2 => n13605, ZN => n11384);
   U2617 : OAI222_X1 port map( A1 => n14811, A2 => n13610, B1 => n648, B2 => 
                           n13607, C1 => n14553, C2 => n13604, ZN => n11383);
   U2618 : OAI222_X1 port map( A1 => n14805, A2 => n13610, B1 => n647, B2 => 
                           n13607, C1 => n14547, C2 => n13604, ZN => n11382);
   U2619 : OAI222_X1 port map( A1 => n14799, A2 => n13610, B1 => n646, B2 => 
                           n13607, C1 => n14541, C2 => n13604, ZN => n11381);
   U2620 : OAI222_X1 port map( A1 => n14793, A2 => n13610, B1 => n645, B2 => 
                           n13607, C1 => n14535, C2 => n13604, ZN => n11380);
   U2621 : OAI222_X1 port map( A1 => n14787, A2 => n13610, B1 => n644, B2 => 
                           n13607, C1 => n14529, C2 => n13604, ZN => n11379);
   U2622 : OAI222_X1 port map( A1 => n14781, A2 => n13610, B1 => n643, B2 => 
                           n13607, C1 => n14523, C2 => n13604, ZN => n11378);
   U2623 : OAI222_X1 port map( A1 => n14775, A2 => n13610, B1 => n642, B2 => 
                           n13607, C1 => n14517, C2 => n13604, ZN => n11377);
   U2624 : OAI222_X1 port map( A1 => n14769, A2 => n13610, B1 => n641, B2 => 
                           n13607, C1 => n14511, C2 => n13604, ZN => n11376);
   U2625 : OAI222_X1 port map( A1 => n14763, A2 => n13610, B1 => n640, B2 => 
                           n13607, C1 => n14712, C2 => n13604, ZN => n11375);
   U2626 : OAI222_X1 port map( A1 => n14757, A2 => n13610, B1 => n639, B2 => 
                           n13607, C1 => n14700, C2 => n13604, ZN => n11374);
   U2627 : OAI222_X1 port map( A1 => n14751, A2 => n13610, B1 => n638, B2 => 
                           n13607, C1 => n14695, C2 => n13604, ZN => n11373);
   U2628 : OAI222_X1 port map( A1 => n14883, A2 => n13629, B1 => n636, B2 => 
                           n13626, C1 => n14625, C2 => n13623, ZN => n11459);
   U2629 : OAI222_X1 port map( A1 => n14877, A2 => n13629, B1 => n635, B2 => 
                           n13626, C1 => n14619, C2 => n13623, ZN => n11458);
   U2630 : OAI222_X1 port map( A1 => n14871, A2 => n13629, B1 => n634, B2 => 
                           n13626, C1 => n14613, C2 => n13623, ZN => n11457);
   U2631 : OAI222_X1 port map( A1 => n14865, A2 => n13629, B1 => n633, B2 => 
                           n13626, C1 => n14607, C2 => n13623, ZN => n11456);
   U2632 : OAI222_X1 port map( A1 => n14859, A2 => n13629, B1 => n632, B2 => 
                           n13626, C1 => n14601, C2 => n13623, ZN => n11455);
   U2633 : OAI222_X1 port map( A1 => n14853, A2 => n13629, B1 => n631, B2 => 
                           n13626, C1 => n14595, C2 => n13623, ZN => n11454);
   U2634 : OAI222_X1 port map( A1 => n14847, A2 => n13629, B1 => n630, B2 => 
                           n13626, C1 => n14589, C2 => n13623, ZN => n11453);
   U2635 : OAI222_X1 port map( A1 => n14841, A2 => n13629, B1 => n629, B2 => 
                           n13626, C1 => n14583, C2 => n13623, ZN => n11452);
   U2636 : OAI222_X1 port map( A1 => n14835, A2 => n13629, B1 => n628, B2 => 
                           n13626, C1 => n14577, C2 => n13623, ZN => n11451);
   U2637 : OAI222_X1 port map( A1 => n14883, A2 => n14294, B1 => n14290, B2 => 
                           n626, C1 => n14624, C2 => n14288, ZN => n9211);
   U2638 : OAI222_X1 port map( A1 => n14877, A2 => n14294, B1 => n14290, B2 => 
                           n625, C1 => n14618, C2 => n14288, ZN => n9209);
   U2639 : OAI222_X1 port map( A1 => n14871, A2 => n14294, B1 => n14290, B2 => 
                           n624, C1 => n14612, C2 => n14288, ZN => n9207);
   U2640 : OAI222_X1 port map( A1 => n14865, A2 => n14294, B1 => n14291, B2 => 
                           n623, C1 => n14606, C2 => n14288, ZN => n9205);
   U2641 : OAI222_X1 port map( A1 => n14859, A2 => n14294, B1 => n14291, B2 => 
                           n622, C1 => n14600, C2 => n14288, ZN => n9203);
   U2642 : OAI222_X1 port map( A1 => n14853, A2 => n14294, B1 => n14291, B2 => 
                           n621, C1 => n14594, C2 => n14288, ZN => n9201);
   U2643 : OAI222_X1 port map( A1 => n14847, A2 => n14294, B1 => n14291, B2 => 
                           n620, C1 => n14588, C2 => n14288, ZN => n9199);
   U2644 : OAI222_X1 port map( A1 => n14841, A2 => n14294, B1 => n14291, B2 => 
                           n619, C1 => n14582, C2 => n14288, ZN => n9197);
   U2645 : OAI222_X1 port map( A1 => n14835, A2 => n14294, B1 => n14291, B2 => 
                           n618, C1 => n14576, C2 => n14288, ZN => n9195);
   U2646 : OAI222_X1 port map( A1 => n14829, A2 => n14294, B1 => n14291, B2 => 
                           n617, C1 => n14570, C2 => n14288, ZN => n9193);
   U2647 : OAI222_X1 port map( A1 => n14817, A2 => n14293, B1 => n14291, B2 => 
                           n615, C1 => n14558, C2 => n14288, ZN => n9189);
   U2648 : OAI222_X1 port map( A1 => n14811, A2 => n14293, B1 => n14291, B2 => 
                           n614, C1 => n14552, C2 => n14287, ZN => n9187);
   U2649 : OAI222_X1 port map( A1 => n14805, A2 => n14293, B1 => n14291, B2 => 
                           n613, C1 => n14546, C2 => n14287, ZN => n9185);
   U2650 : OAI222_X1 port map( A1 => n14799, A2 => n14293, B1 => n14291, B2 => 
                           n612, C1 => n14540, C2 => n14287, ZN => n9183);
   U2651 : OAI222_X1 port map( A1 => n14793, A2 => n14293, B1 => n14292, B2 => 
                           n611, C1 => n14534, C2 => n14287, ZN => n9181);
   U2652 : OAI222_X1 port map( A1 => n14787, A2 => n14293, B1 => n14292, B2 => 
                           n610, C1 => n14528, C2 => n14287, ZN => n9179);
   U2653 : OAI222_X1 port map( A1 => n14781, A2 => n14293, B1 => n14292, B2 => 
                           n609, C1 => n14522, C2 => n14287, ZN => n9177);
   U2654 : OAI222_X1 port map( A1 => n14775, A2 => n14293, B1 => n14292, B2 => 
                           n608, C1 => n14516, C2 => n14287, ZN => n9175);
   U2655 : OAI222_X1 port map( A1 => n14769, A2 => n14293, B1 => n14292, B2 => 
                           n607, C1 => n14510, C2 => n14287, ZN => n9173);
   U2656 : OAI222_X1 port map( A1 => n14763, A2 => n14293, B1 => n14292, B2 => 
                           n606, C1 => n14711, C2 => n14287, ZN => n9171);
   U2657 : OAI222_X1 port map( A1 => n14757, A2 => n14293, B1 => n14292, B2 => 
                           n605, C1 => n14699, C2 => n14287, ZN => n9169);
   U2658 : OAI222_X1 port map( A1 => n14751, A2 => n14293, B1 => n14290, B2 => 
                           n604, C1 => n14695, C2 => n14287, ZN => n9167);
   U2659 : OAI222_X1 port map( A1 => n14883, A2 => n14305, B1 => n14301, B2 => 
                           n602, C1 => n14624, C2 => n14299, ZN => n9251);
   U2660 : OAI222_X1 port map( A1 => n14877, A2 => n14305, B1 => n14301, B2 => 
                           n601, C1 => n14618, C2 => n14299, ZN => n9250);
   U2661 : OAI222_X1 port map( A1 => n14871, A2 => n14305, B1 => n14301, B2 => 
                           n600, C1 => n14612, C2 => n14299, ZN => n9249);
   U2662 : OAI222_X1 port map( A1 => n14865, A2 => n14305, B1 => n14302, B2 => 
                           n599, C1 => n14606, C2 => n14299, ZN => n9248);
   U2663 : OAI222_X1 port map( A1 => n14859, A2 => n14305, B1 => n14302, B2 => 
                           n598, C1 => n14600, C2 => n14299, ZN => n9247);
   U2664 : OAI222_X1 port map( A1 => n14853, A2 => n14305, B1 => n14302, B2 => 
                           n597, C1 => n14594, C2 => n14299, ZN => n9246);
   U2665 : OAI222_X1 port map( A1 => n14847, A2 => n14305, B1 => n14302, B2 => 
                           n596, C1 => n14588, C2 => n14299, ZN => n9245);
   U2666 : OAI222_X1 port map( A1 => n14841, A2 => n14305, B1 => n14302, B2 => 
                           n595, C1 => n14582, C2 => n14299, ZN => n9244);
   U2667 : OAI222_X1 port map( A1 => n14835, A2 => n14305, B1 => n14302, B2 => 
                           n594, C1 => n14576, C2 => n14299, ZN => n9243);
   U2668 : OAI222_X1 port map( A1 => n14829, A2 => n14305, B1 => n14302, B2 => 
                           n593, C1 => n14570, C2 => n14299, ZN => n9242);
   U2669 : OAI222_X1 port map( A1 => n14817, A2 => n14304, B1 => n14302, B2 => 
                           n591, C1 => n14558, C2 => n14299, ZN => n9240);
   U2670 : OAI222_X1 port map( A1 => n14811, A2 => n14304, B1 => n14302, B2 => 
                           n590, C1 => n14552, C2 => n14298, ZN => n9239);
   U2671 : OAI222_X1 port map( A1 => n14805, A2 => n14304, B1 => n14302, B2 => 
                           n589, C1 => n14546, C2 => n14298, ZN => n9238);
   U2672 : OAI222_X1 port map( A1 => n14799, A2 => n14304, B1 => n14302, B2 => 
                           n588, C1 => n14540, C2 => n14298, ZN => n9237);
   U2673 : OAI222_X1 port map( A1 => n14793, A2 => n14304, B1 => n14303, B2 => 
                           n587, C1 => n14534, C2 => n14298, ZN => n9236);
   U2674 : OAI222_X1 port map( A1 => n14787, A2 => n14304, B1 => n14303, B2 => 
                           n586, C1 => n14528, C2 => n14298, ZN => n9235);
   U2675 : OAI222_X1 port map( A1 => n14781, A2 => n14304, B1 => n14303, B2 => 
                           n585, C1 => n14522, C2 => n14298, ZN => n9234);
   U2676 : OAI222_X1 port map( A1 => n14775, A2 => n14304, B1 => n14303, B2 => 
                           n584, C1 => n14516, C2 => n14298, ZN => n9233);
   U2677 : OAI222_X1 port map( A1 => n14769, A2 => n14304, B1 => n14303, B2 => 
                           n583, C1 => n14510, C2 => n14298, ZN => n9232);
   U2678 : OAI222_X1 port map( A1 => n14763, A2 => n14304, B1 => n14303, B2 => 
                           n582, C1 => n14711, C2 => n14298, ZN => n9231);
   U2679 : OAI222_X1 port map( A1 => n14757, A2 => n14304, B1 => n14303, B2 => 
                           n581, C1 => n14699, C2 => n14298, ZN => n9230);
   U2680 : OAI222_X1 port map( A1 => n14751, A2 => n14304, B1 => n14301, B2 => 
                           n580, C1 => n14695, C2 => n14298, ZN => n9229);
   U2681 : OAI222_X1 port map( A1 => n14882, A2 => n14325, B1 => n14322, B2 => 
                           n578, C1 => n14624, C2 => n14319, ZN => n9315);
   U2682 : OAI222_X1 port map( A1 => n14876, A2 => n14325, B1 => n14322, B2 => 
                           n577, C1 => n14618, C2 => n14319, ZN => n9314);
   U2683 : OAI222_X1 port map( A1 => n14870, A2 => n14325, B1 => n14322, B2 => 
                           n576, C1 => n14612, C2 => n14319, ZN => n9313);
   U2684 : OAI222_X1 port map( A1 => n14864, A2 => n14325, B1 => n14322, B2 => 
                           n575, C1 => n14606, C2 => n14319, ZN => n9312);
   U2685 : OAI222_X1 port map( A1 => n14858, A2 => n14325, B1 => n14322, B2 => 
                           n574, C1 => n14600, C2 => n14319, ZN => n9311);
   U2686 : OAI222_X1 port map( A1 => n14852, A2 => n14325, B1 => n14322, B2 => 
                           n573, C1 => n14594, C2 => n14319, ZN => n9310);
   U2687 : OAI222_X1 port map( A1 => n14846, A2 => n14325, B1 => n14322, B2 => 
                           n572, C1 => n14588, C2 => n14319, ZN => n9309);
   U2688 : OAI222_X1 port map( A1 => n14840, A2 => n14325, B1 => n14322, B2 => 
                           n571, C1 => n14582, C2 => n14319, ZN => n9308);
   U2689 : OAI222_X1 port map( A1 => n14834, A2 => n14325, B1 => n14322, B2 => 
                           n570, C1 => n14576, C2 => n14319, ZN => n9307);
   U2690 : OAI222_X1 port map( A1 => n14828, A2 => n14325, B1 => n14322, B2 => 
                           n569, C1 => n14570, C2 => n14319, ZN => n9306);
   U2691 : OAI222_X1 port map( A1 => n14822, A2 => n14325, B1 => n14322, B2 => 
                           n568, C1 => n14564, C2 => n14319, ZN => n9305);
   U2692 : OAI222_X1 port map( A1 => n14816, A2 => n14324, B1 => n14321, B2 => 
                           n567, C1 => n14558, C2 => n14319, ZN => n9304);
   U2693 : OAI222_X1 port map( A1 => n14810, A2 => n14324, B1 => n14321, B2 => 
                           n566, C1 => n14552, C2 => n14318, ZN => n9303);
   U2694 : OAI222_X1 port map( A1 => n14804, A2 => n14324, B1 => n14321, B2 => 
                           n565, C1 => n14546, C2 => n14318, ZN => n9302);
   U2695 : OAI222_X1 port map( A1 => n14798, A2 => n14324, B1 => n14321, B2 => 
                           n564, C1 => n14540, C2 => n14318, ZN => n9301);
   U2696 : OAI222_X1 port map( A1 => n14792, A2 => n14324, B1 => n14321, B2 => 
                           n563, C1 => n14534, C2 => n14318, ZN => n9300);
   U2697 : OAI222_X1 port map( A1 => n14786, A2 => n14324, B1 => n14321, B2 => 
                           n562, C1 => n14528, C2 => n14318, ZN => n9299);
   U2698 : OAI222_X1 port map( A1 => n14780, A2 => n14324, B1 => n14321, B2 => 
                           n561, C1 => n14522, C2 => n14318, ZN => n9298);
   U2699 : OAI222_X1 port map( A1 => n14774, A2 => n14324, B1 => n14321, B2 => 
                           n560, C1 => n14516, C2 => n14318, ZN => n9297);
   U2700 : OAI222_X1 port map( A1 => n14768, A2 => n14324, B1 => n14321, B2 => 
                           n559, C1 => n14510, C2 => n14318, ZN => n9296);
   U2701 : OAI222_X1 port map( A1 => n14763, A2 => n14324, B1 => n14321, B2 => 
                           n558, C1 => n14711, C2 => n14318, ZN => n9295);
   U2702 : OAI222_X1 port map( A1 => n14757, A2 => n14324, B1 => n14321, B2 => 
                           n557, C1 => n14699, C2 => n14318, ZN => n9294);
   U2703 : OAI222_X1 port map( A1 => n14750, A2 => n14324, B1 => n14321, B2 => 
                           n556, C1 => n14696, C2 => n14318, ZN => n9293);
   U2704 : OAI222_X1 port map( A1 => n14882, A2 => n14363, B1 => n14360, B2 => 
                           n530, C1 => n14624, C2 => n14357, ZN => n9443);
   U2705 : OAI222_X1 port map( A1 => n14876, A2 => n14363, B1 => n14360, B2 => 
                           n529, C1 => n14618, C2 => n14357, ZN => n9442);
   U2706 : OAI222_X1 port map( A1 => n14870, A2 => n14363, B1 => n14360, B2 => 
                           n528, C1 => n14612, C2 => n14357, ZN => n9441);
   U2707 : OAI222_X1 port map( A1 => n14864, A2 => n14363, B1 => n14360, B2 => 
                           n527, C1 => n14606, C2 => n14357, ZN => n9440);
   U2708 : OAI222_X1 port map( A1 => n14858, A2 => n14363, B1 => n14360, B2 => 
                           n526, C1 => n14600, C2 => n14357, ZN => n9439);
   U2709 : OAI222_X1 port map( A1 => n14852, A2 => n14363, B1 => n14360, B2 => 
                           n525, C1 => n14594, C2 => n14357, ZN => n9438);
   U2710 : OAI222_X1 port map( A1 => n14846, A2 => n14363, B1 => n14360, B2 => 
                           n524, C1 => n14588, C2 => n14357, ZN => n9437);
   U2711 : OAI222_X1 port map( A1 => n14840, A2 => n14363, B1 => n14360, B2 => 
                           n523, C1 => n14582, C2 => n14357, ZN => n9436);
   U2712 : OAI222_X1 port map( A1 => n14834, A2 => n14363, B1 => n14360, B2 => 
                           n522, C1 => n14576, C2 => n14357, ZN => n9435);
   U2713 : OAI222_X1 port map( A1 => n14828, A2 => n14363, B1 => n14360, B2 => 
                           n521, C1 => n14570, C2 => n14357, ZN => n9434);
   U2714 : OAI222_X1 port map( A1 => n14822, A2 => n14363, B1 => n14360, B2 => 
                           n520, C1 => n14564, C2 => n14357, ZN => n9433);
   U2715 : OAI222_X1 port map( A1 => n14816, A2 => n14362, B1 => n14359, B2 => 
                           n519, C1 => n14558, C2 => n14357, ZN => n9432);
   U2716 : OAI222_X1 port map( A1 => n14810, A2 => n14362, B1 => n14359, B2 => 
                           n518, C1 => n14552, C2 => n14356, ZN => n9431);
   U2717 : OAI222_X1 port map( A1 => n14804, A2 => n14362, B1 => n14359, B2 => 
                           n517, C1 => n14546, C2 => n14356, ZN => n9430);
   U2718 : OAI222_X1 port map( A1 => n14798, A2 => n14362, B1 => n14359, B2 => 
                           n516, C1 => n14540, C2 => n14356, ZN => n9429);
   U2719 : OAI222_X1 port map( A1 => n14792, A2 => n14362, B1 => n14359, B2 => 
                           n515, C1 => n14534, C2 => n14356, ZN => n9428);
   U2720 : OAI222_X1 port map( A1 => n14786, A2 => n14362, B1 => n14359, B2 => 
                           n514, C1 => n14528, C2 => n14356, ZN => n9427);
   U2721 : OAI222_X1 port map( A1 => n14780, A2 => n14362, B1 => n14359, B2 => 
                           n513, C1 => n14522, C2 => n14356, ZN => n9426);
   U2722 : OAI222_X1 port map( A1 => n14774, A2 => n14362, B1 => n14359, B2 => 
                           n512, C1 => n14516, C2 => n14356, ZN => n9425);
   U2723 : OAI222_X1 port map( A1 => n14768, A2 => n14362, B1 => n14359, B2 => 
                           n511, C1 => n14510, C2 => n14356, ZN => n9424);
   U2724 : OAI222_X1 port map( A1 => n14764, A2 => n14362, B1 => n14359, B2 => 
                           n510, C1 => n14712, C2 => n14356, ZN => n9423);
   U2725 : OAI222_X1 port map( A1 => n14758, A2 => n14362, B1 => n14359, B2 => 
                           n509, C1 => n14700, C2 => n14356, ZN => n9422);
   U2726 : OAI222_X1 port map( A1 => n14752, A2 => n14362, B1 => n14359, B2 => 
                           n508, C1 => n14696, C2 => n14356, ZN => n9421);
   U2727 : OAI222_X1 port map( A1 => n14882, A2 => n14390, B1 => n14386, B2 => 
                           n506, C1 => n14624, C2 => n14384, ZN => n9539);
   U2728 : OAI222_X1 port map( A1 => n14876, A2 => n14390, B1 => n14386, B2 => 
                           n505, C1 => n14618, C2 => n14384, ZN => n9538);
   U2729 : OAI222_X1 port map( A1 => n14870, A2 => n14390, B1 => n14386, B2 => 
                           n504, C1 => n14612, C2 => n14384, ZN => n9537);
   U2730 : OAI222_X1 port map( A1 => n14864, A2 => n14390, B1 => n14387, B2 => 
                           n503, C1 => n14606, C2 => n14384, ZN => n9536);
   U2731 : OAI222_X1 port map( A1 => n14858, A2 => n14390, B1 => n14387, B2 => 
                           n502, C1 => n14600, C2 => n14384, ZN => n9535);
   U2732 : OAI222_X1 port map( A1 => n14852, A2 => n14390, B1 => n14387, B2 => 
                           n501, C1 => n14594, C2 => n14384, ZN => n9534);
   U2733 : OAI222_X1 port map( A1 => n14846, A2 => n14390, B1 => n14387, B2 => 
                           n500, C1 => n14588, C2 => n14384, ZN => n9533);
   U2734 : OAI222_X1 port map( A1 => n14840, A2 => n14390, B1 => n14387, B2 => 
                           n499, C1 => n14582, C2 => n14384, ZN => n9532);
   U2735 : OAI222_X1 port map( A1 => n14834, A2 => n14390, B1 => n14387, B2 => 
                           n498, C1 => n14576, C2 => n14384, ZN => n9531);
   U2736 : OAI222_X1 port map( A1 => n14828, A2 => n14390, B1 => n14387, B2 => 
                           n497, C1 => n14570, C2 => n14384, ZN => n9530);
   U2737 : OAI222_X1 port map( A1 => n14816, A2 => n14389, B1 => n14387, B2 => 
                           n495, C1 => n14558, C2 => n14384, ZN => n9528);
   U2738 : OAI222_X1 port map( A1 => n14810, A2 => n14389, B1 => n14387, B2 => 
                           n494, C1 => n14552, C2 => n14383, ZN => n9527);
   U2739 : OAI222_X1 port map( A1 => n14804, A2 => n14389, B1 => n14387, B2 => 
                           n493, C1 => n14546, C2 => n14383, ZN => n9526);
   U2740 : OAI222_X1 port map( A1 => n14798, A2 => n14389, B1 => n14387, B2 => 
                           n492, C1 => n14540, C2 => n14383, ZN => n9525);
   U2741 : OAI222_X1 port map( A1 => n14792, A2 => n14389, B1 => n14388, B2 => 
                           n491, C1 => n14534, C2 => n14383, ZN => n9524);
   U2742 : OAI222_X1 port map( A1 => n14786, A2 => n14389, B1 => n14388, B2 => 
                           n490, C1 => n14528, C2 => n14383, ZN => n9523);
   U2743 : OAI222_X1 port map( A1 => n14780, A2 => n14389, B1 => n14388, B2 => 
                           n489, C1 => n14522, C2 => n14383, ZN => n9522);
   U2744 : OAI222_X1 port map( A1 => n14774, A2 => n14389, B1 => n14388, B2 => 
                           n488, C1 => n14516, C2 => n14383, ZN => n9521);
   U2745 : OAI222_X1 port map( A1 => n14768, A2 => n14389, B1 => n14388, B2 => 
                           n487, C1 => n14510, C2 => n14383, ZN => n9520);
   U2746 : OAI222_X1 port map( A1 => n14762, A2 => n14389, B1 => n14388, B2 => 
                           n486, C1 => n14711, C2 => n14383, ZN => n9519);
   U2747 : OAI222_X1 port map( A1 => n14756, A2 => n14389, B1 => n14388, B2 => 
                           n485, C1 => n14699, C2 => n14383, ZN => n9518);
   U2748 : OAI222_X1 port map( A1 => n14750, A2 => n14389, B1 => n14386, B2 => 
                           n484, C1 => n14696, C2 => n14383, ZN => n9517);
   U2749 : OAI222_X1 port map( A1 => n14882, A2 => n14408, B1 => n14405, B2 => 
                           n482, C1 => n14623, C2 => n14402, ZN => n9603);
   U2750 : OAI222_X1 port map( A1 => n14876, A2 => n14408, B1 => n14405, B2 => 
                           n481, C1 => n14617, C2 => n14402, ZN => n9602);
   U2751 : OAI222_X1 port map( A1 => n14870, A2 => n14408, B1 => n14405, B2 => 
                           n480, C1 => n14611, C2 => n14402, ZN => n9601);
   U2752 : OAI222_X1 port map( A1 => n14864, A2 => n14408, B1 => n14405, B2 => 
                           n479, C1 => n14605, C2 => n14402, ZN => n9600);
   U2753 : OAI222_X1 port map( A1 => n14858, A2 => n14408, B1 => n14405, B2 => 
                           n478, C1 => n14599, C2 => n14402, ZN => n9599);
   U2754 : OAI222_X1 port map( A1 => n14852, A2 => n14408, B1 => n14405, B2 => 
                           n477, C1 => n14593, C2 => n14402, ZN => n9598);
   U2755 : OAI222_X1 port map( A1 => n14846, A2 => n14408, B1 => n14405, B2 => 
                           n476, C1 => n14587, C2 => n14402, ZN => n9597);
   U2756 : OAI222_X1 port map( A1 => n14840, A2 => n14408, B1 => n14405, B2 => 
                           n475, C1 => n14581, C2 => n14402, ZN => n9596);
   U2757 : OAI222_X1 port map( A1 => n14834, A2 => n14408, B1 => n14405, B2 => 
                           n474, C1 => n14575, C2 => n14402, ZN => n9595);
   U2758 : OAI222_X1 port map( A1 => n14828, A2 => n14408, B1 => n14405, B2 => 
                           n473, C1 => n14569, C2 => n14402, ZN => n9594);
   U2759 : OAI222_X1 port map( A1 => n14822, A2 => n14408, B1 => n14405, B2 => 
                           n472, C1 => n14563, C2 => n14402, ZN => n9593);
   U2760 : OAI222_X1 port map( A1 => n14816, A2 => n14407, B1 => n14404, B2 => 
                           n471, C1 => n14557, C2 => n14402, ZN => n9592);
   U2761 : OAI222_X1 port map( A1 => n14810, A2 => n14407, B1 => n14404, B2 => 
                           n470, C1 => n14551, C2 => n14401, ZN => n9591);
   U2762 : OAI222_X1 port map( A1 => n14804, A2 => n14407, B1 => n14404, B2 => 
                           n469, C1 => n14545, C2 => n14401, ZN => n9590);
   U2763 : OAI222_X1 port map( A1 => n14798, A2 => n14407, B1 => n14404, B2 => 
                           n468, C1 => n14539, C2 => n14401, ZN => n9589);
   U2764 : OAI222_X1 port map( A1 => n14792, A2 => n14407, B1 => n14404, B2 => 
                           n467, C1 => n14533, C2 => n14401, ZN => n9588);
   U2765 : OAI222_X1 port map( A1 => n14786, A2 => n14407, B1 => n14404, B2 => 
                           n466, C1 => n14527, C2 => n14401, ZN => n9587);
   U2766 : OAI222_X1 port map( A1 => n14780, A2 => n14407, B1 => n14404, B2 => 
                           n465, C1 => n14521, C2 => n14401, ZN => n9586);
   U2767 : OAI222_X1 port map( A1 => n14774, A2 => n14407, B1 => n14404, B2 => 
                           n464, C1 => n14515, C2 => n14401, ZN => n9585);
   U2768 : OAI222_X1 port map( A1 => n14768, A2 => n14407, B1 => n14404, B2 => 
                           n463, C1 => n14509, C2 => n14401, ZN => n9584);
   U2769 : OAI222_X1 port map( A1 => n14762, A2 => n14407, B1 => n14404, B2 => 
                           n462, C1 => n14711, C2 => n14401, ZN => n9583);
   U2770 : OAI222_X1 port map( A1 => n14756, A2 => n14407, B1 => n14404, B2 => 
                           n461, C1 => n14699, C2 => n14401, ZN => n9582);
   U2771 : OAI222_X1 port map( A1 => n14750, A2 => n14407, B1 => n14404, B2 => 
                           n460, C1 => n14696, C2 => n14401, ZN => n9581);
   U2772 : AOI221_X1 port map( B1 => n14737, B2 => n1775, C1 => n14740, C2 => 
                           n1768, A => n4279, ZN => n4272);
   U2773 : OAI22_X1 port map( A1 => n214, A2 => n4093, B1 => n222, B2 => n13868
                           , ZN => n4279);
   U2774 : AOI221_X1 port map( B1 => n14738, B2 => n2337, C1 => n14741, C2 => 
                           n2313, A => n4834, ZN => n4827);
   U2775 : OAI22_X1 port map( A1 => n1522, A2 => n4093, B1 => n1546, B2 => 
                           n13868, ZN => n4834);
   U2776 : AOI221_X1 port map( B1 => n14738, B2 => n2336, C1 => n14741, C2 => 
                           n2312, A => n4871, ZN => n4864);
   U2777 : OAI22_X1 port map( A1 => n1521, A2 => n4093, B1 => n1545, B2 => 
                           n13868, ZN => n4871);
   U2778 : AOI221_X1 port map( B1 => n14738, B2 => n2335, C1 => n14741, C2 => 
                           n2311, A => n4908, ZN => n4901);
   U2779 : OAI22_X1 port map( A1 => n1520, A2 => n4093, B1 => n1544, B2 => 
                           n13868, ZN => n4908);
   U2780 : AOI221_X1 port map( B1 => n14738, B2 => n2334, C1 => n14741, C2 => 
                           n2310, A => n4945, ZN => n4938);
   U2781 : OAI22_X1 port map( A1 => n1519, A2 => n4093, B1 => n1543, B2 => 
                           n13868, ZN => n4945);
   U2782 : AOI221_X1 port map( B1 => n14738, B2 => n2340, C1 => n14741, C2 => 
                           n2316, A => n4723, ZN => n4716);
   U2783 : OAI22_X1 port map( A1 => n1525, A2 => n13870, B1 => n1549, B2 => 
                           n13869, ZN => n4723);
   U2784 : AOI221_X1 port map( B1 => n14738, B2 => n2339, C1 => n14741, C2 => 
                           n2315, A => n4760, ZN => n4753);
   U2785 : OAI22_X1 port map( A1 => n1524, A2 => n4093, B1 => n1548, B2 => 
                           n13868, ZN => n4760);
   U2786 : AOI221_X1 port map( B1 => n14739, B2 => n2333, C1 => n14742, C2 => 
                           n2309, A => n4982, ZN => n4975);
   U2787 : OAI22_X1 port map( A1 => n1518, A2 => n13870, B1 => n1542, B2 => 
                           n13868, ZN => n4982);
   U2788 : AOI221_X1 port map( B1 => n14739, B2 => n2332, C1 => n14742, C2 => 
                           n2308, A => n5019, ZN => n5012);
   U2789 : OAI22_X1 port map( A1 => n1517, A2 => n4093, B1 => n1541, B2 => 
                           n13868, ZN => n5019);
   U2790 : AOI221_X1 port map( B1 => n14739, B2 => n2331, C1 => n14742, C2 => 
                           n2307, A => n5056, ZN => n5049);
   U2791 : OAI22_X1 port map( A1 => n1516, A2 => n13870, B1 => n1540, B2 => 
                           n13868, ZN => n5056);
   U2792 : AOI221_X1 port map( B1 => n14739, B2 => n2330, C1 => n14742, C2 => 
                           n2306, A => n5093, ZN => n5086);
   U2793 : OAI22_X1 port map( A1 => n1515, A2 => n4093, B1 => n1539, B2 => 
                           n13868, ZN => n5093);
   U2794 : AOI221_X1 port map( B1 => n14739, B2 => n2329, C1 => n14742, C2 => 
                           n2305, A => n5130, ZN => n5123);
   U2795 : OAI22_X1 port map( A1 => n1514, A2 => n13870, B1 => n1538, B2 => 
                           n13868, ZN => n5130);
   U2796 : AOI221_X1 port map( B1 => n14739, B2 => n2328, C1 => n14742, C2 => 
                           n2304, A => n5167, ZN => n5160);
   U2797 : OAI22_X1 port map( A1 => n1513, A2 => n4093, B1 => n1537, B2 => 
                           n13868, ZN => n5167);
   U2798 : AOI221_X1 port map( B1 => n14737, B2 => n1780, C1 => n14740, C2 => 
                           n1773, A => n4092, ZN => n4085);
   U2799 : OAI22_X1 port map( A1 => n219, A2 => n4093, B1 => n227, B2 => n13869
                           , ZN => n4092);
   U2800 : AOI221_X1 port map( B1 => n14737, B2 => n1779, C1 => n14740, C2 => 
                           n1772, A => n4131, ZN => n4124);
   U2801 : OAI22_X1 port map( A1 => n218, A2 => n4093, B1 => n226, B2 => n13868
                           , ZN => n4131);
   U2802 : AOI221_X1 port map( B1 => n14737, B2 => n1778, C1 => n14740, C2 => 
                           n1771, A => n4168, ZN => n4161);
   U2803 : OAI22_X1 port map( A1 => n217, A2 => n4093, B1 => n225, B2 => n13869
                           , ZN => n4168);
   U2804 : AOI221_X1 port map( B1 => n14737, B2 => n1777, C1 => n14740, C2 => 
                           n1770, A => n4205, ZN => n4198);
   U2805 : OAI22_X1 port map( A1 => n216, A2 => n4093, B1 => n224, B2 => n13868
                           , ZN => n4205);
   U2806 : AOI221_X1 port map( B1 => n14737, B2 => n1776, C1 => n14740, C2 => 
                           n1769, A => n4242, ZN => n4235);
   U2807 : OAI22_X1 port map( A1 => n215, A2 => n4093, B1 => n223, B2 => n13869
                           , ZN => n4242);
   U2808 : AOI221_X1 port map( B1 => n14737, B2 => n1774, C1 => n14740, C2 => 
                           n1767, A => n4316, ZN => n4309);
   U2809 : OAI22_X1 port map( A1 => n213, A2 => n13870, B1 => n221, B2 => 
                           n13869, ZN => n4316);
   U2810 : AOI221_X1 port map( B1 => n14737, B2 => n2350, C1 => n14740, C2 => 
                           n2326, A => n4353, ZN => n4346);
   U2811 : OAI22_X1 port map( A1 => n1535, A2 => n13870, B1 => n1559, B2 => 
                           n13869, ZN => n4353);
   U2812 : AOI221_X1 port map( B1 => n14737, B2 => n2349, C1 => n14740, C2 => 
                           n2325, A => n4390, ZN => n4383);
   U2813 : OAI22_X1 port map( A1 => n1534, A2 => n13870, B1 => n1558, B2 => 
                           n13869, ZN => n4390);
   U2814 : AOI221_X1 port map( B1 => n14737, B2 => n2348, C1 => n14740, C2 => 
                           n2324, A => n4427, ZN => n4420);
   U2815 : OAI22_X1 port map( A1 => n1533, A2 => n13870, B1 => n1557, B2 => 
                           n13869, ZN => n4427);
   U2816 : AOI221_X1 port map( B1 => n14737, B2 => n2347, C1 => n14740, C2 => 
                           n2323, A => n4464, ZN => n4457);
   U2817 : OAI22_X1 port map( A1 => n1532, A2 => n13870, B1 => n1556, B2 => 
                           n13869, ZN => n4464);
   U2818 : AOI221_X1 port map( B1 => n14737, B2 => n2346, C1 => n14740, C2 => 
                           n2322, A => n4501, ZN => n4494);
   U2819 : OAI22_X1 port map( A1 => n1531, A2 => n13870, B1 => n1555, B2 => 
                           n13869, ZN => n4501);
   U2820 : AOI221_X1 port map( B1 => n14738, B2 => n2345, C1 => n14741, C2 => 
                           n2321, A => n4538, ZN => n4531);
   U2821 : OAI22_X1 port map( A1 => n1530, A2 => n13870, B1 => n1554, B2 => 
                           n13869, ZN => n4538);
   U2822 : AOI221_X1 port map( B1 => n14738, B2 => n2344, C1 => n14741, C2 => 
                           n2320, A => n4575, ZN => n4568);
   U2823 : OAI22_X1 port map( A1 => n1529, A2 => n13870, B1 => n1553, B2 => 
                           n13869, ZN => n4575);
   U2824 : AOI221_X1 port map( B1 => n14738, B2 => n2343, C1 => n14741, C2 => 
                           n2319, A => n4612, ZN => n4605);
   U2825 : OAI22_X1 port map( A1 => n1528, A2 => n13870, B1 => n1552, B2 => 
                           n13869, ZN => n4612);
   U2826 : AOI221_X1 port map( B1 => n14738, B2 => n2342, C1 => n14741, C2 => 
                           n2318, A => n4649, ZN => n4642);
   U2827 : OAI22_X1 port map( A1 => n1527, A2 => n13870, B1 => n1551, B2 => 
                           n13869, ZN => n4649);
   U2828 : AOI221_X1 port map( B1 => n14738, B2 => n2341, C1 => n14741, C2 => 
                           n2317, A => n4686, ZN => n4679);
   U2829 : OAI22_X1 port map( A1 => n1526, A2 => n13870, B1 => n1550, B2 => 
                           n13869, ZN => n4686);
   U2830 : AOI221_X1 port map( B1 => n13705, B2 => n1780, C1 => n13702, C2 => 
                           n1773, A => n5415, ZN => n5408);
   U2831 : OAI22_X1 port map( A1 => n219, A2 => n13699, B1 => n227, B2 => 
                           n13696, ZN => n5415);
   U2832 : AOI221_X1 port map( B1 => n13705, B2 => n1778, C1 => n13702, C2 => 
                           n1771, A => n5489, ZN => n5482);
   U2833 : OAI22_X1 port map( A1 => n217, A2 => n13699, B1 => n225, B2 => 
                           n13696, ZN => n5489);
   U2834 : AOI221_X1 port map( B1 => n13705, B2 => n1777, C1 => n13702, C2 => 
                           n1770, A => n5526, ZN => n5519);
   U2835 : OAI22_X1 port map( A1 => n216, A2 => n13699, B1 => n224, B2 => 
                           n13696, ZN => n5526);
   U2836 : AOI221_X1 port map( B1 => n13705, B2 => n1776, C1 => n13702, C2 => 
                           n1769, A => n5563, ZN => n5556);
   U2837 : OAI22_X1 port map( A1 => n215, A2 => n13699, B1 => n223, B2 => 
                           n13696, ZN => n5563);
   U2838 : AOI221_X1 port map( B1 => n13705, B2 => n1775, C1 => n13702, C2 => 
                           n1768, A => n5600, ZN => n5593);
   U2839 : OAI22_X1 port map( A1 => n214, A2 => n13699, B1 => n222, B2 => 
                           n13696, ZN => n5600);
   U2840 : AOI221_X1 port map( B1 => n13703, B2 => n2337, C1 => n13700, C2 => 
                           n2313, A => n6155, ZN => n6148);
   U2841 : OAI22_X1 port map( A1 => n1522, A2 => n13697, B1 => n1546, B2 => 
                           n13694, ZN => n6155);
   U2842 : AOI221_X1 port map( B1 => n13703, B2 => n2336, C1 => n13700, C2 => 
                           n2312, A => n6192, ZN => n6185);
   U2843 : OAI22_X1 port map( A1 => n1521, A2 => n13697, B1 => n1545, B2 => 
                           n13694, ZN => n6192);
   U2844 : AOI221_X1 port map( B1 => n13703, B2 => n2335, C1 => n13700, C2 => 
                           n2311, A => n6229, ZN => n6222);
   U2845 : OAI22_X1 port map( A1 => n1520, A2 => n13697, B1 => n1544, B2 => 
                           n13694, ZN => n6229);
   U2846 : AOI221_X1 port map( B1 => n13703, B2 => n2334, C1 => n13700, C2 => 
                           n2310, A => n6266, ZN => n6259);
   U2847 : OAI22_X1 port map( A1 => n1519, A2 => n13697, B1 => n1543, B2 => 
                           n13694, ZN => n6266);
   U2848 : AOI221_X1 port map( B1 => n13703, B2 => n2333, C1 => n13700, C2 => 
                           n2309, A => n6303, ZN => n6296);
   U2849 : OAI22_X1 port map( A1 => n1518, A2 => n13697, B1 => n1542, B2 => 
                           n13694, ZN => n6303);
   U2850 : AOI221_X1 port map( B1 => n13703, B2 => n2332, C1 => n13700, C2 => 
                           n2308, A => n6340, ZN => n6333);
   U2851 : OAI22_X1 port map( A1 => n1517, A2 => n13697, B1 => n1541, B2 => 
                           n13694, ZN => n6340);
   U2852 : AOI221_X1 port map( B1 => n13703, B2 => n2331, C1 => n13700, C2 => 
                           n2307, A => n6377, ZN => n6370);
   U2853 : OAI22_X1 port map( A1 => n1516, A2 => n13697, B1 => n1540, B2 => 
                           n13694, ZN => n6377);
   U2854 : AOI221_X1 port map( B1 => n13703, B2 => n2330, C1 => n13700, C2 => 
                           n2306, A => n6414, ZN => n6407);
   U2855 : OAI22_X1 port map( A1 => n1515, A2 => n13697, B1 => n1539, B2 => 
                           n13694, ZN => n6414);
   U2856 : AOI221_X1 port map( B1 => n13703, B2 => n2329, C1 => n13700, C2 => 
                           n2305, A => n6451, ZN => n6444);
   U2857 : OAI22_X1 port map( A1 => n1514, A2 => n13697, B1 => n1538, B2 => 
                           n13694, ZN => n6451);
   U2858 : AOI221_X1 port map( B1 => n13703, B2 => n2328, C1 => n13700, C2 => 
                           n2304, A => n6488, ZN => n6481);
   U2859 : OAI22_X1 port map( A1 => n1513, A2 => n13697, B1 => n1537, B2 => 
                           n13694, ZN => n6488);
   U2860 : AOI221_X1 port map( B1 => n13704, B2 => n2340, C1 => n13701, C2 => 
                           n2316, A => n6044, ZN => n6037);
   U2861 : OAI22_X1 port map( A1 => n1525, A2 => n13698, B1 => n1549, B2 => 
                           n13695, ZN => n6044);
   U2862 : AOI221_X1 port map( B1 => n13704, B2 => n2339, C1 => n13701, C2 => 
                           n2315, A => n6081, ZN => n6074);
   U2863 : OAI22_X1 port map( A1 => n1524, A2 => n13698, B1 => n1548, B2 => 
                           n13695, ZN => n6081);
   U2864 : AOI221_X1 port map( B1 => n13705, B2 => n1779, C1 => n13702, C2 => 
                           n1772, A => n5452, ZN => n5445);
   U2865 : OAI22_X1 port map( A1 => n218, A2 => n13699, B1 => n226, B2 => 
                           n13696, ZN => n5452);
   U2866 : AOI221_X1 port map( B1 => n13705, B2 => n1774, C1 => n13702, C2 => 
                           n1767, A => n5637, ZN => n5630);
   U2867 : OAI22_X1 port map( A1 => n213, A2 => n13699, B1 => n221, B2 => 
                           n13696, ZN => n5637);
   U2868 : AOI221_X1 port map( B1 => n13704, B2 => n2350, C1 => n13701, C2 => 
                           n2326, A => n5674, ZN => n5667);
   U2869 : OAI22_X1 port map( A1 => n1535, A2 => n13698, B1 => n1559, B2 => 
                           n13695, ZN => n5674);
   U2870 : AOI221_X1 port map( B1 => n13704, B2 => n2349, C1 => n13701, C2 => 
                           n2325, A => n5711, ZN => n5704);
   U2871 : OAI22_X1 port map( A1 => n1534, A2 => n13698, B1 => n1558, B2 => 
                           n13695, ZN => n5711);
   U2872 : AOI221_X1 port map( B1 => n13704, B2 => n2348, C1 => n13701, C2 => 
                           n2324, A => n5748, ZN => n5741);
   U2873 : OAI22_X1 port map( A1 => n1533, A2 => n13698, B1 => n1557, B2 => 
                           n13695, ZN => n5748);
   U2874 : AOI221_X1 port map( B1 => n13704, B2 => n2347, C1 => n13701, C2 => 
                           n2323, A => n5785, ZN => n5778);
   U2875 : OAI22_X1 port map( A1 => n1532, A2 => n13698, B1 => n1556, B2 => 
                           n13695, ZN => n5785);
   U2876 : AOI221_X1 port map( B1 => n13704, B2 => n2346, C1 => n13701, C2 => 
                           n2322, A => n5822, ZN => n5815);
   U2877 : OAI22_X1 port map( A1 => n1531, A2 => n13698, B1 => n1555, B2 => 
                           n13695, ZN => n5822);
   U2878 : AOI221_X1 port map( B1 => n13704, B2 => n2345, C1 => n13701, C2 => 
                           n2321, A => n5859, ZN => n5852);
   U2879 : OAI22_X1 port map( A1 => n1530, A2 => n13698, B1 => n1554, B2 => 
                           n13695, ZN => n5859);
   U2880 : AOI221_X1 port map( B1 => n13704, B2 => n2344, C1 => n13701, C2 => 
                           n2320, A => n5896, ZN => n5889);
   U2881 : OAI22_X1 port map( A1 => n1529, A2 => n13698, B1 => n1553, B2 => 
                           n13695, ZN => n5896);
   U2882 : AOI221_X1 port map( B1 => n13704, B2 => n2343, C1 => n13701, C2 => 
                           n2319, A => n5933, ZN => n5926);
   U2883 : OAI22_X1 port map( A1 => n1528, A2 => n13698, B1 => n1552, B2 => 
                           n13695, ZN => n5933);
   U2884 : AOI221_X1 port map( B1 => n13704, B2 => n2342, C1 => n13701, C2 => 
                           n2318, A => n5970, ZN => n5963);
   U2885 : OAI22_X1 port map( A1 => n1527, A2 => n13698, B1 => n1551, B2 => 
                           n13695, ZN => n5970);
   U2886 : AOI221_X1 port map( B1 => n13704, B2 => n2341, C1 => n13701, C2 => 
                           n2317, A => n6007, ZN => n6000);
   U2887 : OAI22_X1 port map( A1 => n1526, A2 => n13698, B1 => n1550, B2 => 
                           n13695, ZN => n6007);
   U2888 : AOI221_X1 port map( B1 => n14098, B2 => n448, C1 => n14095, C2 => 
                           n424, A => n3545, ZN => n3538);
   U2889 : OAI22_X1 port map( A1 => n2483, A2 => n14092, B1 => n2481, B2 => 
                           n14089, ZN => n3545);
   U2890 : OAI22_X1 port map( A1 => n14000, A2 => n1607, B1 => n13997, B2 => 
                           n1062, ZN => n5207);
   U2891 : OAI22_X1 port map( A1 => n14000, A2 => n268, B1 => n13997, B2 => 
                           n260, ZN => n4000);
   U2892 : OAI22_X1 port map( A1 => n1623, A2 => n3312, B1 => n1644, B2 => 
                           n3313, ZN => n3311);
   U2893 : OAI22_X1 port map( A1 => n1622, A2 => n3312, B1 => n1643, B2 => 
                           n3313, ZN => n3350);
   U2894 : OAI22_X1 port map( A1 => n1621, A2 => n3312, B1 => n1642, B2 => 
                           n3313, ZN => n3387);
   U2895 : OAI22_X1 port map( A1 => n1620, A2 => n3312, B1 => n1641, B2 => 
                           n3313, ZN => n3424);
   U2896 : OAI22_X1 port map( A1 => n1616, A2 => n3312, B1 => n1637, B2 => 
                           n3313, ZN => n3572);
   U2897 : OAI22_X1 port map( A1 => n14224, A2 => n15, B1 => n14221, B2 => n23,
                           ZN => n2806);
   U2898 : OAI22_X1 port map( A1 => n14224, A2 => n14, B1 => n14221, B2 => n22,
                           ZN => n2890);
   U2899 : OAI22_X1 port map( A1 => n14224, A2 => n13, B1 => n14221, B2 => n21,
                           ZN => n2927);
   U2900 : OAI22_X1 port map( A1 => n14224, A2 => n12, B1 => n14221, B2 => n20,
                           ZN => n2964);
   U2901 : OAI22_X1 port map( A1 => n14224, A2 => n11, B1 => n14221, B2 => n19,
                           ZN => n3001);
   U2902 : OAI22_X1 port map( A1 => n14224, A2 => n10, B1 => n14221, B2 => n18,
                           ZN => n3038);
   U2903 : OAI22_X1 port map( A1 => n14224, A2 => n8, B1 => n14221, B2 => n17, 
                           ZN => n3075);
   U2904 : OAI22_X1 port map( A1 => n14224, A2 => n661, B1 => n14221, B2 => 
                           n685, ZN => n3112);
   U2905 : OAI22_X1 port map( A1 => n14251, A2 => n1730, B1 => n14248, B2 => 
                           n64, ZN => n2795);
   U2906 : OAI22_X1 port map( A1 => n14197, A2 => n1756, B1 => n14194, B2 => 
                           n195, ZN => n2821);
   U2907 : OAI22_X1 port map( A1 => n14251, A2 => n57, B1 => n14248, B2 => n63,
                           ZN => n2888);
   U2908 : OAI22_X1 port map( A1 => n14197, A2 => n188, B1 => n14194, B2 => 
                           n194, ZN => n2896);
   U2909 : OAI22_X1 port map( A1 => n14168, A2 => n132, B1 => n14167, B2 => 
                           n138, ZN => n2898);
   U2910 : OAI22_X1 port map( A1 => n14251, A2 => n1729, B1 => n14248, B2 => 
                           n62, ZN => n2925);
   U2911 : OAI22_X1 port map( A1 => n14197, A2 => n1755, B1 => n14194, B2 => 
                           n193, ZN => n2933);
   U2912 : OAI22_X1 port map( A1 => n14251, A2 => n1728, B1 => n14248, B2 => 
                           n61, ZN => n2962);
   U2913 : OAI22_X1 port map( A1 => n14197, A2 => n1754, B1 => n14194, B2 => 
                           n192, ZN => n2970);
   U2914 : OAI22_X1 port map( A1 => n14251, A2 => n1727, B1 => n14248, B2 => 
                           n60, ZN => n2999);
   U2915 : OAI22_X1 port map( A1 => n14197, A2 => n1753, B1 => n14194, B2 => 
                           n191, ZN => n3007);
   U2916 : OAI22_X1 port map( A1 => n14251, A2 => n1726, B1 => n14248, B2 => 
                           n59, ZN => n3036);
   U2917 : OAI22_X1 port map( A1 => n14197, A2 => n1752, B1 => n14194, B2 => 
                           n190, ZN => n3044);
   U2918 : OAI22_X1 port map( A1 => n14251, A2 => n1725, B1 => n14248, B2 => 
                           n58, ZN => n3073);
   U2919 : OAI22_X1 port map( A1 => n14197, A2 => n1751, B1 => n14194, B2 => 
                           n189, ZN => n3081);
   U2920 : OAI22_X1 port map( A1 => n14251, A2 => n2028, B1 => n14248, B2 => 
                           n1144, ZN => n3110);
   U2921 : OAI22_X1 port map( A1 => n14197, A2 => n2137, B1 => n14194, B2 => 
                           n1462, ZN => n3118);
   U2922 : OAI22_X1 port map( A1 => n363, A2 => n13807, B1 => n371, B2 => 
                           n13804, ZN => n5399);
   U2923 : OAI22_X1 port map( A1 => n361, A2 => n13807, B1 => n369, B2 => 
                           n13804, ZN => n5473);
   U2924 : OAI22_X1 port map( A1 => n360, A2 => n13807, B1 => n368, B2 => 
                           n13804, ZN => n5510);
   U2925 : OAI22_X1 port map( A1 => n359, A2 => n13807, B1 => n367, B2 => 
                           n13804, ZN => n5547);
   U2926 : OAI22_X1 port map( A1 => n358, A2 => n13807, B1 => n366, B2 => 
                           n13804, ZN => n5584);
   U2927 : OAI22_X1 port map( A1 => n364, A2 => n13807, B1 => n372, B2 => 
                           n13804, ZN => n5306);
   U2928 : OAI22_X1 port map( A1 => n362, A2 => n13807, B1 => n370, B2 => 
                           n13804, ZN => n5436);
   U2929 : OAI22_X1 port map( A1 => n357, A2 => n13807, B1 => n365, B2 => 
                           n13804, ZN => n5621);
   U2930 : OAI22_X1 port map( A1 => n390, A2 => n13973, B1 => n398, B2 => 
                           n13970, ZN => n4271);
   U2931 : OAI22_X1 port map( A1 => n299, A2 => n13834, B1 => n307, B2 => 
                           n13831, ZN => n5397);
   U2932 : OAI22_X1 port map( A1 => n259, A2 => n13780, B1 => n267, B2 => 
                           n13777, ZN => n5405);
   U2933 : OAI22_X1 port map( A1 => n395, A2 => n13753, B1 => n403, B2 => 
                           n13750, ZN => n5407);
   U2934 : OAI22_X1 port map( A1 => n297, A2 => n13834, B1 => n305, B2 => 
                           n13831, ZN => n5471);
   U2935 : OAI22_X1 port map( A1 => n257, A2 => n13780, B1 => n265, B2 => 
                           n13777, ZN => n5479);
   U2936 : OAI22_X1 port map( A1 => n393, A2 => n13753, B1 => n401, B2 => 
                           n13750, ZN => n5481);
   U2937 : OAI22_X1 port map( A1 => n296, A2 => n13834, B1 => n304, B2 => 
                           n13831, ZN => n5508);
   U2938 : OAI22_X1 port map( A1 => n256, A2 => n13780, B1 => n264, B2 => 
                           n13777, ZN => n5516);
   U2939 : OAI22_X1 port map( A1 => n392, A2 => n13753, B1 => n400, B2 => 
                           n13750, ZN => n5518);
   U2940 : OAI22_X1 port map( A1 => n295, A2 => n13834, B1 => n303, B2 => 
                           n13831, ZN => n5545);
   U2941 : OAI22_X1 port map( A1 => n255, A2 => n13780, B1 => n263, B2 => 
                           n13777, ZN => n5553);
   U2942 : OAI22_X1 port map( A1 => n391, A2 => n13753, B1 => n399, B2 => 
                           n13750, ZN => n5555);
   U2943 : OAI22_X1 port map( A1 => n294, A2 => n13834, B1 => n302, B2 => 
                           n13831, ZN => n5582);
   U2944 : OAI22_X1 port map( A1 => n254, A2 => n13780, B1 => n262, B2 => 
                           n13777, ZN => n5590);
   U2945 : OAI22_X1 port map( A1 => n390, A2 => n13753, B1 => n398, B2 => 
                           n13750, ZN => n5592);
   U2946 : OAI22_X1 port map( A1 => n396, A2 => n13973, B1 => n404, B2 => 
                           n13970, ZN => n4011);
   U2947 : OAI22_X1 port map( A1 => n300, A2 => n13834, B1 => n308, B2 => 
                           n13831, ZN => n5295);
   U2948 : OAI22_X1 port map( A1 => n260, A2 => n13780, B1 => n268, B2 => 
                           n13777, ZN => n5321);
   U2949 : OAI22_X1 port map( A1 => n396, A2 => n13753, B1 => n404, B2 => 
                           n13750, ZN => n5332);
   U2950 : OAI22_X1 port map( A1 => n395, A2 => n13973, B1 => n403, B2 => 
                           n13970, ZN => n4084);
   U2951 : OAI22_X1 port map( A1 => n394, A2 => n13973, B1 => n402, B2 => 
                           n13970, ZN => n4123);
   U2952 : OAI22_X1 port map( A1 => n298, A2 => n13834, B1 => n306, B2 => 
                           n13831, ZN => n5434);
   U2953 : OAI22_X1 port map( A1 => n258, A2 => n13780, B1 => n266, B2 => 
                           n13777, ZN => n5442);
   U2954 : OAI22_X1 port map( A1 => n394, A2 => n13753, B1 => n402, B2 => 
                           n13750, ZN => n5444);
   U2955 : OAI22_X1 port map( A1 => n393, A2 => n13973, B1 => n401, B2 => 
                           n13970, ZN => n4160);
   U2956 : OAI22_X1 port map( A1 => n392, A2 => n13973, B1 => n400, B2 => 
                           n13970, ZN => n4197);
   U2957 : OAI22_X1 port map( A1 => n391, A2 => n13973, B1 => n399, B2 => 
                           n13970, ZN => n4234);
   U2958 : OAI22_X1 port map( A1 => n389, A2 => n13973, B1 => n397, B2 => 
                           n13970, ZN => n4308);
   U2959 : OAI22_X1 port map( A1 => n293, A2 => n13834, B1 => n301, B2 => 
                           n13831, ZN => n5619);
   U2960 : OAI22_X1 port map( A1 => n253, A2 => n13780, B1 => n261, B2 => 
                           n13777, ZN => n5627);
   U2961 : OAI22_X1 port map( A1 => n389, A2 => n13753, B1 => n397, B2 => 
                           n13750, ZN => n5629);
   U2962 : OAI22_X1 port map( A1 => n1089, A2 => n14000, B1 => n1068, B2 => 
                           n13997, ZN => n4972);
   U2963 : OAI22_X1 port map( A1 => n1088, A2 => n14000, B1 => n1067, B2 => 
                           n13997, ZN => n5009);
   U2964 : OAI22_X1 port map( A1 => n1087, A2 => n14000, B1 => n1066, B2 => 
                           n13997, ZN => n5046);
   U2965 : OAI22_X1 port map( A1 => n1707, A2 => n14000, B1 => n1065, B2 => 
                           n13997, ZN => n5083);
   U2966 : OAI22_X1 port map( A1 => n1086, A2 => n14000, B1 => n1064, B2 => 
                           n13997, ZN => n5120);
   U2967 : OAI22_X1 port map( A1 => n1085, A2 => n14000, B1 => n1063, B2 => 
                           n13997, ZN => n5157);
   U2968 : OAI22_X1 port map( A1 => n262, A2 => n13998, B1 => n254, B2 => 
                           n13995, ZN => n4269);
   U2969 : OAI22_X1 port map( A1 => n1650, A2 => n13971, B1 => n1671, B2 => 
                           n13968, ZN => n5209);
   U2970 : OAI22_X1 port map( A1 => n1094, A2 => n13999, B1 => n1073, B2 => 
                           n13996, ZN => n4787);
   U2971 : OAI22_X1 port map( A1 => n1093, A2 => n13999, B1 => n1072, B2 => 
                           n13996, ZN => n4824);
   U2972 : OAI22_X1 port map( A1 => n1657, A2 => n13971, B1 => n1678, B2 => 
                           n13968, ZN => n4826);
   U2973 : OAI22_X1 port map( A1 => n1092, A2 => n13999, B1 => n1071, B2 => 
                           n13996, ZN => n4861);
   U2974 : OAI22_X1 port map( A1 => n1656, A2 => n13971, B1 => n1677, B2 => 
                           n13968, ZN => n4863);
   U2975 : OAI22_X1 port map( A1 => n1091, A2 => n13999, B1 => n1070, B2 => 
                           n13996, ZN => n4898);
   U2976 : OAI22_X1 port map( A1 => n1655, A2 => n13971, B1 => n1676, B2 => 
                           n13968, ZN => n4900);
   U2977 : OAI22_X1 port map( A1 => n1090, A2 => n13999, B1 => n1069, B2 => 
                           n13996, ZN => n4935);
   U2978 : OAI22_X1 port map( A1 => n1654, A2 => n13971, B1 => n1675, B2 => 
                           n13968, ZN => n4937);
   U2979 : OAI22_X1 port map( A1 => n495, A2 => n13832, B1 => n787, B2 => 
                           n13829, ZN => n6100);
   U2980 : OAI22_X1 port map( A1 => n591, A2 => n13805, B1 => n615, B2 => 
                           n13802, ZN => n6102);
   U2981 : OAI22_X1 port map( A1 => n1073, A2 => n13778, B1 => n1094, B2 => 
                           n13775, ZN => n6108);
   U2982 : OAI22_X1 port map( A1 => n494, A2 => n13832, B1 => n785, B2 => 
                           n13829, ZN => n6137);
   U2983 : OAI22_X1 port map( A1 => n590, A2 => n13805, B1 => n614, B2 => 
                           n13802, ZN => n6139);
   U2984 : OAI22_X1 port map( A1 => n1072, A2 => n13778, B1 => n1093, B2 => 
                           n13775, ZN => n6145);
   U2985 : OAI22_X1 port map( A1 => n1657, A2 => n13751, B1 => n1678, B2 => 
                           n13748, ZN => n6147);
   U2986 : OAI22_X1 port map( A1 => n493, A2 => n13832, B1 => n783, B2 => 
                           n13829, ZN => n6174);
   U2987 : OAI22_X1 port map( A1 => n589, A2 => n13805, B1 => n613, B2 => 
                           n13802, ZN => n6176);
   U2988 : OAI22_X1 port map( A1 => n1071, A2 => n13778, B1 => n1092, B2 => 
                           n13775, ZN => n6182);
   U2989 : OAI22_X1 port map( A1 => n1656, A2 => n13751, B1 => n1677, B2 => 
                           n13748, ZN => n6184);
   U2990 : OAI22_X1 port map( A1 => n492, A2 => n13832, B1 => n782, B2 => 
                           n13829, ZN => n6211);
   U2991 : OAI22_X1 port map( A1 => n588, A2 => n13805, B1 => n612, B2 => 
                           n13802, ZN => n6213);
   U2992 : OAI22_X1 port map( A1 => n1070, A2 => n13778, B1 => n1091, B2 => 
                           n13775, ZN => n6219);
   U2993 : OAI22_X1 port map( A1 => n1655, A2 => n13751, B1 => n1676, B2 => 
                           n13748, ZN => n6221);
   U2994 : OAI22_X1 port map( A1 => n491, A2 => n13832, B1 => n781, B2 => 
                           n13829, ZN => n6248);
   U2995 : OAI22_X1 port map( A1 => n587, A2 => n13805, B1 => n611, B2 => 
                           n13802, ZN => n6250);
   U2996 : OAI22_X1 port map( A1 => n1069, A2 => n13778, B1 => n1090, B2 => 
                           n13775, ZN => n6256);
   U2997 : OAI22_X1 port map( A1 => n1654, A2 => n13751, B1 => n1675, B2 => 
                           n13748, ZN => n6258);
   U2998 : OAI22_X1 port map( A1 => n490, A2 => n13832, B1 => n780, B2 => 
                           n13829, ZN => n6285);
   U2999 : OAI22_X1 port map( A1 => n586, A2 => n13805, B1 => n610, B2 => 
                           n13802, ZN => n6287);
   U3000 : OAI22_X1 port map( A1 => n1068, A2 => n13778, B1 => n1089, B2 => 
                           n13775, ZN => n6293);
   U3001 : OAI22_X1 port map( A1 => n1653, A2 => n13751, B1 => n1674, B2 => 
                           n13748, ZN => n6295);
   U3002 : OAI22_X1 port map( A1 => n489, A2 => n13832, B1 => n779, B2 => 
                           n13829, ZN => n6322);
   U3003 : OAI22_X1 port map( A1 => n585, A2 => n13805, B1 => n609, B2 => 
                           n13802, ZN => n6324);
   U3004 : OAI22_X1 port map( A1 => n1067, A2 => n13778, B1 => n1088, B2 => 
                           n13775, ZN => n6330);
   U3005 : OAI22_X1 port map( A1 => n1652, A2 => n13751, B1 => n1673, B2 => 
                           n13748, ZN => n6332);
   U3006 : OAI22_X1 port map( A1 => n488, A2 => n13832, B1 => n778, B2 => 
                           n13829, ZN => n6359);
   U3007 : OAI22_X1 port map( A1 => n584, A2 => n13805, B1 => n608, B2 => 
                           n13802, ZN => n6361);
   U3008 : OAI22_X1 port map( A1 => n1066, A2 => n13778, B1 => n1087, B2 => 
                           n13775, ZN => n6367);
   U3009 : OAI22_X1 port map( A1 => n1651, A2 => n13751, B1 => n1672, B2 => 
                           n13748, ZN => n6369);
   U3010 : OAI22_X1 port map( A1 => n487, A2 => n13832, B1 => n776, B2 => 
                           n13829, ZN => n6396);
   U3011 : OAI22_X1 port map( A1 => n583, A2 => n13805, B1 => n607, B2 => 
                           n13802, ZN => n6398);
   U3012 : OAI22_X1 port map( A1 => n1065, A2 => n13778, B1 => n1707, B2 => 
                           n13775, ZN => n6404);
   U3013 : OAI22_X1 port map( A1 => n1710, A2 => n13751, B1 => n1711, B2 => 
                           n13748, ZN => n6406);
   U3014 : OAI22_X1 port map( A1 => n486, A2 => n13832, B1 => n775, B2 => 
                           n13829, ZN => n6433);
   U3015 : OAI22_X1 port map( A1 => n582, A2 => n13805, B1 => n606, B2 => 
                           n13802, ZN => n6435);
   U3016 : OAI22_X1 port map( A1 => n1064, A2 => n13778, B1 => n1086, B2 => 
                           n13775, ZN => n6441);
   U3017 : OAI22_X1 port map( A1 => n1604, A2 => n13751, B1 => n1606, B2 => 
                           n13748, ZN => n6443);
   U3018 : OAI22_X1 port map( A1 => n485, A2 => n13832, B1 => n773, B2 => 
                           n13829, ZN => n6470);
   U3019 : OAI22_X1 port map( A1 => n581, A2 => n13805, B1 => n605, B2 => 
                           n13802, ZN => n6472);
   U3020 : OAI22_X1 port map( A1 => n1063, A2 => n13778, B1 => n1085, B2 => 
                           n13775, ZN => n6478);
   U3021 : OAI22_X1 port map( A1 => n1603, A2 => n13751, B1 => n1605, B2 => 
                           n13748, ZN => n6480);
   U3022 : OAI22_X1 port map( A1 => n1095, A2 => n13999, B1 => n1074, B2 => 
                           n13996, ZN => n4713);
   U3023 : OAI22_X1 port map( A1 => n1660, A2 => n13972, B1 => n1681, B2 => 
                           n13969, ZN => n4715);
   U3024 : OAI22_X1 port map( A1 => n1868, A2 => n14053, B1 => n472, B2 => 
                           n14050, ZN => n4742);
   U3025 : OAI22_X1 port map( A1 => n1892, A2 => n14026, B1 => n568, B2 => 
                           n14023, ZN => n4744);
   U3026 : OAI22_X1 port map( A1 => n497, A2 => n13833, B1 => n789, B2 => 
                           n13830, ZN => n6026);
   U3027 : OAI22_X1 port map( A1 => n593, A2 => n13806, B1 => n617, B2 => 
                           n13803, ZN => n6028);
   U3028 : OAI22_X1 port map( A1 => n1074, A2 => n13779, B1 => n1095, B2 => 
                           n13776, ZN => n6034);
   U3029 : OAI22_X1 port map( A1 => n1660, A2 => n13752, B1 => n1681, B2 => 
                           n13749, ZN => n6036);
   U3030 : OAI22_X1 port map( A1 => n484, A2 => n13832, B1 => n772, B2 => 
                           n13829, ZN => n6514);
   U3031 : OAI22_X1 port map( A1 => n580, A2 => n13805, B1 => n604, B2 => 
                           n13802, ZN => n6520);
   U3032 : OAI22_X1 port map( A1 => n1062, A2 => n13778, B1 => n1607, B2 => 
                           n13775, ZN => n6528);
   U3033 : OAI22_X1 port map( A1 => n1650, A2 => n13751, B1 => n1671, B2 => 
                           n13748, ZN => n6530);
   U3034 : OAI22_X1 port map( A1 => n1653, A2 => n13971, B1 => n1674, B2 => 
                           n13968, ZN => n4974);
   U3035 : OAI22_X1 port map( A1 => n1652, A2 => n13971, B1 => n1673, B2 => 
                           n13968, ZN => n5011);
   U3036 : OAI22_X1 port map( A1 => n1651, A2 => n13971, B1 => n1672, B2 => 
                           n13968, ZN => n5048);
   U3037 : OAI22_X1 port map( A1 => n1710, A2 => n13971, B1 => n1711, B2 => 
                           n13968, ZN => n5085);
   U3038 : OAI22_X1 port map( A1 => n1604, A2 => n13971, B1 => n1606, B2 => 
                           n13968, ZN => n5122);
   U3039 : OAI22_X1 port map( A1 => n1603, A2 => n13971, B1 => n1605, B2 => 
                           n13968, ZN => n5159);
   U3040 : OAI22_X1 port map( A1 => n14249, A2 => n1731, B1 => n14246, B2 => 
                           n1732, ZN => n6570);
   U3041 : OAI22_X1 port map( A1 => n14222, A2 => n16, B1 => n14219, B2 => n24,
                           ZN => n6575);
   U3042 : OAI22_X1 port map( A1 => n14195, A2 => n1757, B1 => n14192, B2 => 
                           n1758, ZN => n6583);
   U3043 : OAI22_X1 port map( A1 => n14169, A2 => n1741, B1 => n14165, B2 => 
                           n1742, ZN => n6585);
   U3044 : OAI22_X1 port map( A1 => n14123, A2 => n1782, B1 => n14119, B2 => 
                           n1783, ZN => n6594);
   U3045 : OAI22_X1 port map( A1 => n267, A2 => n13998, B1 => n259, B2 => 
                           n13995, ZN => n4082);
   U3046 : OAI22_X1 port map( A1 => n266, A2 => n13998, B1 => n258, B2 => 
                           n13995, ZN => n4121);
   U3047 : OAI22_X1 port map( A1 => n265, A2 => n13998, B1 => n257, B2 => 
                           n13995, ZN => n4158);
   U3048 : OAI22_X1 port map( A1 => n264, A2 => n13998, B1 => n256, B2 => 
                           n13995, ZN => n4195);
   U3049 : OAI22_X1 port map( A1 => n263, A2 => n13998, B1 => n255, B2 => 
                           n13995, ZN => n4232);
   U3050 : OAI22_X1 port map( A1 => n261, A2 => n13998, B1 => n253, B2 => 
                           n13995, ZN => n4306);
   U3051 : OAI22_X1 port map( A1 => n1105, A2 => n13999, B1 => n1084, B2 => 
                           n13996, ZN => n4343);
   U3052 : OAI22_X1 port map( A1 => n1670, A2 => n13972, B1 => n1691, B2 => 
                           n13969, ZN => n4345);
   U3053 : OAI22_X1 port map( A1 => n507, A2 => n13833, B1 => n813, B2 => 
                           n13830, ZN => n5656);
   U3054 : OAI22_X1 port map( A1 => n603, A2 => n13806, B1 => n627, B2 => 
                           n13803, ZN => n5658);
   U3055 : OAI22_X1 port map( A1 => n1084, A2 => n13779, B1 => n1105, B2 => 
                           n13776, ZN => n5664);
   U3056 : OAI22_X1 port map( A1 => n1670, A2 => n13752, B1 => n1691, B2 => 
                           n13749, ZN => n5666);
   U3057 : OAI22_X1 port map( A1 => n1104, A2 => n13998, B1 => n1083, B2 => 
                           n13995, ZN => n4380);
   U3058 : OAI22_X1 port map( A1 => n1669, A2 => n13972, B1 => n1690, B2 => 
                           n13969, ZN => n4382);
   U3059 : OAI22_X1 port map( A1 => n506, A2 => n13833, B1 => n809, B2 => 
                           n13830, ZN => n5693);
   U3060 : OAI22_X1 port map( A1 => n602, A2 => n13806, B1 => n626, B2 => 
                           n13803, ZN => n5695);
   U3061 : OAI22_X1 port map( A1 => n1083, A2 => n13779, B1 => n1104, B2 => 
                           n13776, ZN => n5701);
   U3062 : OAI22_X1 port map( A1 => n1669, A2 => n13752, B1 => n1690, B2 => 
                           n13749, ZN => n5703);
   U3063 : OAI22_X1 port map( A1 => n14250, A2 => n2027, B1 => n14247, B2 => 
                           n1143, ZN => n3147);
   U3064 : OAI22_X1 port map( A1 => n14223, A2 => n660, B1 => n14220, B2 => 
                           n684, ZN => n3149);
   U3065 : OAI22_X1 port map( A1 => n14196, A2 => n2136, B1 => n14193, B2 => 
                           n1461, ZN => n3155);
   U3066 : OAI22_X1 port map( A1 => n1103, A2 => n13998, B1 => n1082, B2 => 
                           n13995, ZN => n4417);
   U3067 : OAI22_X1 port map( A1 => n1668, A2 => n13972, B1 => n1689, B2 => 
                           n13969, ZN => n4419);
   U3068 : OAI22_X1 port map( A1 => n505, A2 => n13833, B1 => n808, B2 => 
                           n13830, ZN => n5730);
   U3069 : OAI22_X1 port map( A1 => n601, A2 => n13806, B1 => n625, B2 => 
                           n13803, ZN => n5732);
   U3070 : OAI22_X1 port map( A1 => n1082, A2 => n13779, B1 => n1103, B2 => 
                           n13776, ZN => n5738);
   U3071 : OAI22_X1 port map( A1 => n1668, A2 => n13752, B1 => n1689, B2 => 
                           n13749, ZN => n5740);
   U3072 : OAI22_X1 port map( A1 => n14250, A2 => n2026, B1 => n14247, B2 => 
                           n1142, ZN => n3184);
   U3073 : OAI22_X1 port map( A1 => n14223, A2 => n659, B1 => n14220, B2 => 
                           n683, ZN => n3186);
   U3074 : OAI22_X1 port map( A1 => n14196, A2 => n2135, B1 => n14193, B2 => 
                           n1460, ZN => n3192);
   U3075 : OAI22_X1 port map( A1 => n1102, A2 => n13998, B1 => n1081, B2 => 
                           n13995, ZN => n4454);
   U3076 : OAI22_X1 port map( A1 => n1667, A2 => n13972, B1 => n1688, B2 => 
                           n13969, ZN => n4456);
   U3077 : OAI22_X1 port map( A1 => n504, A2 => n13833, B1 => n804, B2 => 
                           n13830, ZN => n5767);
   U3078 : OAI22_X1 port map( A1 => n600, A2 => n13806, B1 => n624, B2 => 
                           n13803, ZN => n5769);
   U3079 : OAI22_X1 port map( A1 => n1081, A2 => n13779, B1 => n1102, B2 => 
                           n13776, ZN => n5775);
   U3080 : OAI22_X1 port map( A1 => n1667, A2 => n13752, B1 => n1688, B2 => 
                           n13749, ZN => n5777);
   U3081 : OAI22_X1 port map( A1 => n14250, A2 => n2025, B1 => n14247, B2 => 
                           n1141, ZN => n3221);
   U3082 : OAI22_X1 port map( A1 => n14223, A2 => n658, B1 => n14220, B2 => 
                           n682, ZN => n3223);
   U3083 : OAI22_X1 port map( A1 => n14196, A2 => n2134, B1 => n14193, B2 => 
                           n1459, ZN => n3229);
   U3084 : OAI22_X1 port map( A1 => n1101, A2 => n13998, B1 => n1080, B2 => 
                           n13995, ZN => n4491);
   U3085 : OAI22_X1 port map( A1 => n1666, A2 => n13972, B1 => n1687, B2 => 
                           n13969, ZN => n4493);
   U3086 : OAI22_X1 port map( A1 => n503, A2 => n13833, B1 => n797, B2 => 
                           n13830, ZN => n5804);
   U3087 : OAI22_X1 port map( A1 => n599, A2 => n13806, B1 => n623, B2 => 
                           n13803, ZN => n5806);
   U3088 : OAI22_X1 port map( A1 => n1080, A2 => n13779, B1 => n1101, B2 => 
                           n13776, ZN => n5812);
   U3089 : OAI22_X1 port map( A1 => n1666, A2 => n13752, B1 => n1687, B2 => 
                           n13749, ZN => n5814);
   U3090 : OAI22_X1 port map( A1 => n14250, A2 => n2024, B1 => n14247, B2 => 
                           n1140, ZN => n3258);
   U3091 : OAI22_X1 port map( A1 => n14223, A2 => n657, B1 => n14220, B2 => 
                           n681, ZN => n3260);
   U3092 : OAI22_X1 port map( A1 => n14196, A2 => n2133, B1 => n14193, B2 => 
                           n1458, ZN => n3266);
   U3093 : OAI22_X1 port map( A1 => n14123, A2 => n1564, B1 => n14120, B2 => 
                           n1570, ZN => n3276);
   U3094 : OAI22_X1 port map( A1 => n1100, A2 => n13998, B1 => n1079, B2 => 
                           n13995, ZN => n4528);
   U3095 : OAI22_X1 port map( A1 => n1665, A2 => n13972, B1 => n1686, B2 => 
                           n13969, ZN => n4530);
   U3096 : OAI22_X1 port map( A1 => n502, A2 => n13833, B1 => n796, B2 => 
                           n13830, ZN => n5841);
   U3097 : OAI22_X1 port map( A1 => n598, A2 => n13806, B1 => n622, B2 => 
                           n13803, ZN => n5843);
   U3098 : OAI22_X1 port map( A1 => n1079, A2 => n13779, B1 => n1100, B2 => 
                           n13776, ZN => n5849);
   U3099 : OAI22_X1 port map( A1 => n1665, A2 => n13752, B1 => n1686, B2 => 
                           n13749, ZN => n5851);
   U3100 : OAI22_X1 port map( A1 => n14250, A2 => n1134, B1 => n14247, B2 => 
                           n1139, ZN => n3295);
   U3101 : OAI22_X1 port map( A1 => n14223, A2 => n656, B1 => n14220, B2 => 
                           n680, ZN => n3297);
   U3102 : OAI22_X1 port map( A1 => n14196, A2 => n1452, B1 => n14193, B2 => 
                           n1457, ZN => n3303);
   U3103 : OAI22_X1 port map( A1 => n14169, A2 => n1293, B1 => n14166, B2 => 
                           n1298, ZN => n3305);
   U3104 : OAI22_X1 port map( A1 => n14123, A2 => n1563, B1 => n14120, B2 => 
                           n1569, ZN => n3315);
   U3105 : OAI22_X1 port map( A1 => n1099, A2 => n13999, B1 => n1078, B2 => 
                           n13996, ZN => n4565);
   U3106 : OAI22_X1 port map( A1 => n1664, A2 => n13972, B1 => n1685, B2 => 
                           n13969, ZN => n4567);
   U3107 : OAI22_X1 port map( A1 => n501, A2 => n13833, B1 => n794, B2 => 
                           n13830, ZN => n5878);
   U3108 : OAI22_X1 port map( A1 => n597, A2 => n13806, B1 => n621, B2 => 
                           n13803, ZN => n5880);
   U3109 : OAI22_X1 port map( A1 => n1078, A2 => n13779, B1 => n1099, B2 => 
                           n13776, ZN => n5886);
   U3110 : OAI22_X1 port map( A1 => n1664, A2 => n13752, B1 => n1685, B2 => 
                           n13749, ZN => n5888);
   U3111 : OAI22_X1 port map( A1 => n14250, A2 => n1133, B1 => n14247, B2 => 
                           n1138, ZN => n3334);
   U3112 : OAI22_X1 port map( A1 => n14223, A2 => n655, B1 => n14220, B2 => 
                           n679, ZN => n3336);
   U3113 : OAI22_X1 port map( A1 => n14196, A2 => n1451, B1 => n14193, B2 => 
                           n1456, ZN => n3342);
   U3114 : OAI22_X1 port map( A1 => n14169, A2 => n1292, B1 => n14166, B2 => 
                           n1297, ZN => n3344);
   U3115 : OAI22_X1 port map( A1 => n14123, A2 => n1562, B1 => n14120, B2 => 
                           n1568, ZN => n3352);
   U3116 : OAI22_X1 port map( A1 => n1098, A2 => n13999, B1 => n1077, B2 => 
                           n13996, ZN => n4602);
   U3117 : OAI22_X1 port map( A1 => n1663, A2 => n13972, B1 => n1684, B2 => 
                           n13969, ZN => n4604);
   U3118 : OAI22_X1 port map( A1 => n500, A2 => n13833, B1 => n793, B2 => 
                           n13830, ZN => n5915);
   U3119 : OAI22_X1 port map( A1 => n596, A2 => n13806, B1 => n620, B2 => 
                           n13803, ZN => n5917);
   U3120 : OAI22_X1 port map( A1 => n1077, A2 => n13779, B1 => n1098, B2 => 
                           n13776, ZN => n5923);
   U3121 : OAI22_X1 port map( A1 => n1663, A2 => n13752, B1 => n1684, B2 => 
                           n13749, ZN => n5925);
   U3122 : OAI22_X1 port map( A1 => n14250, A2 => n1132, B1 => n14247, B2 => 
                           n1137, ZN => n3371);
   U3123 : OAI22_X1 port map( A1 => n14223, A2 => n654, B1 => n14220, B2 => 
                           n678, ZN => n3373);
   U3124 : OAI22_X1 port map( A1 => n14196, A2 => n1450, B1 => n14193, B2 => 
                           n1455, ZN => n3379);
   U3125 : OAI22_X1 port map( A1 => n14169, A2 => n1291, B1 => n14166, B2 => 
                           n1296, ZN => n3381);
   U3126 : OAI22_X1 port map( A1 => n14123, A2 => n1561, B1 => n14120, B2 => 
                           n1567, ZN => n3389);
   U3127 : OAI22_X1 port map( A1 => n1097, A2 => n13999, B1 => n1076, B2 => 
                           n13996, ZN => n4639);
   U3128 : OAI22_X1 port map( A1 => n1662, A2 => n13972, B1 => n1683, B2 => 
                           n13969, ZN => n4641);
   U3129 : OAI22_X1 port map( A1 => n499, A2 => n13833, B1 => n792, B2 => 
                           n13830, ZN => n5952);
   U3130 : OAI22_X1 port map( A1 => n595, A2 => n13806, B1 => n619, B2 => 
                           n13803, ZN => n5954);
   U3131 : OAI22_X1 port map( A1 => n1076, A2 => n13779, B1 => n1097, B2 => 
                           n13776, ZN => n5960);
   U3132 : OAI22_X1 port map( A1 => n1662, A2 => n13752, B1 => n1683, B2 => 
                           n13749, ZN => n5962);
   U3133 : OAI22_X1 port map( A1 => n14250, A2 => n1131, B1 => n14247, B2 => 
                           n1136, ZN => n3408);
   U3134 : OAI22_X1 port map( A1 => n14223, A2 => n653, B1 => n14220, B2 => 
                           n677, ZN => n3410);
   U3135 : OAI22_X1 port map( A1 => n14196, A2 => n1449, B1 => n14193, B2 => 
                           n1454, ZN => n3416);
   U3136 : OAI22_X1 port map( A1 => n14169, A2 => n1290, B1 => n14166, B2 => 
                           n1295, ZN => n3418);
   U3137 : OAI22_X1 port map( A1 => n14123, A2 => n1560, B1 => n14120, B2 => 
                           n1566, ZN => n3426);
   U3138 : OAI22_X1 port map( A1 => n1096, A2 => n13999, B1 => n1075, B2 => 
                           n13996, ZN => n4676);
   U3139 : OAI22_X1 port map( A1 => n1661, A2 => n13972, B1 => n1682, B2 => 
                           n13969, ZN => n4678);
   U3140 : OAI22_X1 port map( A1 => n498, A2 => n13833, B1 => n790, B2 => 
                           n13830, ZN => n5989);
   U3141 : OAI22_X1 port map( A1 => n594, A2 => n13806, B1 => n618, B2 => 
                           n13803, ZN => n5991);
   U3142 : OAI22_X1 port map( A1 => n1075, A2 => n13779, B1 => n1096, B2 => 
                           n13776, ZN => n5997);
   U3143 : OAI22_X1 port map( A1 => n1661, A2 => n13752, B1 => n1682, B2 => 
                           n13749, ZN => n5999);
   U3144 : OAI22_X1 port map( A1 => n14250, A2 => n1130, B1 => n14247, B2 => 
                           n1135, ZN => n3445);
   U3145 : OAI22_X1 port map( A1 => n14223, A2 => n652, B1 => n14220, B2 => 
                           n676, ZN => n3447);
   U3146 : OAI22_X1 port map( A1 => n14196, A2 => n1448, B1 => n14193, B2 => 
                           n1453, ZN => n3453);
   U3147 : OAI22_X1 port map( A1 => n14169, A2 => n1289, B1 => n14166, B2 => 
                           n1294, ZN => n3455);
   U3148 : OAI22_X1 port map( A1 => n14250, A2 => n2023, B1 => n14247, B2 => 
                           n2042, ZN => n3482);
   U3149 : OAI22_X1 port map( A1 => n14223, A2 => n651, B1 => n14220, B2 => 
                           n675, ZN => n3484);
   U3150 : OAI22_X1 port map( A1 => n14196, A2 => n2132, B1 => n14193, B2 => 
                           n2279, ZN => n3490);
   U3151 : OAI22_X1 port map( A1 => n14169, A2 => n2080, B1 => n14166, B2 => 
                           n2094, ZN => n3492);
   U3152 : OAI22_X1 port map( A1 => n14123, A2 => n2364, B1 => n14120, B2 => 
                           n2378, ZN => n3500);
   U3153 : OAI22_X1 port map( A1 => n14250, A2 => n2022, B1 => n14247, B2 => 
                           n2041, ZN => n3519);
   U3154 : OAI22_X1 port map( A1 => n14223, A2 => n650, B1 => n14220, B2 => 
                           n674, ZN => n3521);
   U3155 : OAI22_X1 port map( A1 => n14196, A2 => n2131, B1 => n14193, B2 => 
                           n2278, ZN => n3527);
   U3156 : OAI22_X1 port map( A1 => n14169, A2 => n2079, B1 => n14166, B2 => 
                           n2093, ZN => n3529);
   U3157 : OAI22_X1 port map( A1 => n14123, A2 => n2363, B1 => n14120, B2 => 
                           n2377, ZN => n3537);
   U3158 : OAI22_X1 port map( A1 => n14250, A2 => n2021, B1 => n14247, B2 => 
                           n2040, ZN => n3556);
   U3159 : OAI22_X1 port map( A1 => n14223, A2 => n649, B1 => n14220, B2 => 
                           n673, ZN => n3558);
   U3160 : OAI22_X1 port map( A1 => n14196, A2 => n2130, B1 => n14193, B2 => 
                           n2149, ZN => n3564);
   U3161 : OAI22_X1 port map( A1 => n14169, A2 => n2078, B1 => n14166, B2 => 
                           n2092, ZN => n3566);
   U3162 : OAI22_X1 port map( A1 => n14123, A2 => n2362, B1 => n14120, B2 => 
                           n2376, ZN => n3574);
   U3163 : OAI22_X1 port map( A1 => n14249, A2 => n2020, B1 => n14246, B2 => 
                           n2039, ZN => n3593);
   U3164 : OAI22_X1 port map( A1 => n14222, A2 => n648, B1 => n14219, B2 => 
                           n672, ZN => n3595);
   U3165 : OAI22_X1 port map( A1 => n14195, A2 => n2129, B1 => n14192, B2 => 
                           n2148, ZN => n3601);
   U3166 : OAI22_X1 port map( A1 => n14169, A2 => n2077, B1 => n14165, B2 => 
                           n2091, ZN => n3603);
   U3167 : OAI22_X1 port map( A1 => n14123, A2 => n2361, B1 => n14119, B2 => 
                           n2375, ZN => n3611);
   U3168 : OAI22_X1 port map( A1 => n14249, A2 => n2019, B1 => n14246, B2 => 
                           n2038, ZN => n3630);
   U3169 : OAI22_X1 port map( A1 => n14222, A2 => n647, B1 => n14219, B2 => 
                           n671, ZN => n3632);
   U3170 : OAI22_X1 port map( A1 => n14195, A2 => n2128, B1 => n14192, B2 => 
                           n2147, ZN => n3638);
   U3171 : OAI22_X1 port map( A1 => n14169, A2 => n2076, B1 => n14165, B2 => 
                           n2090, ZN => n3640);
   U3172 : OAI22_X1 port map( A1 => n14123, A2 => n2360, B1 => n14119, B2 => 
                           n2374, ZN => n3648);
   U3173 : OAI22_X1 port map( A1 => n14249, A2 => n2018, B1 => n14246, B2 => 
                           n2037, ZN => n3667);
   U3174 : OAI22_X1 port map( A1 => n14222, A2 => n646, B1 => n14219, B2 => 
                           n670, ZN => n3669);
   U3175 : OAI22_X1 port map( A1 => n14195, A2 => n2127, B1 => n14192, B2 => 
                           n2146, ZN => n3675);
   U3176 : OAI22_X1 port map( A1 => n14169, A2 => n2075, B1 => n14165, B2 => 
                           n2089, ZN => n3677);
   U3177 : OAI22_X1 port map( A1 => n14123, A2 => n2359, B1 => n14119, B2 => 
                           n2373, ZN => n3685);
   U3178 : OAI22_X1 port map( A1 => n14249, A2 => n2017, B1 => n14246, B2 => 
                           n2036, ZN => n3704);
   U3179 : OAI22_X1 port map( A1 => n14222, A2 => n645, B1 => n14219, B2 => 
                           n669, ZN => n3706);
   U3180 : OAI22_X1 port map( A1 => n14195, A2 => n2126, B1 => n14192, B2 => 
                           n2145, ZN => n3712);
   U3181 : OAI22_X1 port map( A1 => n14170, A2 => n2074, B1 => n14165, B2 => 
                           n2088, ZN => n3714);
   U3182 : OAI22_X1 port map( A1 => n14124, A2 => n2358, B1 => n14119, B2 => 
                           n2372, ZN => n3722);
   U3183 : OAI22_X1 port map( A1 => n14249, A2 => n2016, B1 => n14246, B2 => 
                           n2035, ZN => n3741);
   U3184 : OAI22_X1 port map( A1 => n14222, A2 => n644, B1 => n14219, B2 => 
                           n668, ZN => n3743);
   U3185 : OAI22_X1 port map( A1 => n14195, A2 => n2125, B1 => n14192, B2 => 
                           n2144, ZN => n3749);
   U3186 : OAI22_X1 port map( A1 => n14170, A2 => n2073, B1 => n14165, B2 => 
                           n2087, ZN => n3751);
   U3187 : OAI22_X1 port map( A1 => n14124, A2 => n2357, B1 => n14119, B2 => 
                           n2371, ZN => n3759);
   U3188 : OAI22_X1 port map( A1 => n14249, A2 => n2015, B1 => n14246, B2 => 
                           n2034, ZN => n3778);
   U3189 : OAI22_X1 port map( A1 => n14222, A2 => n643, B1 => n14219, B2 => 
                           n667, ZN => n3780);
   U3190 : OAI22_X1 port map( A1 => n14195, A2 => n2124, B1 => n14192, B2 => 
                           n2143, ZN => n3786);
   U3191 : OAI22_X1 port map( A1 => n14170, A2 => n2072, B1 => n14165, B2 => 
                           n2086, ZN => n3788);
   U3192 : OAI22_X1 port map( A1 => n14124, A2 => n2356, B1 => n14119, B2 => 
                           n2370, ZN => n3796);
   U3193 : OAI22_X1 port map( A1 => n14249, A2 => n2014, B1 => n14246, B2 => 
                           n2033, ZN => n3815);
   U3194 : OAI22_X1 port map( A1 => n14222, A2 => n642, B1 => n14219, B2 => 
                           n666, ZN => n3817);
   U3195 : OAI22_X1 port map( A1 => n14195, A2 => n2123, B1 => n14192, B2 => 
                           n2142, ZN => n3823);
   U3196 : OAI22_X1 port map( A1 => n14170, A2 => n2071, B1 => n14165, B2 => 
                           n2085, ZN => n3825);
   U3197 : OAI22_X1 port map( A1 => n14124, A2 => n2355, B1 => n14119, B2 => 
                           n2369, ZN => n3833);
   U3198 : OAI22_X1 port map( A1 => n14249, A2 => n2013, B1 => n14246, B2 => 
                           n2032, ZN => n3852);
   U3199 : OAI22_X1 port map( A1 => n14222, A2 => n641, B1 => n14219, B2 => 
                           n665, ZN => n3854);
   U3200 : OAI22_X1 port map( A1 => n14195, A2 => n2122, B1 => n14192, B2 => 
                           n2141, ZN => n3860);
   U3201 : OAI22_X1 port map( A1 => n14170, A2 => n2070, B1 => n14165, B2 => 
                           n2084, ZN => n3862);
   U3202 : OAI22_X1 port map( A1 => n14124, A2 => n2354, B1 => n14119, B2 => 
                           n2368, ZN => n3870);
   U3203 : OAI22_X1 port map( A1 => n14249, A2 => n2012, B1 => n14246, B2 => 
                           n2031, ZN => n3889);
   U3204 : OAI22_X1 port map( A1 => n14222, A2 => n640, B1 => n14219, B2 => 
                           n664, ZN => n3891);
   U3205 : OAI22_X1 port map( A1 => n14195, A2 => n2121, B1 => n14192, B2 => 
                           n2140, ZN => n3897);
   U3206 : OAI22_X1 port map( A1 => n14170, A2 => n2069, B1 => n14165, B2 => 
                           n2083, ZN => n3899);
   U3207 : OAI22_X1 port map( A1 => n14124, A2 => n2353, B1 => n14119, B2 => 
                           n2367, ZN => n3907);
   U3208 : OAI22_X1 port map( A1 => n14249, A2 => n2011, B1 => n14246, B2 => 
                           n2030, ZN => n3926);
   U3209 : OAI22_X1 port map( A1 => n14222, A2 => n639, B1 => n14219, B2 => 
                           n663, ZN => n3928);
   U3210 : OAI22_X1 port map( A1 => n14195, A2 => n2120, B1 => n14192, B2 => 
                           n2139, ZN => n3934);
   U3211 : OAI22_X1 port map( A1 => n14170, A2 => n2068, B1 => n14165, B2 => 
                           n2082, ZN => n3936);
   U3212 : OAI22_X1 port map( A1 => n14124, A2 => n2352, B1 => n14119, B2 => 
                           n2366, ZN => n3944);
   U3213 : OAI22_X1 port map( A1 => n14249, A2 => n2010, B1 => n14246, B2 => 
                           n2029, ZN => n5248);
   U3214 : OAI22_X1 port map( A1 => n14222, A2 => n638, B1 => n14219, B2 => 
                           n662, ZN => n5250);
   U3215 : OAI22_X1 port map( A1 => n14195, A2 => n2119, B1 => n14192, B2 => 
                           n2138, ZN => n5256);
   U3216 : OAI22_X1 port map( A1 => n14169, A2 => n2067, B1 => n14165, B2 => 
                           n2081, ZN => n5258);
   U3217 : OAI22_X1 port map( A1 => n14123, A2 => n2351, B1 => n14119, B2 => 
                           n2365, ZN => n5266);
   U3218 : NAND4_X1 port map( A1 => n4737, A2 => n4738, A3 => n4739, A4 => 
                           n4740, ZN => n4736);
   U3219 : AOI221_X1 port map( B1 => n14032, B2 => n592, C1 => n14029, C2 => 
                           n616, A => n4744, ZN => n4737);
   U3220 : AOI221_X1 port map( B1 => n14059, B2 => n496, C1 => n14056, C2 => 
                           n788, A => n4742, ZN => n4739);
   U3221 : AOI221_X1 port map( B1 => n14047, B2 => n1025, C1 => n14044, C2 => 
                           n544, A => n4743, ZN => n4738);
   U3222 : NOR3_X1 port map( A1 => n2544, A2 => n2545, A3 => n2543, ZN => n5226
                           );
   U3223 : NOR3_X1 port map( A1 => n2550, A2 => n2551, A3 => n2549, ZN => n6547
                           );
   U3224 : NOR3_X2 port map( A1 => n2547, A2 => n2548, A3 => n2546, ZN => n5189
                           );
   U3225 : NOR3_X2 port map( A1 => n2553, A2 => n2554, A3 => n2552, ZN => n6510
                           );
   U3226 : OAI221_X1 port map( B1 => n2702, B2 => n6607, C1 => n14962, C2 => 
                           n13568, A => n14746, ZN => n6628);
   U3227 : OAI221_X1 port map( B1 => n14952, B2 => n13631, C1 => n2667, C2 => 
                           n6607, A => n14746, ZN => n6604);
   U3228 : OAI221_X1 port map( B1 => n14952, B2 => n14309, C1 => n2748, C2 => 
                           n14307, A => n14747, ZN => n2767);
   U3229 : OAI221_X1 port map( B1 => n14953, B2 => n13613, C1 => n2677, C2 => 
                           n6607, A => n14746, ZN => n6613);
   U3230 : OAI221_X1 port map( B1 => n14952, B2 => n14287, C1 => n2748, C2 => 
                           n14118, A => n14746, ZN => n2775);
   U3231 : OAI221_X1 port map( B1 => n14952, B2 => n14298, C1 => n2748, C2 => 
                           n14297, A => n14747, ZN => n2771);
   U3232 : OAI221_X1 port map( B1 => n14951, B2 => n14318, C1 => n2748, C2 => 
                           n2765, A => n14747, ZN => n2763);
   U3233 : OAI221_X1 port map( B1 => n14951, B2 => n14327, C1 => n2748, C2 => 
                           n2761, A => n14747, ZN => n2759);
   U3234 : OAI221_X1 port map( B1 => n14951, B2 => n14336, C1 => n2748, C2 => 
                           n2757, A => n14747, ZN => n2755);
   U3235 : OAI221_X1 port map( B1 => n14951, B2 => n14345, C1 => n2748, C2 => 
                           n2753, A => n14747, ZN => n2751);
   U3236 : OAI221_X1 port map( B1 => n14950, B2 => n14356, C1 => n2748, C2 => 
                           n14354, A => n14747, ZN => n2746);
   U3237 : OAI221_X1 port map( B1 => n14954, B2 => n13577, C1 => n2697, C2 => 
                           n6607, A => n14746, ZN => n6625);
   U3238 : OAI221_X1 port map( B1 => n14954, B2 => n13586, C1 => n2692, C2 => 
                           n6607, A => n14746, ZN => n6622);
   U3239 : OAI221_X1 port map( B1 => n14953, B2 => n13595, C1 => n2687, C2 => 
                           n6607, A => n14746, ZN => n6619);
   U3240 : OAI221_X1 port map( B1 => n14953, B2 => n13604, C1 => n2682, C2 => 
                           n6607, A => n14746, ZN => n6616);
   U3241 : OAI221_X1 port map( B1 => n14953, B2 => n13622, C1 => n2672, C2 => 
                           n6607, A => n14746, ZN => n6610);
   U3242 : NOR2_X1 port map( A1 => n2587, A2 => n2588, ZN => n6576);
   U3243 : NOR2_X1 port map( A1 => n2586, A2 => n2589, ZN => n6775);
   U3244 : NAND2_X1 port map( A1 => n2744, A2 => n2529, ZN => n2707);
   U3245 : INV_X1 port map( A => n6607, ZN => n2527);
   U3246 : NAND2_X1 port map( A1 => n2573, A2 => n6591, ZN => n3312);
   U3247 : NAND2_X1 port map( A1 => n2577, A2 => n6591, ZN => n3313);
   U3248 : NAND2_X1 port map( A1 => n5198, A2 => n5189, ZN => n3982);
   U3249 : NAND2_X1 port map( A1 => n5198, A2 => n5192, ZN => n3981);
   U3250 : NAND2_X1 port map( A1 => n5198, A2 => n5196, ZN => n3986);
   U3251 : NAND2_X1 port map( A1 => n5198, A2 => n5195, ZN => n3987);
   U3252 : NAND2_X1 port map( A1 => n6519, A2 => n6510, ZN => n5303);
   U3253 : NAND2_X1 port map( A1 => n6519, A2 => n6513, ZN => n5302);
   U3254 : NAND2_X1 port map( A1 => n6519, A2 => n6511, ZN => n5307);
   U3255 : NAND2_X1 port map( A1 => n6519, A2 => n6508, ZN => n5308);
   U3256 : NAND2_X1 port map( A1 => n5205, A2 => n5192, ZN => n4037);
   U3257 : NAND2_X1 port map( A1 => n5205, A2 => n5189, ZN => n4036);
   U3258 : NAND2_X1 port map( A1 => n5205, A2 => n5196, ZN => n3997);
   U3259 : NAND2_X1 port map( A1 => n5205, A2 => n5195, ZN => n3995);
   U3260 : NAND2_X1 port map( A1 => n5205, A2 => n5190, ZN => n3996);
   U3261 : NAND2_X1 port map( A1 => n5215, A2 => n5194, ZN => n4023);
   U3262 : NAND2_X1 port map( A1 => n5215, A2 => n5191, ZN => n4021);
   U3263 : NAND2_X1 port map( A1 => n5215, A2 => n5195, ZN => n4022);
   U3264 : NAND2_X1 port map( A1 => n5215, A2 => n5187, ZN => n4028);
   U3265 : NAND2_X1 port map( A1 => n5215, A2 => n5192, ZN => n4062);
   U3266 : NAND2_X1 port map( A1 => n5215, A2 => n5189, ZN => n4063);
   U3267 : NAND2_X1 port map( A1 => n6536, A2 => n6516, ZN => n5344);
   U3268 : NAND2_X1 port map( A1 => n6536, A2 => n6512, ZN => n5342);
   U3269 : NAND2_X1 port map( A1 => n6536, A2 => n6517, ZN => n5343);
   U3270 : NAND2_X1 port map( A1 => n6536, A2 => n6508, ZN => n5349);
   U3272 : NAND2_X1 port map( A1 => n6536, A2 => n6510, ZN => n5385);
   U3273 : NAND2_X1 port map( A1 => n6536, A2 => n6513, ZN => n5386);
   U3274 : BUF_X1 port map( A => n2521, Z => n14747);
   U3275 : BUF_X1 port map( A => n2521, Z => n14748);
   U3276 : BUF_X1 port map( A => n2521, Z => n14743);
   U3277 : BUF_X1 port map( A => n2521, Z => n14744);
   U3278 : BUF_X1 port map( A => n2521, Z => n14745);
   U3279 : BUF_X1 port map( A => n2521, Z => n14746);
   U3280 : BUF_X1 port map( A => n4043, Z => n13920);
   U3281 : INV_X1 port map( A => n2748, ZN => n2529);
   U3282 : BUF_X1 port map( A => n2799, Z => n14240);
   U3283 : BUF_X1 port map( A => n2805, Z => n14225);
   U3284 : BUF_X1 port map( A => n2799, Z => n14241);
   U3285 : NAND2_X1 port map( A1 => n6574, A2 => n6709, ZN => n2724);
   U3286 : NAND2_X1 port map( A1 => n6576, A2 => n6709, ZN => n2714);
   U3287 : BUF_X1 port map( A => n4043, Z => n13921);
   U3288 : NAND2_X1 port map( A1 => n6574, A2 => n6775, ZN => n2719);
   U3289 : NAND2_X1 port map( A1 => n5206, A2 => n5195, ZN => n4001);
   U3290 : NAND2_X1 port map( A1 => n5206, A2 => n5194, ZN => n4002);
   U3291 : NAND2_X1 port map( A1 => n5206, A2 => n5190, ZN => n4008);
   U3292 : NAND2_X1 port map( A1 => n5206, A2 => n5196, ZN => n4006);
   U3293 : NAND2_X1 port map( A1 => n5206, A2 => n5187, ZN => n4007);
   U3294 : NAND2_X1 port map( A1 => n6526, A2 => n6515, ZN => n5318);
   U3295 : NAND2_X1 port map( A1 => n6526, A2 => n6517, ZN => n5316);
   U3296 : NAND2_X1 port map( A1 => n6526, A2 => n6511, ZN => n5317);
   U3297 : NAND2_X1 port map( A1 => n6527, A2 => n6516, ZN => n5322);
   U3298 : NAND2_X1 port map( A1 => n6527, A2 => n6517, ZN => n5323);
   U3299 : NAND2_X1 port map( A1 => n6527, A2 => n6511, ZN => n5329);
   U3300 : NAND2_X1 port map( A1 => n6527, A2 => n6515, ZN => n5327);
   U3301 : NAND2_X1 port map( A1 => n6527, A2 => n6508, ZN => n5328);
   U3302 : NAND2_X1 port map( A1 => n6526, A2 => n6512, ZN => n5359);
   U3303 : NAND2_X1 port map( A1 => n6526, A2 => n6516, ZN => n5360);
   U3304 : BUF_X1 port map( A => n5374, Z => n13670);
   U3305 : BUF_X1 port map( A => n4051, Z => n13902);
   U3306 : BUF_X1 port map( A => n4051, Z => n13903);
   U3307 : BUF_X1 port map( A => n5374, Z => n13671);
   U3308 : BUF_X1 port map( A => n2639, Z => n14633);
   U3309 : BUF_X1 port map( A => n2640, Z => n14627);
   U3310 : BUF_X1 port map( A => n2641, Z => n14621);
   U3311 : BUF_X1 port map( A => n2642, Z => n14615);
   U3312 : BUF_X1 port map( A => n2643, Z => n14609);
   U3313 : BUF_X1 port map( A => n2644, Z => n14603);
   U3314 : BUF_X1 port map( A => n2645, Z => n14597);
   U3315 : BUF_X1 port map( A => n2646, Z => n14591);
   U3316 : BUF_X1 port map( A => n2647, Z => n14585);
   U3317 : BUF_X1 port map( A => n2648, Z => n14579);
   U3318 : BUF_X1 port map( A => n2649, Z => n14573);
   U3319 : BUF_X1 port map( A => n2650, Z => n14567);
   U3320 : BUF_X1 port map( A => n2651, Z => n14561);
   U3321 : BUF_X1 port map( A => n2652, Z => n14555);
   U3322 : BUF_X1 port map( A => n2653, Z => n14549);
   U3323 : BUF_X1 port map( A => n2654, Z => n14543);
   U3324 : BUF_X1 port map( A => n2655, Z => n14537);
   U3325 : BUF_X1 port map( A => n2656, Z => n14531);
   U3326 : BUF_X1 port map( A => n2657, Z => n14525);
   U3327 : BUF_X1 port map( A => n2658, Z => n14519);
   U3328 : BUF_X1 port map( A => n2659, Z => n14513);
   U3329 : BUF_X1 port map( A => n2626, Z => n14702);
   U3330 : BUF_X1 port map( A => n2627, Z => n14693);
   U3331 : BUF_X1 port map( A => n2639, Z => n14632);
   U3332 : BUF_X1 port map( A => n2640, Z => n14626);
   U3333 : BUF_X1 port map( A => n2641, Z => n14620);
   U3334 : BUF_X1 port map( A => n2642, Z => n14614);
   U3335 : BUF_X1 port map( A => n2643, Z => n14608);
   U3336 : BUF_X1 port map( A => n2644, Z => n14602);
   U3337 : BUF_X1 port map( A => n2645, Z => n14596);
   U3338 : BUF_X1 port map( A => n2646, Z => n14590);
   U3339 : BUF_X1 port map( A => n2647, Z => n14584);
   U3340 : BUF_X1 port map( A => n2648, Z => n14578);
   U3341 : BUF_X1 port map( A => n2649, Z => n14572);
   U3342 : BUF_X1 port map( A => n2650, Z => n14566);
   U3343 : BUF_X1 port map( A => n2651, Z => n14560);
   U3344 : BUF_X1 port map( A => n2652, Z => n14554);
   U3345 : BUF_X1 port map( A => n2653, Z => n14548);
   U3346 : BUF_X1 port map( A => n2654, Z => n14542);
   U3347 : BUF_X1 port map( A => n2655, Z => n14536);
   U3348 : BUF_X1 port map( A => n2656, Z => n14530);
   U3349 : BUF_X1 port map( A => n2657, Z => n14524);
   U3350 : BUF_X1 port map( A => n2658, Z => n14518);
   U3351 : BUF_X1 port map( A => n2659, Z => n14512);
   U3352 : BUF_X1 port map( A => n2626, Z => n14701);
   U3353 : BUF_X1 port map( A => n2627, Z => n14694);
   U3354 : BUF_X1 port map( A => n2627, Z => n14692);
   U3355 : BUF_X1 port map( A => n2649, Z => n14571);
   U3356 : BUF_X1 port map( A => n2650, Z => n14565);
   U3357 : BUF_X1 port map( A => n2651, Z => n14559);
   U3358 : BUF_X1 port map( A => n2652, Z => n14553);
   U3359 : BUF_X1 port map( A => n2653, Z => n14547);
   U3360 : BUF_X1 port map( A => n2654, Z => n14541);
   U3361 : BUF_X1 port map( A => n2655, Z => n14535);
   U3362 : BUF_X1 port map( A => n2656, Z => n14529);
   U3363 : BUF_X1 port map( A => n2657, Z => n14523);
   U3364 : BUF_X1 port map( A => n2658, Z => n14517);
   U3365 : BUF_X1 port map( A => n2659, Z => n14511);
   U3366 : BUF_X1 port map( A => n2639, Z => n14631);
   U3367 : BUF_X1 port map( A => n2640, Z => n14625);
   U3368 : BUF_X1 port map( A => n2641, Z => n14619);
   U3369 : BUF_X1 port map( A => n2642, Z => n14613);
   U3370 : BUF_X1 port map( A => n2643, Z => n14607);
   U3371 : BUF_X1 port map( A => n2644, Z => n14601);
   U3372 : BUF_X1 port map( A => n2645, Z => n14595);
   U3373 : BUF_X1 port map( A => n2646, Z => n14589);
   U3374 : BUF_X1 port map( A => n2647, Z => n14583);
   U3375 : BUF_X1 port map( A => n2648, Z => n14577);
   U3376 : BUF_X1 port map( A => n2627, Z => n14695);
   U3377 : BUF_X1 port map( A => n2626, Z => n14700);
   U3378 : BUF_X1 port map( A => n2639, Z => n14630);
   U3379 : BUF_X1 port map( A => n2640, Z => n14624);
   U3380 : BUF_X1 port map( A => n2641, Z => n14618);
   U3381 : BUF_X1 port map( A => n2642, Z => n14612);
   U3382 : BUF_X1 port map( A => n2643, Z => n14606);
   U3383 : BUF_X1 port map( A => n2644, Z => n14600);
   U3384 : BUF_X1 port map( A => n2645, Z => n14594);
   U3385 : BUF_X1 port map( A => n2646, Z => n14588);
   U3386 : BUF_X1 port map( A => n2647, Z => n14582);
   U3387 : BUF_X1 port map( A => n2648, Z => n14576);
   U3388 : BUF_X1 port map( A => n2649, Z => n14570);
   U3389 : BUF_X1 port map( A => n2650, Z => n14564);
   U3390 : BUF_X1 port map( A => n2651, Z => n14558);
   U3391 : BUF_X1 port map( A => n2652, Z => n14552);
   U3392 : BUF_X1 port map( A => n2653, Z => n14546);
   U3393 : BUF_X1 port map( A => n2654, Z => n14540);
   U3394 : BUF_X1 port map( A => n2655, Z => n14534);
   U3395 : BUF_X1 port map( A => n2656, Z => n14528);
   U3396 : BUF_X1 port map( A => n2657, Z => n14522);
   U3397 : BUF_X1 port map( A => n2658, Z => n14516);
   U3398 : BUF_X1 port map( A => n2659, Z => n14510);
   U3399 : BUF_X1 port map( A => n2626, Z => n14699);
   U3400 : BUF_X1 port map( A => n2627, Z => n14696);
   U3401 : BUF_X1 port map( A => n2639, Z => n14629);
   U3402 : BUF_X1 port map( A => n2640, Z => n14623);
   U3403 : BUF_X1 port map( A => n2641, Z => n14617);
   U3404 : BUF_X1 port map( A => n2642, Z => n14611);
   U3405 : BUF_X1 port map( A => n2643, Z => n14605);
   U3406 : BUF_X1 port map( A => n2644, Z => n14599);
   U3407 : BUF_X1 port map( A => n2645, Z => n14593);
   U3408 : BUF_X1 port map( A => n2646, Z => n14587);
   U3409 : BUF_X1 port map( A => n2647, Z => n14581);
   U3410 : BUF_X1 port map( A => n2648, Z => n14575);
   U3411 : BUF_X1 port map( A => n2649, Z => n14569);
   U3412 : BUF_X1 port map( A => n2650, Z => n14563);
   U3413 : BUF_X1 port map( A => n2651, Z => n14557);
   U3414 : BUF_X1 port map( A => n2652, Z => n14551);
   U3415 : BUF_X1 port map( A => n2653, Z => n14545);
   U3416 : BUF_X1 port map( A => n2654, Z => n14539);
   U3417 : BUF_X1 port map( A => n2655, Z => n14533);
   U3418 : BUF_X1 port map( A => n2656, Z => n14527);
   U3419 : BUF_X1 port map( A => n2657, Z => n14521);
   U3420 : BUF_X1 port map( A => n2658, Z => n14515);
   U3421 : BUF_X1 port map( A => n2659, Z => n14509);
   U3422 : BUF_X1 port map( A => n2626, Z => n14698);
   U3423 : BUF_X1 port map( A => n2631, Z => n14678);
   U3424 : BUF_X1 port map( A => n2632, Z => n14672);
   U3425 : BUF_X1 port map( A => n2633, Z => n14666);
   U3426 : BUF_X1 port map( A => n2634, Z => n14660);
   U3427 : BUF_X1 port map( A => n2635, Z => n14654);
   U3428 : BUF_X1 port map( A => n2636, Z => n14648);
   U3429 : BUF_X1 port map( A => n2637, Z => n14642);
   U3430 : BUF_X1 port map( A => n2638, Z => n14636);
   U3431 : BUF_X1 port map( A => n2631, Z => n14677);
   U3432 : BUF_X1 port map( A => n2632, Z => n14671);
   U3433 : BUF_X1 port map( A => n2633, Z => n14665);
   U3434 : BUF_X1 port map( A => n2634, Z => n14659);
   U3435 : BUF_X1 port map( A => n2635, Z => n14653);
   U3436 : BUF_X1 port map( A => n2636, Z => n14647);
   U3437 : BUF_X1 port map( A => n2637, Z => n14641);
   U3438 : BUF_X1 port map( A => n2638, Z => n14635);
   U3439 : BUF_X1 port map( A => n2631, Z => n14681);
   U3440 : BUF_X1 port map( A => n2632, Z => n14675);
   U3441 : BUF_X1 port map( A => n2633, Z => n14669);
   U3442 : BUF_X1 port map( A => n2634, Z => n14663);
   U3443 : BUF_X1 port map( A => n2635, Z => n14657);
   U3444 : BUF_X1 port map( A => n2636, Z => n14651);
   U3445 : BUF_X1 port map( A => n2637, Z => n14645);
   U3446 : BUF_X1 port map( A => n2638, Z => n14639);
   U3447 : BUF_X1 port map( A => n2631, Z => n14680);
   U3448 : BUF_X1 port map( A => n2632, Z => n14674);
   U3449 : BUF_X1 port map( A => n2633, Z => n14668);
   U3450 : BUF_X1 port map( A => n2634, Z => n14662);
   U3451 : BUF_X1 port map( A => n2635, Z => n14656);
   U3452 : BUF_X1 port map( A => n2636, Z => n14650);
   U3453 : BUF_X1 port map( A => n2637, Z => n14644);
   U3454 : BUF_X1 port map( A => n2638, Z => n14638);
   U3455 : BUF_X1 port map( A => n2631, Z => n14679);
   U3456 : BUF_X1 port map( A => n2632, Z => n14673);
   U3457 : BUF_X1 port map( A => n2633, Z => n14667);
   U3458 : BUF_X1 port map( A => n2634, Z => n14661);
   U3459 : BUF_X1 port map( A => n2635, Z => n14655);
   U3460 : BUF_X1 port map( A => n2636, Z => n14649);
   U3461 : BUF_X1 port map( A => n2637, Z => n14643);
   U3462 : BUF_X1 port map( A => n2638, Z => n14637);
   U3463 : BUF_X1 port map( A => n2623, Z => n14714);
   U3464 : BUF_X1 port map( A => n2623, Z => n14713);
   U3465 : BUF_X1 port map( A => n2623, Z => n14712);
   U3466 : BUF_X1 port map( A => n2623, Z => n14711);
   U3467 : BUF_X1 port map( A => n2623, Z => n14710);
   U3468 : BUF_X1 port map( A => n2803, Z => n14232);
   U3469 : BUF_X1 port map( A => n2803, Z => n14231);
   U3470 : BUF_X1 port map( A => n5275, Z => n13865);
   U3471 : BUF_X1 port map( A => n3954, Z => n14085);
   U3472 : BUF_X1 port map( A => n2623, Z => n14715);
   U3473 : BUF_X1 port map( A => n2805, Z => n14226);
   U3474 : BUF_X1 port map( A => n2627, Z => n14697);
   U3475 : BUF_X1 port map( A => n2626, Z => n14703);
   U3476 : BUF_X1 port map( A => n5375, Z => n13667);
   U3477 : BUF_X1 port map( A => n4052, Z => n13899);
   U3478 : BUF_X1 port map( A => n4052, Z => n13900);
   U3479 : BUF_X1 port map( A => n5375, Z => n13668);
   U3480 : BUF_X1 port map( A => n3954, Z => n14086);
   U3481 : BUF_X1 port map( A => n5275, Z => n13866);
   U3482 : BUF_X1 port map( A => n2659, Z => n14514);
   U3483 : BUF_X1 port map( A => n2639, Z => n14634);
   U3484 : BUF_X1 port map( A => n2640, Z => n14628);
   U3485 : BUF_X1 port map( A => n2641, Z => n14622);
   U3486 : BUF_X1 port map( A => n2642, Z => n14616);
   U3487 : BUF_X1 port map( A => n2643, Z => n14610);
   U3488 : BUF_X1 port map( A => n2644, Z => n14604);
   U3489 : BUF_X1 port map( A => n2645, Z => n14598);
   U3490 : BUF_X1 port map( A => n2646, Z => n14592);
   U3491 : BUF_X1 port map( A => n2647, Z => n14586);
   U3492 : BUF_X1 port map( A => n2648, Z => n14580);
   U3493 : BUF_X1 port map( A => n2649, Z => n14574);
   U3494 : BUF_X1 port map( A => n2650, Z => n14568);
   U3495 : BUF_X1 port map( A => n2651, Z => n14562);
   U3496 : BUF_X1 port map( A => n2652, Z => n14556);
   U3497 : BUF_X1 port map( A => n2653, Z => n14550);
   U3498 : BUF_X1 port map( A => n2654, Z => n14544);
   U3499 : BUF_X1 port map( A => n2655, Z => n14538);
   U3500 : BUF_X1 port map( A => n2656, Z => n14532);
   U3501 : BUF_X1 port map( A => n2657, Z => n14526);
   U3502 : BUF_X1 port map( A => n2658, Z => n14520);
   U3503 : BUF_X1 port map( A => n2631, Z => n14682);
   U3504 : BUF_X1 port map( A => n2632, Z => n14676);
   U3505 : BUF_X1 port map( A => n2633, Z => n14670);
   U3506 : BUF_X1 port map( A => n2634, Z => n14664);
   U3507 : BUF_X1 port map( A => n2635, Z => n14658);
   U3508 : BUF_X1 port map( A => n2636, Z => n14652);
   U3509 : BUF_X1 port map( A => n2637, Z => n14646);
   U3510 : BUF_X1 port map( A => n2638, Z => n14640);
   U3511 : BUF_X1 port map( A => n2802, Z => n14235);
   U3512 : BUF_X1 port map( A => n2802, Z => n14234);
   U3513 : NAND2_X1 port map( A1 => n5186, A2 => n5187, ZN => n3971);
   U3514 : NAND2_X1 port map( A1 => n5186, A2 => n5190, ZN => n3969);
   U3515 : NAND2_X1 port map( A1 => n5188, A2 => n5189, ZN => n3970);
   U3516 : NAND2_X1 port map( A1 => n5188, A2 => n5187, ZN => n3980);
   U3517 : NAND2_X1 port map( A1 => n5188, A2 => n5195, ZN => n3975);
   U3518 : NAND2_X1 port map( A1 => n5188, A2 => n5194, ZN => n3976);
   U3519 : NAND2_X1 port map( A1 => n5186, A2 => n5195, ZN => n4012);
   U3520 : NAND2_X1 port map( A1 => n5186, A2 => n5196, ZN => n4013);
   U3521 : NAND2_X1 port map( A1 => n5217, A2 => n5195, ZN => n4034);
   U3522 : NAND2_X1 port map( A1 => n5217, A2 => n5194, ZN => n4032);
   U3523 : NAND2_X1 port map( A1 => n5217, A2 => n5196, ZN => n4033);
   U3524 : NAND2_X1 port map( A1 => n5217, A2 => n5189, ZN => n4027);
   U3525 : NAND2_X1 port map( A1 => n6507, A2 => n6508, ZN => n5292);
   U3526 : NAND2_X1 port map( A1 => n6507, A2 => n6511, ZN => n5290);
   U3527 : NAND2_X1 port map( A1 => n6509, A2 => n6510, ZN => n5291);
   U3528 : NAND2_X1 port map( A1 => n6509, A2 => n6508, ZN => n5301);
   U3529 : NAND2_X1 port map( A1 => n6509, A2 => n6515, ZN => n5296);
   U3530 : NAND2_X1 port map( A1 => n6509, A2 => n6511, ZN => n5297);
   U3531 : NAND2_X1 port map( A1 => n6507, A2 => n6517, ZN => n5333);
   U3532 : NAND2_X1 port map( A1 => n6507, A2 => n6515, ZN => n5334);
   U3533 : NAND2_X1 port map( A1 => n6538, A2 => n6517, ZN => n5355);
   U3534 : NAND2_X1 port map( A1 => n6538, A2 => n6516, ZN => n5353);
   U3535 : NAND2_X1 port map( A1 => n6538, A2 => n6515, ZN => n5354);
   U3536 : NAND2_X1 port map( A1 => n6538, A2 => n6510, ZN => n5348);
   U3537 : NAND2_X1 port map( A1 => n14941, A2 => n2531, ZN => n5278);
   U3538 : NAND2_X1 port map( A1 => ENABLE, A2 => n2530, ZN => n3957);
   U3539 : BUF_X1 port map( A => n5371, Z => n13676);
   U3540 : BUF_X1 port map( A => n5365, Z => n13691);
   U3541 : BUF_X1 port map( A => n2798, Z => n14243);
   U3542 : BUF_X1 port map( A => n2804, Z => n14228);
   U3543 : BUF_X1 port map( A => n4042, Z => n13923);
   U3544 : BUF_X1 port map( A => n4048, Z => n13908);
   U3545 : BUF_X1 port map( A => n4042, Z => n13924);
   U3546 : BUF_X1 port map( A => n4048, Z => n13909);
   U3547 : BUF_X1 port map( A => n5365, Z => n13692);
   U3548 : BUF_X1 port map( A => n5371, Z => n13677);
   U3549 : BUF_X1 port map( A => n2798, Z => n14244);
   U3550 : BUF_X1 port map( A => n2804, Z => n14229);
   U3551 : NAND2_X1 port map( A1 => n5226, A2 => n5191, ZN => n4058);
   U3552 : NAND2_X1 port map( A1 => n5226, A2 => n5192, ZN => n4056);
   U3553 : NAND2_X1 port map( A1 => n5226, A2 => n5194, ZN => n4057);
   U3554 : NAND2_X1 port map( A1 => n6547, A2 => n6512, ZN => n5381);
   U3555 : NAND2_X1 port map( A1 => n6547, A2 => n6513, ZN => n5379);
   U3556 : NAND2_X1 port map( A1 => n6547, A2 => n6516, ZN => n5380);
   U3557 : BUF_X1 port map( A => n2808, Z => n14220);
   U3558 : BUF_X1 port map( A => n2808, Z => n14219);
   U3559 : BUF_X1 port map( A => n5366, Z => n13688);
   U3560 : BUF_X1 port map( A => n5366, Z => n13689);
   U3561 : BUF_X1 port map( A => n2807, Z => n14223);
   U3562 : BUF_X1 port map( A => n2807, Z => n14222);
   U3563 : NAND2_X1 port map( A1 => n2744, A2 => n2576, ZN => n2761);
   U3564 : NAND2_X1 port map( A1 => n2744, A2 => n2572, ZN => n2757);
   U3565 : BUF_X1 port map( A => n5370, Z => n13679);
   U3566 : BUF_X1 port map( A => n4047, Z => n13911);
   U3567 : BUF_X1 port map( A => n4047, Z => n13912);
   U3568 : BUF_X1 port map( A => n5370, Z => n13680);
   U3569 : NOR2_X1 port map( A1 => n2537, A2 => n2538, ZN => n6714);
   U3570 : BUF_X1 port map( A => n2799, Z => n14242);
   U3571 : NAND2_X1 port map( A1 => n6720, A2 => n6572, ZN => n2702);
   U3572 : BUF_X1 port map( A => n5374, Z => n13672);
   U3573 : BUF_X1 port map( A => n2803, Z => n14233);
   U3574 : BUF_X1 port map( A => n5368, Z => n13685);
   U3575 : BUF_X1 port map( A => n4045, Z => n13917);
   U3576 : BUF_X1 port map( A => n4045, Z => n13918);
   U3577 : BUF_X1 port map( A => n5368, Z => n13686);
   U3578 : NOR2_X1 port map( A1 => n2536, A2 => n2535, ZN => n6777);
   U3579 : BUF_X1 port map( A => n5369, Z => n13682);
   U3580 : BUF_X1 port map( A => n4046, Z => n13914);
   U3581 : BUF_X1 port map( A => n4046, Z => n13915);
   U3582 : BUF_X1 port map( A => n5369, Z => n13683);
   U3583 : BUF_X1 port map( A => n5375, Z => n13669);
   U3584 : BUF_X1 port map( A => n4051, Z => n13904);
   U3585 : BUF_X1 port map( A => n2802, Z => n14236);
   U3586 : BUF_X1 port map( A => n4052, Z => n13901);
   U3587 : NAND2_X1 port map( A1 => n6572, A2 => n6775, ZN => n2739);
   U3588 : BUF_X1 port map( A => n5371, Z => n13678);
   U3589 : BUF_X1 port map( A => n5365, Z => n13693);
   U3590 : NAND2_X1 port map( A1 => n6709, A2 => n6572, ZN => n2661);
   U3591 : BUF_X1 port map( A => n4048, Z => n13910);
   U3592 : BUF_X1 port map( A => n2798, Z => n14245);
   U3593 : BUF_X1 port map( A => n2804, Z => n14230);
   U3594 : BUF_X1 port map( A => n4042, Z => n13925);
   U3595 : NAND2_X1 port map( A1 => n6573, A2 => n6709, ZN => n2734);
   U3596 : BUF_X1 port map( A => n2808, Z => n14221);
   U3597 : NAND2_X1 port map( A1 => n6576, A2 => n6715, ZN => n2667);
   U3598 : NAND2_X1 port map( A1 => n5205, A2 => n5191, ZN => n4093);
   U3599 : NAND2_X1 port map( A1 => n6573, A2 => n6775, ZN => n2729);
   U3600 : NAND2_X1 port map( A1 => n6573, A2 => n6720, ZN => n2692);
   U3601 : NAND2_X1 port map( A1 => n6574, A2 => n6720, ZN => n2682);
   U3602 : BUF_X1 port map( A => n2807, Z => n14224);
   U3603 : BUF_X1 port map( A => n2805, Z => n14227);
   U3604 : BUF_X1 port map( A => n5366, Z => n13690);
   U3605 : NAND2_X1 port map( A1 => n6574, A2 => n6715, ZN => n2677);
   U3606 : NAND2_X1 port map( A1 => n6573, A2 => n6715, ZN => n2687);
   U3607 : NAND2_X1 port map( A1 => n6720, A2 => n6576, ZN => n2672);
   U3608 : NAND2_X1 port map( A1 => n6715, A2 => n6572, ZN => n2697);
   U3609 : AND2_X1 port map( A1 => n6719, A2 => n6713, ZN => n2673);
   U3610 : AND2_X1 port map( A1 => n6713, A2 => n6724, ZN => n2678);
   U3611 : AND2_X1 port map( A1 => n6713, A2 => n6707, ZN => n2683);
   U3612 : AND2_X1 port map( A1 => n6713, A2 => n6714, ZN => n2668);
   U3613 : AND2_X1 port map( A1 => n6736, A2 => n6719, ZN => n2693);
   U3614 : AND2_X1 port map( A1 => n6736, A2 => n6707, ZN => n2703);
   U3615 : AND2_X1 port map( A1 => n6736, A2 => n6724, ZN => n2698);
   U3616 : AND2_X1 port map( A1 => n6736, A2 => n6714, ZN => n2688);
   U3617 : BUF_X1 port map( A => n4047, Z => n13913);
   U3618 : BUF_X1 port map( A => n5370, Z => n13681);
   U3619 : BUF_X1 port map( A => n4045, Z => n13919);
   U3620 : BUF_X1 port map( A => n5368, Z => n13687);
   U3621 : BUF_X1 port map( A => n4046, Z => n13916);
   U3622 : BUF_X1 port map( A => n5369, Z => n13684);
   U3623 : INV_X1 port map( A => n6601, ZN => n2563);
   U3624 : NAND2_X1 port map( A1 => n2744, A2 => n2571, ZN => n2765);
   U3625 : NAND2_X1 port map( A1 => n2744, A2 => n2577, ZN => n2753);
   U3626 : BUF_X1 port map( A => n5275, Z => n13867);
   U3627 : BUF_X1 port map( A => n3954, Z => n14087);
   U3628 : AND2_X1 port map( A1 => n6708, A2 => n6724, ZN => n2740);
   U3629 : AND2_X1 port map( A1 => n2744, A2 => n2570, ZN => n13222);
   U3630 : AND2_X1 port map( A1 => n6707, A2 => n6708, ZN => n2662);
   U3631 : NAND2_X1 port map( A1 => n6601, A2 => n2578, ZN => n2870);
   U3632 : AND2_X1 port map( A1 => n6601, A2 => n2585, ZN => n13223);
   U3633 : AND2_X1 port map( A1 => n6719, A2 => n6708, ZN => n2735);
   U3634 : AND2_X1 port map( A1 => n6714, A2 => n6708, ZN => n2730);
   U3635 : AND2_X1 port map( A1 => n6777, A2 => n6707, ZN => n2725);
   U3636 : AND2_X1 port map( A1 => n6777, A2 => n6724, ZN => n2720);
   U3637 : AND2_X1 port map( A1 => n6777, A2 => n6719, ZN => n2715);
   U3638 : NAND2_X1 port map( A1 => n2584, A2 => n6591, ZN => n2852);
   U3639 : NAND2_X1 port map( A1 => n2579, A2 => n6591, ZN => n2853);
   U3640 : NAND2_X1 port map( A1 => n2583, A2 => n6591, ZN => n2851);
   U3641 : NAND2_X1 port map( A1 => n2572, A2 => n6591, ZN => n2844);
   U3642 : NAND2_X1 port map( A1 => n2576, A2 => n6591, ZN => n2842);
   U3643 : NAND2_X1 port map( A1 => n2575, A2 => n6591, ZN => n2843);
   U3644 : NAND2_X1 port map( A1 => n2574, A2 => n6591, ZN => n2876);
   U3645 : NAND2_X1 port map( A1 => n2570, A2 => n6591, ZN => n2877);
   U3646 : BUF_X1 port map( A => n4043, Z => n13922);
   U3647 : AND2_X1 port map( A1 => n2744, A2 => n2575, ZN => n13224);
   U3648 : NAND2_X1 port map( A1 => n2578, A2 => n6591, ZN => n2846);
   U3649 : NAND2_X1 port map( A1 => n2582, A2 => n6591, ZN => n2847);
   U3650 : NAND2_X1 port map( A1 => n2663, A2 => n2740, ZN => n2624);
   U3651 : NAND2_X1 port map( A1 => n2662, A2 => n2663, ZN => n2630);
   U3652 : AND2_X1 port map( A1 => n2744, A2 => n2574, ZN => n13225);
   U3653 : AND2_X1 port map( A1 => n5198, A2 => n5191, ZN => n3977);
   U3654 : AND2_X1 port map( A1 => n5198, A2 => n5194, ZN => n3978);
   U3655 : AND2_X1 port map( A1 => n5198, A2 => n5190, ZN => n3983);
   U3656 : AND2_X1 port map( A1 => n5198, A2 => n5187, ZN => n3984);
   U3657 : AND2_X1 port map( A1 => n6519, A2 => n6512, ZN => n5298);
   U3658 : AND2_X1 port map( A1 => n6519, A2 => n6516, ZN => n5299);
   U3659 : AND2_X1 port map( A1 => n6519, A2 => n6515, ZN => n5304);
   U3660 : AND2_X1 port map( A1 => n6519, A2 => n6517, ZN => n5305);
   U3661 : NAND2_X1 port map( A1 => n6685, A2 => n2698, ZN => n6751);
   U3662 : NAND2_X1 port map( A1 => n6685, A2 => n2673, ZN => n6718);
   U3663 : NAND2_X1 port map( A1 => n6685, A2 => n2735, ZN => n6700);
   U3664 : NAND2_X1 port map( A1 => n6685, A2 => n2703, ZN => n6759);
   U3665 : NAND2_X1 port map( A1 => n6685, A2 => n2693, ZN => n6747);
   U3666 : NAND2_X1 port map( A1 => n6685, A2 => n2688, ZN => n6735);
   U3667 : NAND2_X1 port map( A1 => n6685, A2 => n2683, ZN => n6730);
   U3668 : NAND2_X1 port map( A1 => n6685, A2 => n2678, ZN => n6723);
   U3669 : NAND2_X1 port map( A1 => n6685, A2 => n2668, ZN => n6712);
   U3670 : NAND2_X1 port map( A1 => n6685, A2 => n2662, ZN => n6706);
   U3671 : NAND2_X1 port map( A1 => n6685, A2 => n2740, ZN => n6703);
   U3672 : NAND2_X1 port map( A1 => n6685, A2 => n2730, ZN => n6697);
   U3673 : NAND2_X1 port map( A1 => n6685, A2 => n2725, ZN => n6694);
   U3674 : NAND2_X1 port map( A1 => n6685, A2 => n2720, ZN => n6691);
   U3675 : NAND2_X1 port map( A1 => n6685, A2 => n2715, ZN => n6688);
   U3676 : NAND2_X1 port map( A1 => n6685, A2 => n2709, ZN => n6683);
   U3677 : NAND2_X1 port map( A1 => n6634, A2 => n2688, ZN => n6670);
   U3678 : NAND2_X1 port map( A1 => n6634, A2 => n2725, ZN => n6643);
   U3679 : NAND2_X1 port map( A1 => n6634, A2 => n2703, ZN => n6679);
   U3680 : NAND2_X1 port map( A1 => n6634, A2 => n2698, ZN => n6676);
   U3681 : NAND2_X1 port map( A1 => n6634, A2 => n2693, ZN => n6673);
   U3682 : NAND2_X1 port map( A1 => n6634, A2 => n2683, ZN => n6667);
   U3683 : NAND2_X1 port map( A1 => n6634, A2 => n2678, ZN => n6664);
   U3684 : NAND2_X1 port map( A1 => n6634, A2 => n2673, ZN => n6661);
   U3685 : NAND2_X1 port map( A1 => n6634, A2 => n2668, ZN => n6658);
   U3686 : NAND2_X1 port map( A1 => n6634, A2 => n2662, ZN => n6655);
   U3687 : NAND2_X1 port map( A1 => n6634, A2 => n2740, ZN => n6652);
   U3688 : NAND2_X1 port map( A1 => n6634, A2 => n2735, ZN => n6649);
   U3689 : NAND2_X1 port map( A1 => n6634, A2 => n2730, ZN => n6646);
   U3690 : NAND2_X1 port map( A1 => n6634, A2 => n2720, ZN => n6640);
   U3691 : NAND2_X1 port map( A1 => n6634, A2 => n2715, ZN => n6637);
   U3692 : NAND2_X1 port map( A1 => n6634, A2 => n2709, ZN => n6632);
   U3693 : AND2_X1 port map( A1 => n5205, A2 => n5187, ZN => n3992);
   U3694 : AND2_X1 port map( A1 => n5215, A2 => n5190, ZN => n4019);
   U3695 : AND2_X1 port map( A1 => n5215, A2 => n5196, ZN => n4018);
   U3696 : AND2_X1 port map( A1 => n6536, A2 => n6515, ZN => n5339);
   U3697 : AND2_X1 port map( A1 => n6536, A2 => n6511, ZN => n5340);
   U3698 : NAND2_X1 port map( A1 => n2582, A2 => n6601, ZN => n2872);
   U3699 : NAND2_X1 port map( A1 => n2579, A2 => n6601, ZN => n2871);
   U3700 : NAND2_X1 port map( A1 => n2683, A2 => n2663, ZN => n2681);
   U3701 : NAND2_X1 port map( A1 => n2678, A2 => n2663, ZN => n2676);
   U3702 : NAND2_X1 port map( A1 => n2720, A2 => n2663, ZN => n6797);
   U3703 : NAND2_X1 port map( A1 => n2735, A2 => n2663, ZN => n6825);
   U3704 : NAND2_X1 port map( A1 => n2703, A2 => n2663, ZN => n2701);
   U3705 : NAND2_X1 port map( A1 => n2698, A2 => n2663, ZN => n2696);
   U3706 : NAND2_X1 port map( A1 => n2693, A2 => n2663, ZN => n2691);
   U3707 : NAND2_X1 port map( A1 => n2688, A2 => n2663, ZN => n2686);
   U3708 : NAND2_X1 port map( A1 => n2673, A2 => n2663, ZN => n2671);
   U3709 : NAND2_X1 port map( A1 => n2668, A2 => n2663, ZN => n2666);
   U3710 : NAND2_X1 port map( A1 => n2730, A2 => n2663, ZN => n6819);
   U3711 : NAND2_X1 port map( A1 => n2725, A2 => n2663, ZN => n6807);
   U3712 : NAND2_X1 port map( A1 => n2715, A2 => n2663, ZN => n6784);
   U3713 : NAND2_X1 port map( A1 => n2709, A2 => n2663, ZN => n6772);
   U3714 : AND2_X1 port map( A1 => n5206, A2 => n5189, ZN => n3993);
   U3715 : AND2_X1 port map( A1 => n5206, A2 => n5192, ZN => n3998);
   U3716 : AND2_X1 port map( A1 => n5206, A2 => n5191, ZN => n3999);
   U3717 : AND2_X1 port map( A1 => n6526, A2 => n6508, ZN => n5313);
   U3718 : AND2_X1 port map( A1 => n6527, A2 => n6510, ZN => n5314);
   U3719 : AND2_X1 port map( A1 => n6527, A2 => n6512, ZN => n5319);
   U3720 : AND2_X1 port map( A1 => n6527, A2 => n6513, ZN => n5320);
   U3721 : AND2_X1 port map( A1 => n6526, A2 => n6513, ZN => n5356);
   U3722 : AND2_X1 port map( A1 => n6526, A2 => n6510, ZN => n5357);
   U3723 : AND2_X1 port map( A1 => n5188, A2 => n5192, ZN => n3966);
   U3724 : AND2_X1 port map( A1 => n5188, A2 => n5191, ZN => n3967);
   U3725 : AND2_X1 port map( A1 => n5188, A2 => n5196, ZN => n3972);
   U3726 : AND2_X1 port map( A1 => n5188, A2 => n5190, ZN => n3973);
   U3727 : AND2_X1 port map( A1 => n5186, A2 => n5194, ZN => n4009);
   U3728 : AND2_X1 port map( A1 => n5186, A2 => n5191, ZN => n4010);
   U3729 : AND2_X1 port map( A1 => n5186, A2 => n5189, ZN => n4003);
   U3730 : AND2_X1 port map( A1 => n5186, A2 => n5192, ZN => n4004);
   U3731 : AND2_X1 port map( A1 => n5217, A2 => n5187, ZN => n4030);
   U3732 : AND2_X1 port map( A1 => n5217, A2 => n5190, ZN => n4029);
   U3733 : AND2_X1 port map( A1 => n5217, A2 => n5191, ZN => n4025);
   U3734 : AND2_X1 port map( A1 => n5217, A2 => n5192, ZN => n4024);
   U3735 : AND2_X1 port map( A1 => n6509, A2 => n6513, ZN => n5287);
   U3736 : AND2_X1 port map( A1 => n6509, A2 => n6512, ZN => n5288);
   U3737 : AND2_X1 port map( A1 => n6509, A2 => n6517, ZN => n5293);
   U3738 : AND2_X1 port map( A1 => n6509, A2 => n6516, ZN => n5294);
   U3739 : AND2_X1 port map( A1 => n6507, A2 => n6516, ZN => n5330);
   U3740 : AND2_X1 port map( A1 => n6507, A2 => n6512, ZN => n5331);
   U3741 : AND2_X1 port map( A1 => n6507, A2 => n6510, ZN => n5324);
   U3742 : AND2_X1 port map( A1 => n6507, A2 => n6513, ZN => n5325);
   U3743 : AND2_X1 port map( A1 => n6538, A2 => n6511, ZN => n5350);
   U3744 : AND2_X1 port map( A1 => n6538, A2 => n6508, ZN => n5351);
   U3745 : AND2_X1 port map( A1 => n6538, A2 => n6513, ZN => n5345);
   U3746 : AND2_X1 port map( A1 => n6538, A2 => n6512, ZN => n5346);
   U3747 : AND2_X1 port map( A1 => n6547, A2 => n6508, ZN => n5382);
   U3748 : AND2_X1 port map( A1 => n5226, A2 => n5196, ZN => n4054);
   U3749 : AND2_X1 port map( A1 => n5226, A2 => n5195, ZN => n4053);
   U3750 : AND2_X1 port map( A1 => n5226, A2 => n5187, ZN => n4060);
   U3751 : AND2_X1 port map( A1 => n5226, A2 => n5190, ZN => n4059);
   U3752 : AND2_X1 port map( A1 => n6547, A2 => n6517, ZN => n5376);
   U3753 : AND2_X1 port map( A1 => n6547, A2 => n6515, ZN => n5377);
   U3754 : AND2_X1 port map( A1 => n6547, A2 => n6511, ZN => n5383);
   U3755 : NAND2_X1 port map( A1 => n6569, A2 => n2578, ZN => n2792);
   U3756 : NAND2_X1 port map( A1 => n6569, A2 => n2577, ZN => n2791);
   U3757 : NAND2_X1 port map( A1 => n6569, A2 => n2585, ZN => n2790);
   U3758 : NAND2_X1 port map( A1 => n6569, A2 => n2581, ZN => n2801);
   U3759 : NAND2_X1 port map( A1 => n6569, A2 => n2580, ZN => n2797);
   U3760 : NAND2_X1 port map( A1 => n6569, A2 => n2584, ZN => n2796);
   U3761 : NAND2_X1 port map( A1 => n6582, A2 => n2572, ZN => n2818);
   U3762 : NAND2_X1 port map( A1 => n6582, A2 => n2576, ZN => n2816);
   U3763 : NAND2_X1 port map( A1 => n6582, A2 => n2577, ZN => n2817);
   U3764 : NAND2_X1 port map( A1 => n6582, A2 => n2581, ZN => n2829);
   U3765 : NAND2_X1 port map( A1 => n6582, A2 => n2584, ZN => n2828);
   U3766 : NAND2_X1 port map( A1 => n6569, A2 => n2574, ZN => n2827);
   U3767 : NAND2_X1 port map( A1 => n6582, A2 => n2579, ZN => n2823);
   U3768 : NAND2_X1 port map( A1 => n6582, A2 => n2583, ZN => n2822);
   U3769 : NAND2_X1 port map( A1 => n6569, A2 => n2572, ZN => n2833);
   U3770 : NAND2_X1 port map( A1 => n6569, A2 => n2576, ZN => n2834);
   U3771 : NAND2_X1 port map( A1 => n6582, A2 => n2571, ZN => n2857);
   U3772 : NAND2_X1 port map( A1 => n6582, A2 => n2575, ZN => n2858);
   U3773 : NAND2_X1 port map( A1 => n6608, A2 => n2668, ZN => n6606);
   U3774 : NAND2_X1 port map( A1 => n6608, A2 => n2678, ZN => n6614);
   U3775 : NAND2_X1 port map( A1 => n6608, A2 => n2703, ZN => n6629);
   U3776 : NAND2_X1 port map( A1 => n6608, A2 => n2698, ZN => n6626);
   U3777 : NAND2_X1 port map( A1 => n6608, A2 => n2693, ZN => n6623);
   U3778 : NAND2_X1 port map( A1 => n6608, A2 => n2688, ZN => n6620);
   U3779 : NAND2_X1 port map( A1 => n6608, A2 => n2683, ZN => n6617);
   U3780 : NAND2_X1 port map( A1 => n6608, A2 => n2673, ZN => n6611);
   U3781 : AND2_X1 port map( A1 => n2580, A2 => n6591, ZN => n2849);
   U3782 : AND2_X1 port map( A1 => n2585, A2 => n6591, ZN => n2839);
   U3783 : AND2_X1 port map( A1 => n2571, A2 => n6591, ZN => n2840);
   U3784 : AND2_X1 port map( A1 => n2581, A2 => n6591, ZN => n2855);
   U3785 : AND2_X1 port map( A1 => n6569, A2 => n2573, ZN => n2788);
   U3786 : AND2_X1 port map( A1 => n6569, A2 => n2583, ZN => n2787);
   U3787 : AND2_X1 port map( A1 => n6569, A2 => n2582, ZN => n2794);
   U3788 : AND2_X1 port map( A1 => n6569, A2 => n2579, ZN => n2793);
   U3789 : AND2_X1 port map( A1 => n6582, A2 => n2573, ZN => n2814);
   U3790 : AND2_X1 port map( A1 => n6582, A2 => n2582, ZN => n2813);
   U3791 : AND2_X1 port map( A1 => n6582, A2 => n2580, ZN => n2825);
   U3792 : AND2_X1 port map( A1 => n6569, A2 => n2571, ZN => n2824);
   U3793 : AND2_X1 port map( A1 => n6582, A2 => n2585, ZN => n2820);
   U3794 : AND2_X1 port map( A1 => n6582, A2 => n2578, ZN => n2819);
   U3795 : AND2_X1 port map( A1 => n6569, A2 => n2570, ZN => n2831);
   U3796 : AND2_X1 port map( A1 => n6569, A2 => n2575, ZN => n2830);
   U3797 : AND2_X1 port map( A1 => n6582, A2 => n2570, ZN => n2848);
   U3798 : AND2_X1 port map( A1 => n6582, A2 => n2574, ZN => n2854);
   U3799 : BUF_X1 port map( A => n2778, Z => n14275);
   U3800 : BUF_X1 port map( A => n2778, Z => n14273);
   U3801 : BUF_X1 port map( A => n2778, Z => n14274);
   U3802 : INV_X1 port map( A => n14941, ZN => n14966);
   U3803 : AOI221_X1 port map( B1 => n7108, B2 => n14728, C1 => n833, C2 => 
                           n14725, A => n6599, ZN => n6598);
   U3804 : OAI222_X1 port map( A1 => n14118, A2 => n372, B1 => n7684, B2 => 
                           n14307, C1 => n14296, C2 => n364, ZN => n6599);
   U3805 : AOI221_X1 port map( B1 => n6771, B2 => n14728, C1 => n837, C2 => 
                           n14727, A => n2911, ZN => n2910);
   U3806 : OAI222_X1 port map( A1 => n14118, A2 => n370, B1 => n7672, B2 => 
                           n14307, C1 => n14296, C2 => n362, ZN => n2911);
   U3807 : AOI221_X1 port map( B1 => n6778, B2 => n14728, C1 => n839, C2 => 
                           n14727, A => n2948, ZN => n2947);
   U3808 : OAI222_X1 port map( A1 => n14117, A2 => n369, B1 => n7666, B2 => 
                           n14307, C1 => n14296, C2 => n361, ZN => n2948);
   U3809 : AOI221_X1 port map( B1 => n6787, B2 => n14728, C1 => n841, C2 => 
                           n14727, A => n2985, ZN => n2984);
   U3810 : OAI222_X1 port map( A1 => n14118, A2 => n368, B1 => n7660, B2 => 
                           n14307, C1 => n14296, C2 => n360, ZN => n2985);
   U3811 : AOI221_X1 port map( B1 => n6799, B2 => n14728, C1 => n843, C2 => 
                           n14727, A => n3022, ZN => n3021);
   U3812 : OAI222_X1 port map( A1 => n14117, A2 => n367, B1 => n7654, B2 => 
                           n14307, C1 => n14296, C2 => n359, ZN => n3022);
   U3813 : AOI221_X1 port map( B1 => n6817, B2 => n14728, C1 => n845, C2 => 
                           n14727, A => n3059, ZN => n3058);
   U3814 : OAI222_X1 port map( A1 => n14118, A2 => n366, B1 => n7648, B2 => 
                           n14307, C1 => n14296, C2 => n358, ZN => n3059);
   U3815 : AOI221_X1 port map( B1 => n6826, B2 => n14728, C1 => n847, C2 => 
                           n14727, A => n3096, ZN => n3095);
   U3816 : OAI222_X1 port map( A1 => n14117, A2 => n365, B1 => n7642, B2 => 
                           n14307, C1 => n14296, C2 => n357, ZN => n3096);
   U3817 : AOI221_X1 port map( B1 => n6853, B2 => n14728, C1 => n851, C2 => 
                           n14726, A => n3170, ZN => n3169);
   U3818 : OAI222_X1 port map( A1 => n14118, A2 => n626, B1 => n7630, B2 => 
                           n14307, C1 => n14296, C2 => n602, ZN => n3170);
   U3819 : AOI221_X1 port map( B1 => n6868, B2 => n14728, C1 => n853, C2 => 
                           n14726, A => n3207, ZN => n3206);
   U3820 : OAI222_X1 port map( A1 => n14117, A2 => n625, B1 => n7624, B2 => 
                           n14308, C1 => n14296, C2 => n601, ZN => n3207);
   U3821 : AOI221_X1 port map( B1 => n6880, B2 => n14729, C1 => n855, C2 => 
                           n14726, A => n3244, ZN => n3243);
   U3822 : OAI222_X1 port map( A1 => n14118, A2 => n624, B1 => n7618, B2 => 
                           n14307, C1 => n14296, C2 => n600, ZN => n3244);
   U3823 : AOI221_X1 port map( B1 => n8893, B2 => n13925, C1 => n8861, C2 => 
                           n13920, A => n4044, ZN => n4041);
   U3824 : OAI222_X1 port map( A1 => n6726, A2 => n13919, B1 => n6728, B2 => 
                           n13916, C1 => n6727, C2 => n13913, ZN => n4044);
   U3825 : AOI221_X1 port map( B1 => n13693, B2 => n8893, C1 => n13690, C2 => 
                           n8861, A => n5367, ZN => n5364);
   U3826 : OAI222_X1 port map( A1 => n6726, A2 => n13687, B1 => n6728, B2 => 
                           n13684, C1 => n6727, C2 => n13681, ZN => n5367);
   U3827 : OAI222_X1 port map( A1 => n6885, A2 => n13988, B1 => n6887, B2 => 
                           n13985, C1 => n6886, C2 => n13982, ZN => n4270);
   U3828 : OAI222_X1 port map( A1 => n6765, A2 => n13768, B1 => n6767, B2 => 
                           n13765, C1 => n6766, C2 => n13762, ZN => n5406);
   U3829 : OAI222_X1 port map( A1 => n6813, A2 => n13768, B1 => n6815, B2 => 
                           n13765, C1 => n6814, C2 => n13762, ZN => n5480);
   U3830 : OAI222_X1 port map( A1 => n6837, A2 => n13768, B1 => n6839, B2 => 
                           n13765, C1 => n6838, C2 => n13762, ZN => n5517);
   U3831 : OAI222_X1 port map( A1 => n6861, A2 => n13768, B1 => n6863, B2 => 
                           n13765, C1 => n6862, C2 => n13762, ZN => n5554);
   U3832 : OAI222_X1 port map( A1 => n6885, A2 => n13768, B1 => n6887, B2 => 
                           n13765, C1 => n6886, C2 => n13762, ZN => n5591);
   U3833 : OAI222_X1 port map( A1 => n7488, A2 => n14067, B1 => n7490, B2 => 
                           n14064, C1 => n7489, C2 => n14061, ZN => n5185);
   U3834 : OAI222_X1 port map( A1 => n7485, A2 => n13986, B1 => n7487, B2 => 
                           n13983, C1 => n7486, C2 => n13980, ZN => n5208);
   U3835 : OAI222_X1 port map( A1 => n7248, A2 => n14067, B1 => n7250, B2 => 
                           n14064, C1 => n7249, C2 => n14061, ZN => n4815);
   U3836 : OAI222_X1 port map( A1 => n7245, A2 => n13986, B1 => n7247, B2 => 
                           n13983, C1 => n7246, C2 => n13980, ZN => n4825);
   U3837 : OAI222_X1 port map( A1 => n7272, A2 => n14067, B1 => n7274, B2 => 
                           n14064, C1 => n7273, C2 => n14061, ZN => n4852);
   U3838 : OAI222_X1 port map( A1 => n7269, A2 => n13986, B1 => n7271, B2 => 
                           n13983, C1 => n7270, C2 => n13980, ZN => n4862);
   U3839 : OAI222_X1 port map( A1 => n7296, A2 => n14067, B1 => n7298, B2 => 
                           n14064, C1 => n7297, C2 => n14061, ZN => n4889);
   U3840 : OAI222_X1 port map( A1 => n7293, A2 => n13986, B1 => n7295, B2 => 
                           n13983, C1 => n7294, C2 => n13980, ZN => n4899);
   U3841 : OAI222_X1 port map( A1 => n7320, A2 => n14067, B1 => n7322, B2 => 
                           n14064, C1 => n7321, C2 => n14061, ZN => n4926);
   U3842 : OAI222_X1 port map( A1 => n7317, A2 => n13986, B1 => n7319, B2 => 
                           n13983, C1 => n7318, C2 => n13980, ZN => n4936);
   U3843 : OAI222_X1 port map( A1 => n7248, A2 => n13847, B1 => n7250, B2 => 
                           n13844, C1 => n7249, C2 => n13841, ZN => n6136);
   U3844 : OAI222_X1 port map( A1 => n7245, A2 => n13766, B1 => n7247, B2 => 
                           n13763, C1 => n7246, C2 => n13760, ZN => n6146);
   U3845 : OAI222_X1 port map( A1 => n7272, A2 => n13847, B1 => n7274, B2 => 
                           n13844, C1 => n7273, C2 => n13841, ZN => n6173);
   U3846 : OAI222_X1 port map( A1 => n7269, A2 => n13766, B1 => n7271, B2 => 
                           n13763, C1 => n7270, C2 => n13760, ZN => n6183);
   U3847 : OAI222_X1 port map( A1 => n7296, A2 => n13847, B1 => n7298, B2 => 
                           n13844, C1 => n7297, C2 => n13841, ZN => n6210);
   U3848 : OAI222_X1 port map( A1 => n7293, A2 => n13766, B1 => n7295, B2 => 
                           n13763, C1 => n7294, C2 => n13760, ZN => n6220);
   U3849 : OAI222_X1 port map( A1 => n7320, A2 => n13847, B1 => n7322, B2 => 
                           n13844, C1 => n7321, C2 => n13841, ZN => n6247);
   U3850 : OAI222_X1 port map( A1 => n7317, A2 => n13766, B1 => n7319, B2 => 
                           n13763, C1 => n7318, C2 => n13760, ZN => n6257);
   U3851 : OAI222_X1 port map( A1 => n7344, A2 => n13847, B1 => n7346, B2 => 
                           n13844, C1 => n7345, C2 => n13841, ZN => n6284);
   U3852 : OAI222_X1 port map( A1 => n7341, A2 => n13766, B1 => n7343, B2 => 
                           n13763, C1 => n7342, C2 => n13760, ZN => n6294);
   U3853 : OAI222_X1 port map( A1 => n7368, A2 => n13847, B1 => n7370, B2 => 
                           n13844, C1 => n7369, C2 => n13841, ZN => n6321);
   U3854 : OAI222_X1 port map( A1 => n7365, A2 => n13766, B1 => n7367, B2 => 
                           n13763, C1 => n7366, C2 => n13760, ZN => n6331);
   U3855 : OAI222_X1 port map( A1 => n7392, A2 => n13847, B1 => n7394, B2 => 
                           n13844, C1 => n7393, C2 => n13841, ZN => n6358);
   U3856 : OAI222_X1 port map( A1 => n7389, A2 => n13766, B1 => n7391, B2 => 
                           n13763, C1 => n7390, C2 => n13760, ZN => n6368);
   U3857 : OAI222_X1 port map( A1 => n7416, A2 => n13847, B1 => n7418, B2 => 
                           n13844, C1 => n7417, C2 => n13841, ZN => n6395);
   U3858 : OAI222_X1 port map( A1 => n7413, A2 => n13766, B1 => n7415, B2 => 
                           n13763, C1 => n7414, C2 => n13760, ZN => n6405);
   U3859 : OAI222_X1 port map( A1 => n7440, A2 => n13847, B1 => n7442, B2 => 
                           n13844, C1 => n7441, C2 => n13841, ZN => n6432);
   U3860 : OAI222_X1 port map( A1 => n7437, A2 => n13766, B1 => n7439, B2 => 
                           n13763, C1 => n7438, C2 => n13760, ZN => n6442);
   U3861 : OAI222_X1 port map( A1 => n7464, A2 => n13847, B1 => n7466, B2 => 
                           n13844, C1 => n7465, C2 => n13841, ZN => n6469);
   U3862 : OAI222_X1 port map( A1 => n7461, A2 => n13766, B1 => n7463, B2 => 
                           n13763, C1 => n7462, C2 => n13760, ZN => n6479);
   U3863 : OAI222_X1 port map( A1 => n7176, A2 => n14068, B1 => n7178, B2 => 
                           n14065, C1 => n7177, C2 => n14062, ZN => n4704);
   U3864 : OAI222_X1 port map( A1 => n7173, A2 => n13987, B1 => n7175, B2 => 
                           n13984, C1 => n7174, C2 => n13981, ZN => n4714);
   U3865 : OAI222_X1 port map( A1 => n7176, A2 => n13848, B1 => n7178, B2 => 
                           n13845, C1 => n7177, C2 => n13842, ZN => n6025);
   U3866 : OAI222_X1 port map( A1 => n7173, A2 => n13767, B1 => n7175, B2 => 
                           n13764, C1 => n7174, C2 => n13761, ZN => n6035);
   U3867 : OAI222_X1 port map( A1 => n7488, A2 => n13847, B1 => n7490, B2 => 
                           n13844, C1 => n7489, C2 => n13841, ZN => n6506);
   U3868 : OAI222_X1 port map( A1 => n7485, A2 => n13766, B1 => n7487, B2 => 
                           n13763, C1 => n7486, C2 => n13760, ZN => n6529);
   U3869 : OAI222_X1 port map( A1 => n7344, A2 => n14067, B1 => n7346, B2 => 
                           n14064, C1 => n7345, C2 => n14061, ZN => n4963);
   U3870 : OAI222_X1 port map( A1 => n7341, A2 => n13986, B1 => n7343, B2 => 
                           n13983, C1 => n7342, C2 => n13980, ZN => n4973);
   U3871 : OAI222_X1 port map( A1 => n7368, A2 => n14067, B1 => n7370, B2 => 
                           n14064, C1 => n7369, C2 => n14061, ZN => n5000);
   U3872 : OAI222_X1 port map( A1 => n7365, A2 => n13986, B1 => n7367, B2 => 
                           n13983, C1 => n7366, C2 => n13980, ZN => n5010);
   U3873 : OAI222_X1 port map( A1 => n7392, A2 => n14067, B1 => n7394, B2 => 
                           n14064, C1 => n7393, C2 => n14061, ZN => n5037);
   U3874 : OAI222_X1 port map( A1 => n7389, A2 => n13986, B1 => n7391, B2 => 
                           n13983, C1 => n7390, C2 => n13980, ZN => n5047);
   U3875 : OAI222_X1 port map( A1 => n7416, A2 => n14067, B1 => n7418, B2 => 
                           n14064, C1 => n7417, C2 => n14061, ZN => n5074);
   U3876 : OAI222_X1 port map( A1 => n7413, A2 => n13986, B1 => n7415, B2 => 
                           n13983, C1 => n7414, C2 => n13980, ZN => n5084);
   U3877 : OAI222_X1 port map( A1 => n7440, A2 => n14067, B1 => n7442, B2 => 
                           n14064, C1 => n7441, C2 => n14061, ZN => n5111);
   U3878 : OAI222_X1 port map( A1 => n7437, A2 => n13986, B1 => n7439, B2 => 
                           n13983, C1 => n7438, C2 => n13980, ZN => n5121);
   U3879 : OAI222_X1 port map( A1 => n7464, A2 => n14067, B1 => n7466, B2 => 
                           n14064, C1 => n7465, C2 => n14061, ZN => n5148);
   U3880 : OAI222_X1 port map( A1 => n7461, A2 => n13986, B1 => n7463, B2 => 
                           n13983, C1 => n7462, C2 => n13980, ZN => n5158);
   U3881 : OAI222_X1 port map( A1 => n6744, A2 => n14069, B1 => n6746, B2 => 
                           n14066, C1 => n6745, C2 => n14063, ZN => n3968);
   U3882 : OAI222_X1 port map( A1 => n6741, A2 => n13988, B1 => n6743, B2 => 
                           n13985, C1 => n6742, C2 => n13982, ZN => n4005);
   U3883 : OAI222_X1 port map( A1 => n6744, A2 => n13849, B1 => n6746, B2 => 
                           n13846, C1 => n6745, C2 => n13843, ZN => n5289);
   U3884 : OAI222_X1 port map( A1 => n6741, A2 => n13768, B1 => n6743, B2 => 
                           n13765, C1 => n6742, C2 => n13762, ZN => n5326);
   U3885 : OAI222_X1 port map( A1 => n6765, A2 => n13988, B1 => n6767, B2 => 
                           n13985, C1 => n6766, C2 => n13982, ZN => n4083);
   U3886 : OAI222_X1 port map( A1 => n6789, A2 => n13988, B1 => n6791, B2 => 
                           n13985, C1 => n6790, C2 => n13982, ZN => n4122);
   U3887 : OAI222_X1 port map( A1 => n6789, A2 => n13768, B1 => n6791, B2 => 
                           n13765, C1 => n6790, C2 => n13762, ZN => n5443);
   U3888 : OAI222_X1 port map( A1 => n6813, A2 => n13988, B1 => n6815, B2 => 
                           n13985, C1 => n6814, C2 => n13982, ZN => n4159);
   U3889 : OAI222_X1 port map( A1 => n6837, A2 => n13988, B1 => n6839, B2 => 
                           n13985, C1 => n6838, C2 => n13982, ZN => n4196);
   U3890 : OAI222_X1 port map( A1 => n6861, A2 => n13988, B1 => n6863, B2 => 
                           n13985, C1 => n6862, C2 => n13982, ZN => n4233);
   U3891 : OAI222_X1 port map( A1 => n6909, A2 => n13988, B1 => n6911, B2 => 
                           n13985, C1 => n6910, C2 => n13982, ZN => n4307);
   U3892 : OAI222_X1 port map( A1 => n6909, A2 => n13768, B1 => n6911, B2 => 
                           n13765, C1 => n6910, C2 => n13762, ZN => n5628);
   U3893 : OAI222_X1 port map( A1 => n6933, A2 => n13987, B1 => n6935, B2 => 
                           n13984, C1 => n6934, C2 => n13981, ZN => n4344);
   U3894 : OAI222_X1 port map( A1 => n6933, A2 => n13767, B1 => n6935, B2 => 
                           n13764, C1 => n6934, C2 => n13761, ZN => n5665);
   U3895 : OAI222_X1 port map( A1 => n6957, A2 => n13987, B1 => n6959, B2 => 
                           n13984, C1 => n6958, C2 => n13981, ZN => n4381);
   U3896 : OAI222_X1 port map( A1 => n6957, A2 => n13767, B1 => n6959, B2 => 
                           n13764, C1 => n6958, C2 => n13761, ZN => n5702);
   U3897 : OAI222_X1 port map( A1 => n6981, A2 => n13987, B1 => n6983, B2 => 
                           n13984, C1 => n6982, C2 => n13981, ZN => n4418);
   U3898 : OAI222_X1 port map( A1 => n6981, A2 => n13767, B1 => n6983, B2 => 
                           n13764, C1 => n6982, C2 => n13761, ZN => n5739);
   U3899 : OAI222_X1 port map( A1 => n7005, A2 => n13987, B1 => n7007, B2 => 
                           n13984, C1 => n7006, C2 => n13981, ZN => n4455);
   U3900 : OAI222_X1 port map( A1 => n7005, A2 => n13767, B1 => n7007, B2 => 
                           n13764, C1 => n7006, C2 => n13761, ZN => n5776);
   U3901 : OAI222_X1 port map( A1 => n7029, A2 => n13987, B1 => n7031, B2 => 
                           n13984, C1 => n7030, C2 => n13981, ZN => n4492);
   U3902 : OAI222_X1 port map( A1 => n7029, A2 => n13767, B1 => n7031, B2 => 
                           n13764, C1 => n7030, C2 => n13761, ZN => n5813);
   U3903 : OAI222_X1 port map( A1 => n1715, A2 => n13987, B1 => n7055, B2 => 
                           n13984, C1 => n7054, C2 => n13981, ZN => n4529);
   U3904 : OAI222_X1 port map( A1 => n1715, A2 => n13767, B1 => n7055, B2 => 
                           n13764, C1 => n7054, C2 => n13761, ZN => n5850);
   U3905 : OAI222_X1 port map( A1 => n1714, A2 => n13987, B1 => n7079, B2 => 
                           n13984, C1 => n7078, C2 => n13981, ZN => n4566);
   U3906 : OAI222_X1 port map( A1 => n1714, A2 => n13767, B1 => n7079, B2 => 
                           n13764, C1 => n7078, C2 => n13761, ZN => n5887);
   U3907 : OAI222_X1 port map( A1 => n1713, A2 => n13987, B1 => n7103, B2 => 
                           n13984, C1 => n7102, C2 => n13981, ZN => n4603);
   U3908 : OAI222_X1 port map( A1 => n1713, A2 => n13767, B1 => n7103, B2 => 
                           n13764, C1 => n7102, C2 => n13761, ZN => n5924);
   U3909 : OAI222_X1 port map( A1 => n1712, A2 => n13987, B1 => n7127, B2 => 
                           n13984, C1 => n7126, C2 => n13981, ZN => n4640);
   U3910 : OAI222_X1 port map( A1 => n1712, A2 => n13767, B1 => n7127, B2 => 
                           n13764, C1 => n7126, C2 => n13761, ZN => n5961);
   U3911 : OAI222_X1 port map( A1 => n7149, A2 => n13987, B1 => n7151, B2 => 
                           n13984, C1 => n7150, C2 => n13981, ZN => n4677);
   U3912 : OAI222_X1 port map( A1 => n7149, A2 => n13767, B1 => n7151, B2 => 
                           n13764, C1 => n7150, C2 => n13761, ZN => n5998);
   U3913 : OAI222_X1 port map( A1 => n829, A2 => n14139, B1 => n7851, B2 => 
                           n14135, C1 => n828, C2 => n14133, ZN => n3536);
   U3914 : OAI222_X1 port map( A1 => n7814, A2 => n14156, B1 => n404, B2 => 
                           n14153, C1 => n7815, C2 => n14150, ZN => n6590);
   U3915 : OAI222_X1 port map( A1 => n7810, A2 => n14158, B1 => n403, B2 => 
                           n14155, C1 => n7811, C2 => n14152, ZN => n2841);
   U3916 : OAI222_X1 port map( A1 => n7806, A2 => n14158, B1 => n402, B2 => 
                           n14155, C1 => n7807, C2 => n14152, ZN => n2903);
   U3917 : OAI222_X1 port map( A1 => n7802, A2 => n14158, B1 => n401, B2 => 
                           n14155, C1 => n7803, C2 => n14152, ZN => n2940);
   U3918 : OAI222_X1 port map( A1 => n7798, A2 => n14158, B1 => n400, B2 => 
                           n14155, C1 => n7799, C2 => n14152, ZN => n2977);
   U3919 : OAI222_X1 port map( A1 => n7794, A2 => n14158, B1 => n399, B2 => 
                           n14155, C1 => n7795, C2 => n14152, ZN => n3014);
   U3920 : OAI222_X1 port map( A1 => n7790, A2 => n14158, B1 => n398, B2 => 
                           n14155, C1 => n7791, C2 => n14152, ZN => n3051);
   U3921 : OAI222_X1 port map( A1 => n7786, A2 => n14158, B1 => n397, B2 => 
                           n14155, C1 => n7787, C2 => n14152, ZN => n3088);
   U3922 : OAI222_X1 port map( A1 => n7782, A2 => n14158, B1 => n1691, B2 => 
                           n14155, C1 => n7783, C2 => n14152, ZN => n3125);
   U3923 : OAI222_X1 port map( A1 => n7778, A2 => n14157, B1 => n1690, B2 => 
                           n14154, C1 => n7779, C2 => n14151, ZN => n3162);
   U3924 : OAI222_X1 port map( A1 => n7774, A2 => n14157, B1 => n1689, B2 => 
                           n14154, C1 => n7775, C2 => n14151, ZN => n3199);
   U3925 : OAI222_X1 port map( A1 => n7770, A2 => n14157, B1 => n1688, B2 => 
                           n14154, C1 => n7771, C2 => n14151, ZN => n3236);
   U3926 : OAI222_X1 port map( A1 => n7766, A2 => n14157, B1 => n1687, B2 => 
                           n14154, C1 => n7767, C2 => n14151, ZN => n3273);
   U3927 : OAI222_X1 port map( A1 => n7762, A2 => n14157, B1 => n1686, B2 => 
                           n14154, C1 => n7763, C2 => n14151, ZN => n3310);
   U3928 : OAI222_X1 port map( A1 => n7758, A2 => n14157, B1 => n1685, B2 => 
                           n14154, C1 => n7759, C2 => n14151, ZN => n3349);
   U3929 : OAI222_X1 port map( A1 => n7754, A2 => n14157, B1 => n1684, B2 => 
                           n14154, C1 => n7755, C2 => n14151, ZN => n3386);
   U3930 : OAI222_X1 port map( A1 => n7750, A2 => n14157, B1 => n1683, B2 => 
                           n14154, C1 => n7751, C2 => n14151, ZN => n3423);
   U3931 : OAI222_X1 port map( A1 => n7746, A2 => n14157, B1 => n1682, B2 => 
                           n14154, C1 => n7747, C2 => n14151, ZN => n3460);
   U3932 : OAI222_X1 port map( A1 => n7742, A2 => n14157, B1 => n1681, B2 => 
                           n14154, C1 => n7743, C2 => n14151, ZN => n3497);
   U3933 : OAI222_X1 port map( A1 => n7734, A2 => n14157, B1 => n1679, B2 => 
                           n14154, C1 => n7735, C2 => n14151, ZN => n3571);
   U3934 : OAI222_X1 port map( A1 => n7730, A2 => n14156, B1 => n1678, B2 => 
                           n14153, C1 => n7731, C2 => n14150, ZN => n3608);
   U3935 : OAI222_X1 port map( A1 => n7726, A2 => n14156, B1 => n1677, B2 => 
                           n14153, C1 => n7727, C2 => n14150, ZN => n3645);
   U3936 : OAI222_X1 port map( A1 => n7722, A2 => n14156, B1 => n1676, B2 => 
                           n14153, C1 => n7723, C2 => n14150, ZN => n3682);
   U3937 : OAI222_X1 port map( A1 => n7718, A2 => n14156, B1 => n1675, B2 => 
                           n14153, C1 => n7719, C2 => n14150, ZN => n3719);
   U3938 : OAI222_X1 port map( A1 => n7714, A2 => n14156, B1 => n1674, B2 => 
                           n14153, C1 => n7715, C2 => n14150, ZN => n3756);
   U3939 : OAI222_X1 port map( A1 => n7710, A2 => n14156, B1 => n1673, B2 => 
                           n14153, C1 => n7711, C2 => n14150, ZN => n3793);
   U3940 : OAI222_X1 port map( A1 => n7706, A2 => n14156, B1 => n1672, B2 => 
                           n14153, C1 => n7707, C2 => n14150, ZN => n3830);
   U3941 : OAI222_X1 port map( A1 => n7702, A2 => n14156, B1 => n1711, B2 => 
                           n14153, C1 => n7703, C2 => n14150, ZN => n3867);
   U3942 : OAI222_X1 port map( A1 => n7698, A2 => n14156, B1 => n1606, B2 => 
                           n14153, C1 => n7699, C2 => n14150, ZN => n3904);
   U3943 : OAI222_X1 port map( A1 => n7694, A2 => n14156, B1 => n1605, B2 => 
                           n14153, C1 => n7695, C2 => n14150, ZN => n3941);
   U3944 : OAI222_X1 port map( A1 => n7690, A2 => n14156, B1 => n1671, B2 => 
                           n14153, C1 => n7691, C2 => n14150, ZN => n5263);
   U3945 : AOI221_X1 port map( B1 => n13801, B2 => n8321, C1 => n13798, C2 => 
                           n8289, A => n5315, ZN => n5312);
   U3946 : OAI222_X1 port map( A1 => n1782, A2 => n13795, B1 => n6740, B2 => 
                           n13792, C1 => n1783, C2 => n13789, ZN => n5315);
   U3947 : AOI221_X1 port map( B1 => n13855, B2 => n8124, C1 => n13852, C2 => 
                           n8092, A => n5618, ZN => n5617);
   U3948 : OAI222_X1 port map( A1 => n6912, A2 => n13849, B1 => n6914, B2 => 
                           n13846, C1 => n405, C2 => n13843, ZN => n5618);
   U3949 : AOI221_X1 port map( B1 => n13801, B2 => n8314, C1 => n13798, C2 => 
                           n8282, A => n5626, ZN => n5625);
   U3950 : OAI222_X1 port map( A1 => n6906, A2 => n13795, B1 => n6908, B2 => 
                           n13792, C1 => n229, C2 => n13789, ZN => n5626);
   U3951 : AOI221_X1 port map( B1 => n7051, B2 => n14730, C1 => n883, C2 => 
                           n14725, A => n3764, ZN => n3763);
   U3952 : OAI222_X1 port map( A1 => n14117, A2 => n610, B1 => n7534, B2 => 
                           n14307, C1 => n14296, C2 => n586, ZN => n3764);
   U3953 : AOI221_X1 port map( B1 => n13966, B2 => n8615, C1 => n13964, C2 => 
                           n8583, A => n4942, ZN => n4941);
   U3954 : OAI222_X1 port map( A1 => n2074, A2 => n13961, B1 => n7310, B2 => 
                           n13956, C1 => n2088, C2 => n13955, ZN => n4942);
   U3955 : AOI221_X1 port map( B1 => n13967, B2 => n8614, C1 => n13964, C2 => 
                           n8582, A => n4979, ZN => n4978);
   U3956 : OAI222_X1 port map( A1 => n2073, A2 => n13961, B1 => n7334, B2 => 
                           n13956, C1 => n2087, C2 => n13955, ZN => n4979);
   U3957 : AOI221_X1 port map( B1 => n13967, B2 => n8613, C1 => n13964, C2 => 
                           n8581, A => n5016, ZN => n5015);
   U3958 : OAI222_X1 port map( A1 => n2072, A2 => n13961, B1 => n7358, B2 => 
                           n13956, C1 => n2086, C2 => n13955, ZN => n5016);
   U3959 : AOI221_X1 port map( B1 => n13967, B2 => n8612, C1 => n13964, C2 => 
                           n8580, A => n5053, ZN => n5052);
   U3960 : OAI222_X1 port map( A1 => n2071, A2 => n13961, B1 => n7382, B2 => 
                           n13956, C1 => n2085, C2 => n13955, ZN => n5053);
   U3961 : AOI221_X1 port map( B1 => n13967, B2 => n8611, C1 => n13964, C2 => 
                           n8579, A => n5090, ZN => n5089);
   U3962 : OAI222_X1 port map( A1 => n2070, A2 => n13961, B1 => n7406, B2 => 
                           n13956, C1 => n2084, C2 => n13955, ZN => n5090);
   U3963 : AOI221_X1 port map( B1 => n13967, B2 => n8610, C1 => n13964, C2 => 
                           n8578, A => n5127, ZN => n5126);
   U3964 : OAI222_X1 port map( A1 => n2069, A2 => n13961, B1 => n7430, B2 => 
                           n13956, C1 => n2083, C2 => n13955, ZN => n5127);
   U3965 : OAI222_X1 port map( A1 => n928, A2 => n14040, B1 => n743, B2 => 
                           n14037, C1 => n519, C2 => n14034, ZN => n4780);
   U3966 : OAI222_X1 port map( A1 => n928, A2 => n13820, B1 => n743, B2 => 
                           n13817, C1 => n519, C2 => n13814, ZN => n6101);
   U3967 : OAI222_X1 port map( A1 => n930, A2 => n14041, B1 => n807, B2 => 
                           n14038, C1 => n520, C2 => n14035, ZN => n4743);
   U3968 : OAI222_X1 port map( A1 => n930, A2 => n13821, B1 => n807, B2 => 
                           n13818, C1 => n520, C2 => n13815, ZN => n6064);
   U3969 : AOI221_X1 port map( B1 => n13938, B2 => n8443, C1 => n13935, C2 => 
                           n8411, A => n4278, ZN => n4273);
   U3970 : OAI222_X1 port map( A1 => n1752, A2 => n13932, B1 => n6881, B2 => 
                           n13931, C1 => n190, C2 => n13926, ZN => n4278);
   U3971 : AOI221_X1 port map( B1 => n13897, B2 => n8747, C1 => n13894, C2 => 
                           n8715, A => n4804, ZN => n4799);
   U3972 : OAI222_X1 port map( A1 => n2021, A2 => n13891, B1 => n2054, B2 => 
                           n13887, C1 => n2040, C2 => n13885, ZN => n4804);
   U3973 : AOI221_X1 port map( B1 => n13897, B2 => n8746, C1 => n13894, C2 => 
                           n8714, A => n4841, ZN => n4836);
   U3974 : OAI222_X1 port map( A1 => n2020, A2 => n13891, B1 => n2053, B2 => 
                           n13887, C1 => n2039, C2 => n13885, ZN => n4841);
   U3975 : AOI221_X1 port map( B1 => n13897, B2 => n8745, C1 => n13894, C2 => 
                           n8713, A => n4878, ZN => n4873);
   U3976 : OAI222_X1 port map( A1 => n2019, A2 => n13891, B1 => n7259, B2 => 
                           n13887, C1 => n2038, C2 => n13885, ZN => n4878);
   U3977 : AOI221_X1 port map( B1 => n13897, B2 => n8744, C1 => n13894, C2 => 
                           n8712, A => n4915, ZN => n4910);
   U3978 : OAI222_X1 port map( A1 => n2018, A2 => n13891, B1 => n7283, B2 => 
                           n13887, C1 => n2037, C2 => n13885, ZN => n4915);
   U3979 : AOI221_X1 port map( B1 => n13799, B2 => n8301, C1 => n13796, C2 => 
                           n8269, A => n6107, ZN => n6106);
   U3980 : OAI222_X1 port map( A1 => n2362, A2 => n13793, B1 => n2390, B2 => 
                           n13790, C1 => n2376, C2 => n13787, ZN => n6107);
   U3981 : AOI221_X1 port map( B1 => n13799, B2 => n8300, C1 => n13796, C2 => 
                           n8268, A => n6144, ZN => n6143);
   U3982 : OAI222_X1 port map( A1 => n2361, A2 => n13793, B1 => n7244, B2 => 
                           n13790, C1 => n2375, C2 => n13787, ZN => n6144);
   U3983 : AOI221_X1 port map( B1 => n13799, B2 => n8299, C1 => n13796, C2 => 
                           n8267, A => n6181, ZN => n6180);
   U3984 : OAI222_X1 port map( A1 => n2360, A2 => n13793, B1 => n7268, B2 => 
                           n13790, C1 => n2374, C2 => n13787, ZN => n6181);
   U3985 : AOI221_X1 port map( B1 => n13799, B2 => n8298, C1 => n13796, C2 => 
                           n8266, A => n6218, ZN => n6217);
   U3986 : OAI222_X1 port map( A1 => n2359, A2 => n13793, B1 => n7292, B2 => 
                           n13790, C1 => n2373, C2 => n13787, ZN => n6218);
   U3987 : AOI221_X1 port map( B1 => n13799, B2 => n8297, C1 => n13796, C2 => 
                           n8265, A => n6255, ZN => n6254);
   U3988 : OAI222_X1 port map( A1 => n2358, A2 => n13793, B1 => n7316, B2 => 
                           n13790, C1 => n2372, C2 => n13787, ZN => n6255);
   U3989 : AOI221_X1 port map( B1 => n13799, B2 => n8296, C1 => n13796, C2 => 
                           n8264, A => n6292, ZN => n6291);
   U3990 : OAI222_X1 port map( A1 => n2357, A2 => n13793, B1 => n7340, B2 => 
                           n13790, C1 => n2371, C2 => n13787, ZN => n6292);
   U3991 : AOI221_X1 port map( B1 => n13799, B2 => n8295, C1 => n13796, C2 => 
                           n8263, A => n6329, ZN => n6328);
   U3992 : OAI222_X1 port map( A1 => n2356, A2 => n13793, B1 => n7364, B2 => 
                           n13790, C1 => n2370, C2 => n13787, ZN => n6329);
   U3993 : AOI221_X1 port map( B1 => n13799, B2 => n8294, C1 => n13796, C2 => 
                           n8262, A => n6366, ZN => n6365);
   U3994 : OAI222_X1 port map( A1 => n2355, A2 => n13793, B1 => n7388, B2 => 
                           n13790, C1 => n2369, C2 => n13787, ZN => n6366);
   U3995 : AOI221_X1 port map( B1 => n13799, B2 => n8293, C1 => n13796, C2 => 
                           n8261, A => n6403, ZN => n6402);
   U3996 : OAI222_X1 port map( A1 => n2354, A2 => n13793, B1 => n7412, B2 => 
                           n13790, C1 => n2368, C2 => n13787, ZN => n6403);
   U3997 : AOI221_X1 port map( B1 => n13799, B2 => n8292, C1 => n13796, C2 => 
                           n8260, A => n6440, ZN => n6439);
   U3998 : OAI222_X1 port map( A1 => n2353, A2 => n13793, B1 => n7436, B2 => 
                           n13790, C1 => n2367, C2 => n13787, ZN => n6440);
   U3999 : AOI221_X1 port map( B1 => n13799, B2 => n8291, C1 => n13796, C2 => 
                           n8259, A => n6477, ZN => n6476);
   U4000 : OAI222_X1 port map( A1 => n2352, A2 => n13793, B1 => n7460, B2 => 
                           n13790, C1 => n2366, C2 => n13787, ZN => n6477);
   U4001 : AOI221_X1 port map( B1 => n14020, B2 => n8303, C1 => n14017, C2 => 
                           n8271, A => n4712, ZN => n4711);
   U4002 : OAI222_X1 port map( A1 => n2364, A2 => n14014, B1 => n7172, B2 => 
                           n14011, C1 => n2378, C2 => n14008, ZN => n4712);
   U4003 : AOI221_X1 port map( B1 => n13939, B2 => n8431, C1 => n13936, C2 => 
                           n8399, A => n4722, ZN => n4717);
   U4004 : OAI222_X1 port map( A1 => n2132, A2 => n13933, B1 => n7169, B2 => 
                           n13930, C1 => n2279, C2 => n13927, ZN => n4722);
   U4005 : AOI221_X1 port map( B1 => n14020, B2 => n8302, C1 => n14017, C2 => 
                           n8270, A => n4749, ZN => n4748);
   U4006 : OAI222_X1 port map( A1 => n2363, A2 => n14014, B1 => n7196, B2 => 
                           n14011, C1 => n2377, C2 => n14008, ZN => n4749);
   U4007 : AOI221_X1 port map( B1 => n13939, B2 => n8430, C1 => n13936, C2 => 
                           n8398, A => n4759, ZN => n4754);
   U4008 : OAI222_X1 port map( A1 => n2131, A2 => n13933, B1 => n7193, B2 => 
                           n13930, C1 => n2278, C2 => n13927, ZN => n4759);
   U4009 : AOI221_X1 port map( B1 => n13940, B2 => n8419, C1 => n13935, C2 => 
                           n8387, A => n5166, ZN => n5161);
   U4010 : OAI222_X1 port map( A1 => n2120, A2 => n13932, B1 => n7457, B2 => 
                           n13929, C1 => n2139, C2 => n13926, ZN => n5166);
   U4011 : AOI221_X1 port map( B1 => n13938, B2 => n8448, C1 => n13935, C2 => 
                           n8416, A => n4091, ZN => n4086);
   U4012 : OAI222_X1 port map( A1 => n1756, A2 => n13932, B1 => n6761, B2 => 
                           n13931, C1 => n195, C2 => n13926, ZN => n4091);
   U4013 : AOI221_X1 port map( B1 => n13938, B2 => n8447, C1 => n13935, C2 => 
                           n8415, A => n4130, ZN => n4125);
   U4014 : OAI222_X1 port map( A1 => n188, A2 => n13932, B1 => n6785, B2 => 
                           n13931, C1 => n194, C2 => n13926, ZN => n4130);
   U4015 : AOI221_X1 port map( B1 => n13938, B2 => n8446, C1 => n13935, C2 => 
                           n8414, A => n4167, ZN => n4162);
   U4016 : OAI222_X1 port map( A1 => n1755, A2 => n13932, B1 => n6809, B2 => 
                           n13931, C1 => n193, C2 => n13926, ZN => n4167);
   U4017 : AOI221_X1 port map( B1 => n13938, B2 => n8445, C1 => n13935, C2 => 
                           n8413, A => n4204, ZN => n4199);
   U4018 : OAI222_X1 port map( A1 => n1754, A2 => n13932, B1 => n6833, B2 => 
                           n13931, C1 => n192, C2 => n13926, ZN => n4204);
   U4019 : AOI221_X1 port map( B1 => n13938, B2 => n8444, C1 => n13935, C2 => 
                           n8412, A => n4241, ZN => n4236);
   U4020 : OAI222_X1 port map( A1 => n1753, A2 => n13932, B1 => n6857, B2 => 
                           n13931, C1 => n191, C2 => n13926, ZN => n4241);
   U4021 : AOI221_X1 port map( B1 => n13938, B2 => n8442, C1 => n13935, C2 => 
                           n8410, A => n4315, ZN => n4310);
   U4022 : OAI222_X1 port map( A1 => n1751, A2 => n13932, B1 => n6905, B2 => 
                           n13931, C1 => n189, C2 => n13926, ZN => n4315);
   U4023 : AOI221_X1 port map( B1 => n14020, B2 => n8313, C1 => n14017, C2 => 
                           n8281, A => n4342, ZN => n4341);
   U4024 : OAI222_X1 port map( A1 => n6930, A2 => n14014, B1 => n6932, B2 => 
                           n14011, C1 => n1574, C2 => n14008, ZN => n4342);
   U4025 : AOI221_X1 port map( B1 => n13939, B2 => n8441, C1 => n13936, C2 => 
                           n8409, A => n4352, ZN => n4347);
   U4026 : OAI222_X1 port map( A1 => n2137, A2 => n13933, B1 => n6929, B2 => 
                           n13930, C1 => n1462, C2 => n13927, ZN => n4352);
   U4027 : AOI221_X1 port map( B1 => n13854, B2 => n8123, C1 => n13851, C2 => 
                           n8091, A => n5655, ZN => n5654);
   U4028 : OAI222_X1 port map( A1 => n6936, A2 => n13848, B1 => n6938, B2 => 
                           n13845, C1 => n1706, C2 => n13842, ZN => n5655);
   U4029 : AOI221_X1 port map( B1 => n13938, B2 => n8440, C1 => n13935, C2 => 
                           n8408, A => n4389, ZN => n4384);
   U4030 : OAI222_X1 port map( A1 => n2136, A2 => n13932, B1 => n6953, B2 => 
                           n13930, C1 => n1461, C2 => n13926, ZN => n4389);
   U4031 : AOI221_X1 port map( B1 => n13854, B2 => n8122, C1 => n13851, C2 => 
                           n8090, A => n5692, ZN => n5691);
   U4032 : OAI222_X1 port map( A1 => n6960, A2 => n13848, B1 => n6962, B2 => 
                           n13845, C1 => n1705, C2 => n13842, ZN => n5692);
   U4033 : AOI221_X1 port map( B1 => n13938, B2 => n8439, C1 => n13935, C2 => 
                           n8407, A => n4426, ZN => n4421);
   U4034 : OAI222_X1 port map( A1 => n2135, A2 => n13932, B1 => n6977, B2 => 
                           n13930, C1 => n1460, C2 => n13926, ZN => n4426);
   U4035 : AOI221_X1 port map( B1 => n13854, B2 => n8121, C1 => n13851, C2 => 
                           n8089, A => n5729, ZN => n5728);
   U4036 : OAI222_X1 port map( A1 => n6984, A2 => n13848, B1 => n6986, B2 => 
                           n13845, C1 => n1704, C2 => n13842, ZN => n5729);
   U4037 : AOI221_X1 port map( B1 => n13938, B2 => n8438, C1 => n13935, C2 => 
                           n8406, A => n4463, ZN => n4458);
   U4038 : OAI222_X1 port map( A1 => n2134, A2 => n13932, B1 => n7001, B2 => 
                           n13930, C1 => n1459, C2 => n13926, ZN => n4463);
   U4039 : AOI221_X1 port map( B1 => n13854, B2 => n8120, C1 => n13851, C2 => 
                           n8088, A => n5766, ZN => n5765);
   U4040 : OAI222_X1 port map( A1 => n7008, A2 => n13848, B1 => n7010, B2 => 
                           n13845, C1 => n1703, C2 => n13842, ZN => n5766);
   U4041 : AOI221_X1 port map( B1 => n14019, B2 => n8309, C1 => n14017, C2 => 
                           n8277, A => n4490, ZN => n4489);
   U4042 : OAI222_X1 port map( A1 => n1564, A2 => n14014, B1 => n7028, B2 => 
                           n14011, C1 => n1570, C2 => n14008, ZN => n4490);
   U4043 : AOI221_X1 port map( B1 => n13938, B2 => n8437, C1 => n13936, C2 => 
                           n8405, A => n4500, ZN => n4495);
   U4044 : OAI222_X1 port map( A1 => n2133, A2 => n13933, B1 => n7025, B2 => 
                           n13930, C1 => n1458, C2 => n13927, ZN => n4500);
   U4045 : AOI221_X1 port map( B1 => n13854, B2 => n8119, C1 => n13851, C2 => 
                           n8087, A => n5803, ZN => n5802);
   U4046 : OAI222_X1 port map( A1 => n1696, A2 => n13848, B1 => n7034, B2 => 
                           n13845, C1 => n1702, C2 => n13842, ZN => n5803);
   U4047 : AOI221_X1 port map( B1 => n14019, B2 => n8308, C1 => n14017, C2 => 
                           n8276, A => n4527, ZN => n4526);
   U4048 : OAI222_X1 port map( A1 => n1563, A2 => n14014, B1 => n7052, B2 => 
                           n14011, C1 => n1569, C2 => n14008, ZN => n4527);
   U4049 : AOI221_X1 port map( B1 => n13938, B2 => n8436, C1 => n13936, C2 => 
                           n8404, A => n4537, ZN => n4532);
   U4050 : OAI222_X1 port map( A1 => n1452, A2 => n13933, B1 => n7049, B2 => 
                           n13930, C1 => n1457, C2 => n13927, ZN => n4537);
   U4051 : AOI221_X1 port map( B1 => n13854, B2 => n8118, C1 => n13851, C2 => 
                           n8086, A => n5840, ZN => n5839);
   U4052 : OAI222_X1 port map( A1 => n1695, A2 => n13848, B1 => n7058, B2 => 
                           n13845, C1 => n1701, C2 => n13842, ZN => n5840);
   U4053 : AOI221_X1 port map( B1 => n14020, B2 => n8307, C1 => n14017, C2 => 
                           n8275, A => n4564, ZN => n4563);
   U4054 : OAI222_X1 port map( A1 => n1562, A2 => n14014, B1 => n7076, B2 => 
                           n14011, C1 => n1568, C2 => n14008, ZN => n4564);
   U4055 : AOI221_X1 port map( B1 => n13939, B2 => n8435, C1 => n13936, C2 => 
                           n8403, A => n4574, ZN => n4569);
   U4056 : OAI222_X1 port map( A1 => n1451, A2 => n13933, B1 => n7073, B2 => 
                           n13930, C1 => n1456, C2 => n13927, ZN => n4574);
   U4057 : AOI221_X1 port map( B1 => n13854, B2 => n8117, C1 => n13851, C2 => 
                           n8085, A => n5877, ZN => n5876);
   U4058 : OAI222_X1 port map( A1 => n1694, A2 => n13848, B1 => n7082, B2 => 
                           n13845, C1 => n1700, C2 => n13842, ZN => n5877);
   U4059 : AOI221_X1 port map( B1 => n14020, B2 => n8306, C1 => n14017, C2 => 
                           n8274, A => n4601, ZN => n4600);
   U4060 : OAI222_X1 port map( A1 => n1561, A2 => n14014, B1 => n7100, B2 => 
                           n14011, C1 => n1567, C2 => n14008, ZN => n4601);
   U4061 : AOI221_X1 port map( B1 => n13939, B2 => n8434, C1 => n13936, C2 => 
                           n8402, A => n4611, ZN => n4606);
   U4062 : OAI222_X1 port map( A1 => n1450, A2 => n13933, B1 => n7097, B2 => 
                           n13930, C1 => n1455, C2 => n13927, ZN => n4611);
   U4063 : AOI221_X1 port map( B1 => n13854, B2 => n8116, C1 => n13851, C2 => 
                           n8084, A => n5914, ZN => n5913);
   U4064 : OAI222_X1 port map( A1 => n1693, A2 => n13848, B1 => n7106, B2 => 
                           n13845, C1 => n1699, C2 => n13842, ZN => n5914);
   U4065 : AOI221_X1 port map( B1 => n14020, B2 => n8305, C1 => n14017, C2 => 
                           n8273, A => n4638, ZN => n4637);
   U4066 : OAI222_X1 port map( A1 => n1560, A2 => n14014, B1 => n7124, B2 => 
                           n14011, C1 => n1566, C2 => n14008, ZN => n4638);
   U4067 : AOI221_X1 port map( B1 => n13939, B2 => n8433, C1 => n13936, C2 => 
                           n8401, A => n4648, ZN => n4643);
   U4068 : OAI222_X1 port map( A1 => n1449, A2 => n13933, B1 => n7121, B2 => 
                           n13930, C1 => n1454, C2 => n13927, ZN => n4648);
   U4069 : AOI221_X1 port map( B1 => n13854, B2 => n8115, C1 => n13851, C2 => 
                           n8083, A => n5951, ZN => n5950);
   U4070 : OAI222_X1 port map( A1 => n1692, A2 => n13848, B1 => n7130, B2 => 
                           n13845, C1 => n1698, C2 => n13842, ZN => n5951);
   U4071 : AOI221_X1 port map( B1 => n14020, B2 => n8304, C1 => n14017, C2 => 
                           n8272, A => n4675, ZN => n4674);
   U4072 : OAI222_X1 port map( A1 => n7146, A2 => n14014, B1 => n7148, B2 => 
                           n14011, C1 => n1565, C2 => n14008, ZN => n4675);
   U4073 : AOI221_X1 port map( B1 => n13939, B2 => n8432, C1 => n13936, C2 => 
                           n8400, A => n4685, ZN => n4680);
   U4074 : OAI222_X1 port map( A1 => n1448, A2 => n13933, B1 => n7145, B2 => 
                           n13930, C1 => n1453, C2 => n13927, ZN => n4685);
   U4075 : AOI221_X1 port map( B1 => n13854, B2 => n8114, C1 => n13851, C2 => 
                           n8082, A => n5988, ZN => n5987);
   U4076 : OAI222_X1 port map( A1 => n7152, A2 => n13848, B1 => n7154, B2 => 
                           n13845, C1 => n1697, C2 => n13842, ZN => n5988);
   U4077 : AOI221_X1 port map( B1 => n8608, B2 => n13967, C1 => n8576, C2 => 
                           n13962, A => n5214, ZN => n5213);
   U4078 : OAI222_X1 port map( A1 => n13959, A2 => n2067, B1 => n7478, B2 => 
                           n13956, C1 => n13953, C2 => n2081, ZN => n5214);
   U4079 : AOI221_X1 port map( B1 => n8736, B2 => n13898, C1 => n8704, C2 => 
                           n13893, A => n5227, ZN => n5221);
   U4080 : OAI222_X1 port map( A1 => n13890, A2 => n2010, B1 => n7475, B2 => 
                           n13887, C1 => n13884, C2 => n2029, ZN => n5227);
   U4081 : AOI221_X1 port map( B1 => n8639, B2 => n13967, C1 => n8607, C2 => 
                           n13962, A => n4020, ZN => n4017);
   U4082 : OAI222_X1 port map( A1 => n13959, A2 => n1741, B1 => n6734, B2 => 
                           n13958, C1 => n13953, C2 => n1742, ZN => n4020);
   U4083 : AOI221_X1 port map( B1 => n8449, B2 => n13940, C1 => n8417, C2 => 
                           n13935, A => n4031, ZN => n4015);
   U4084 : OAI222_X1 port map( A1 => n13932, A2 => n1757, B1 => n6737, B2 => 
                           n13931, C1 => n13926, C2 => n1758, ZN => n4031);
   U4085 : AOI221_X1 port map( B1 => n6843, B2 => n14729, C1 => n849, C2 => 
                           n14727, A => n3133, ZN => n3132);
   U4086 : OAI222_X1 port map( A1 => n14117, A2 => n627, B1 => n7636, B2 => 
                           n14308, C1 => n14297, C2 => n603, ZN => n3133);
   U4087 : AOI221_X1 port map( B1 => n14143, B2 => n2401, C1 => n14141, C2 => 
                           n1987, A => n3164, ZN => n3159);
   U4088 : OAI222_X1 port map( A1 => n14137, A2 => n1083, B1 => n7881, B2 => 
                           n14135, C1 => n14131, C2 => n1104, ZN => n3164);
   U4089 : AOI221_X1 port map( B1 => n14143, B2 => n2400, C1 => n14141, C2 => 
                           n1986, A => n3201, ZN => n3196);
   U4090 : OAI222_X1 port map( A1 => n14137, A2 => n1082, B1 => n7878, B2 => 
                           n14135, C1 => n14131, C2 => n1103, ZN => n3201);
   U4091 : AOI221_X1 port map( B1 => n14143, B2 => n2399, C1 => n14141, C2 => 
                           n1985, A => n3238, ZN => n3233);
   U4092 : OAI222_X1 port map( A1 => n14137, A2 => n1081, B1 => n7875, B2 => 
                           n14135, C1 => n14131, C2 => n1102, ZN => n3238);
   U4093 : AOI221_X1 port map( B1 => n14143, B2 => n2398, C1 => n14141, C2 => 
                           n1984, A => n3275, ZN => n3270);
   U4094 : OAI222_X1 port map( A1 => n14137, A2 => n1080, B1 => n7872, B2 => 
                           n14135, C1 => n14131, C2 => n1101, ZN => n3275);
   U4095 : AOI221_X1 port map( B1 => n14144, B2 => n2397, C1 => n14141, C2 => 
                           n1983, A => n3314, ZN => n3307);
   U4096 : OAI222_X1 port map( A1 => n14138, A2 => n1079, B1 => n7869, B2 => 
                           n14135, C1 => n14132, C2 => n1100, ZN => n3314);
   U4097 : AOI221_X1 port map( B1 => n14144, B2 => n2396, C1 => n14141, C2 => 
                           n1982, A => n3351, ZN => n3346);
   U4098 : OAI222_X1 port map( A1 => n14138, A2 => n1078, B1 => n7866, B2 => 
                           n14135, C1 => n14132, C2 => n1099, ZN => n3351);
   U4099 : AOI221_X1 port map( B1 => n14144, B2 => n2395, C1 => n14141, C2 => 
                           n1981, A => n3388, ZN => n3383);
   U4100 : OAI222_X1 port map( A1 => n14138, A2 => n1077, B1 => n7863, B2 => 
                           n14135, C1 => n14132, C2 => n1098, ZN => n3388);
   U4101 : AOI221_X1 port map( B1 => n14144, B2 => n2394, C1 => n14141, C2 => 
                           n1980, A => n3425, ZN => n3420);
   U4102 : OAI222_X1 port map( A1 => n14138, A2 => n1076, B1 => n7860, B2 => 
                           n14135, C1 => n14132, C2 => n1097, ZN => n3425);
   U4103 : AOI221_X1 port map( B1 => n14144, B2 => n2393, C1 => n14141, C2 => 
                           n1979, A => n3462, ZN => n3457);
   U4104 : OAI222_X1 port map( A1 => n14138, A2 => n1075, B1 => n7857, B2 => 
                           n14135, C1 => n14132, C2 => n1096, ZN => n3462);
   U4105 : AOI221_X1 port map( B1 => n14144, B2 => n2392, C1 => n14141, C2 => 
                           n1978, A => n3499, ZN => n3494);
   U4106 : OAI222_X1 port map( A1 => n14138, A2 => n1074, B1 => n7854, B2 => 
                           n14135, C1 => n14132, C2 => n1095, ZN => n3499);
   U4107 : AOI221_X1 port map( B1 => n7036, B2 => n14729, C1 => n879, C2 => 
                           n14725, A => n3690, ZN => n3689);
   U4108 : OAI222_X1 port map( A1 => n14118, A2 => n612, B1 => n7546, B2 => 
                           n14308, C1 => n14297, C2 => n588, ZN => n3690);
   U4109 : AOI221_X1 port map( B1 => n7044, B2 => n14730, C1 => n881, C2 => 
                           n14725, A => n3727, ZN => n3726);
   U4110 : OAI222_X1 port map( A1 => n14118, A2 => n611, B1 => n7540, B2 => 
                           n14308, C1 => n14297, C2 => n587, ZN => n3727);
   U4111 : AOI221_X1 port map( B1 => n6754, B2 => n14728, C1 => n835, C2 => 
                           n14727, A => n2863, ZN => n2862);
   U4112 : OAI222_X1 port map( A1 => n14117, A2 => n371, B1 => n7678, B2 => 
                           n14307, C1 => n14296, C2 => n363, ZN => n2863);
   U4113 : AOI221_X1 port map( B1 => n6893, B2 => n14729, C1 => n857, C2 => 
                           n14726, A => n3281, ZN => n3280);
   U4114 : OAI222_X1 port map( A1 => n14117, A2 => n623, B1 => n7612, B2 => 
                           n14307, C1 => n14296, C2 => n599, ZN => n3281);
   U4115 : AOI221_X1 port map( B1 => n6907, B2 => n14729, C1 => n859, C2 => 
                           n14726, A => n3320, ZN => n3319);
   U4116 : OAI222_X1 port map( A1 => n14117, A2 => n622, B1 => n7606, B2 => 
                           n14308, C1 => n14297, C2 => n598, ZN => n3320);
   U4117 : AOI221_X1 port map( B1 => n6919, B2 => n14729, C1 => n861, C2 => 
                           n14726, A => n3357, ZN => n3356);
   U4118 : OAI222_X1 port map( A1 => n14117, A2 => n621, B1 => n7600, B2 => 
                           n14308, C1 => n14297, C2 => n597, ZN => n3357);
   U4119 : AOI221_X1 port map( B1 => n6937, B2 => n14729, C1 => n863, C2 => 
                           n14726, A => n3394, ZN => n3393);
   U4120 : OAI222_X1 port map( A1 => n14117, A2 => n620, B1 => n7594, B2 => 
                           n14308, C1 => n14297, C2 => n596, ZN => n3394);
   U4121 : AOI221_X1 port map( B1 => n6946, B2 => n14729, C1 => n865, C2 => 
                           n14726, A => n3431, ZN => n3430);
   U4122 : OAI222_X1 port map( A1 => n14117, A2 => n619, B1 => n7588, B2 => 
                           n14308, C1 => n14297, C2 => n595, ZN => n3431);
   U4123 : AOI221_X1 port map( B1 => n6963, B2 => n14729, C1 => n867, C2 => 
                           n14726, A => n3468, ZN => n3467);
   U4124 : OAI222_X1 port map( A1 => n14117, A2 => n618, B1 => n7582, B2 => 
                           n14308, C1 => n14297, C2 => n594, ZN => n3468);
   U4125 : AOI221_X1 port map( B1 => n6973, B2 => n14729, C1 => n869, C2 => 
                           n14726, A => n3505, ZN => n3504);
   U4126 : OAI222_X1 port map( A1 => n14117, A2 => n617, B1 => n7576, B2 => 
                           n14308, C1 => n14297, C2 => n593, ZN => n3505);
   U4127 : AOI221_X1 port map( B1 => n14728, B2 => n1000, C1 => n873, C2 => 
                           n14726, A => n3579, ZN => n3578);
   U4128 : OAI222_X1 port map( A1 => n14117, A2 => n615, B1 => n7564, B2 => 
                           n14308, C1 => n14297, C2 => n591, ZN => n3579);
   U4129 : AOI221_X1 port map( B1 => n7013, B2 => n14729, C1 => n875, C2 => 
                           n14725, A => n3616, ZN => n3615);
   U4130 : OAI222_X1 port map( A1 => n14117, A2 => n614, B1 => n7558, B2 => 
                           n14308, C1 => n14297, C2 => n590, ZN => n3616);
   U4131 : AOI221_X1 port map( B1 => n7026, B2 => n14729, C1 => n877, C2 => 
                           n14725, A => n3653, ZN => n3652);
   U4132 : OAI222_X1 port map( A1 => n14117, A2 => n613, B1 => n7552, B2 => 
                           n14308, C1 => n14297, C2 => n589, ZN => n3653);
   U4133 : AOI221_X1 port map( B1 => n7060, B2 => n14730, C1 => n885, C2 => 
                           n14725, A => n3801, ZN => n3800);
   U4134 : OAI222_X1 port map( A1 => n14118, A2 => n609, B1 => n7528, B2 => 
                           n14308, C1 => n14297, C2 => n585, ZN => n3801);
   U4135 : AOI221_X1 port map( B1 => n7068, B2 => n14730, C1 => n887, C2 => 
                           n14725, A => n3838, ZN => n3837);
   U4136 : OAI222_X1 port map( A1 => n14118, A2 => n608, B1 => n7522, B2 => 
                           n14307, C1 => n14296, C2 => n584, ZN => n3838);
   U4137 : AOI221_X1 port map( B1 => n7075, B2 => n14730, C1 => n889, C2 => 
                           n14725, A => n3875, ZN => n3874);
   U4138 : OAI222_X1 port map( A1 => n14118, A2 => n607, B1 => n7516, B2 => 
                           n14308, C1 => n14297, C2 => n583, ZN => n3875);
   U4139 : AOI221_X1 port map( B1 => n7084, B2 => n14730, C1 => n891, C2 => 
                           n14725, A => n3912, ZN => n3911);
   U4140 : OAI222_X1 port map( A1 => n14118, A2 => n606, B1 => n7510, B2 => 
                           n14307, C1 => n14296, C2 => n582, ZN => n3912);
   U4141 : AOI221_X1 port map( B1 => n7092, B2 => n14730, C1 => n893, C2 => 
                           n14725, A => n3949, ZN => n3948);
   U4142 : OAI222_X1 port map( A1 => n14118, A2 => n605, B1 => n7504, B2 => 
                           n14308, C1 => n14297, C2 => n581, ZN => n3949);
   U4143 : AOI221_X1 port map( B1 => n7099, B2 => n14730, C1 => n895, C2 => 
                           n14725, A => n5271, ZN => n5270);
   U4144 : OAI222_X1 port map( A1 => n14118, A2 => n604, B1 => n7498, B2 => 
                           n14307, C1 => n14296, C2 => n580, ZN => n5271);
   U4145 : AOI221_X1 port map( B1 => n14728, B2 => n1001, C1 => n871, C2 => 
                           n14726, A => n3542, ZN => n3541);
   U4146 : OAI222_X1 port map( A1 => n801, A2 => n14118, B1 => n14307, B2 => 
                           n1892, C1 => n802, C2 => n14297, ZN => n3542);
   U4147 : AOI221_X1 port map( B1 => n14075, B2 => n8125, C1 => n14072, C2 => 
                           n8093, A => n4260, ZN => n4259);
   U4148 : OAI222_X1 port map( A1 => n6888, A2 => n14069, B1 => n6890, B2 => 
                           n14066, C1 => n406, C2 => n14063, ZN => n4260);
   U4149 : AOI221_X1 port map( B1 => n14019, B2 => n8315, C1 => n14016, C2 => 
                           n8283, A => n4268, ZN => n4267);
   U4150 : OAI222_X1 port map( A1 => n6882, A2 => n14013, B1 => n6884, B2 => 
                           n14012, C1 => n230, C2 => n14007, ZN => n4268);
   U4151 : AOI221_X1 port map( B1 => n13965, B2 => n8633, C1 => n13962, C2 => 
                           n8601, A => n4276, ZN => n4275);
   U4152 : OAI222_X1 port map( A1 => n6876, A2 => n13959, B1 => n6878, B2 => 
                           n13958, C1 => n134, C2 => n13953, ZN => n4276);
   U4153 : AOI221_X1 port map( B1 => n13923, B2 => n8887, C1 => n13920, C2 => 
                           n8855, A => n4284, ZN => n4283);
   U4154 : OAI222_X1 port map( A1 => n6870, A2 => n13919, B1 => n6872, B2 => 
                           n13916, C1 => n2, C2 => n13913, ZN => n4284);
   U4155 : AOI221_X1 port map( B1 => n13855, B2 => n8130, C1 => n13852, C2 => 
                           n8098, A => n5396, ZN => n5395);
   U4156 : OAI222_X1 port map( A1 => n6768, A2 => n13849, B1 => n6770, B2 => 
                           n13846, C1 => n411, C2 => n13843, ZN => n5396);
   U4157 : AOI221_X1 port map( B1 => n13801, B2 => n8320, C1 => n13798, C2 => 
                           n8288, A => n5404, ZN => n5403);
   U4158 : OAI222_X1 port map( A1 => n6762, A2 => n13795, B1 => n6764, B2 => 
                           n13792, C1 => n235, C2 => n13789, ZN => n5404);
   U4159 : AOI221_X1 port map( B1 => n13747, B2 => n8638, C1 => n13744, C2 => 
                           n8606, A => n5412, ZN => n5411);
   U4160 : OAI222_X1 port map( A1 => n6756, A2 => n13741, B1 => n6758, B2 => 
                           n13738, C1 => n139, C2 => n13735, ZN => n5412);
   U4161 : AOI221_X1 port map( B1 => n13693, B2 => n8892, C1 => n13690, C2 => 
                           n8860, A => n5420, ZN => n5419);
   U4162 : OAI222_X1 port map( A1 => n6750, A2 => n13687, B1 => n6752, B2 => 
                           n13684, C1 => n7, C2 => n13681, ZN => n5420);
   U4163 : AOI221_X1 port map( B1 => n13855, B2 => n8128, C1 => n13852, C2 => 
                           n8096, A => n5470, ZN => n5469);
   U4164 : OAI222_X1 port map( A1 => n6816, A2 => n13849, B1 => n6818, B2 => 
                           n13846, C1 => n409, C2 => n13843, ZN => n5470);
   U4165 : AOI221_X1 port map( B1 => n13801, B2 => n8318, C1 => n13798, C2 => 
                           n8286, A => n5478, ZN => n5477);
   U4166 : OAI222_X1 port map( A1 => n6810, A2 => n13795, B1 => n6812, B2 => 
                           n13792, C1 => n233, C2 => n13789, ZN => n5478);
   U4167 : AOI221_X1 port map( B1 => n13747, B2 => n8636, C1 => n13744, C2 => 
                           n8604, A => n5486, ZN => n5485);
   U4168 : OAI222_X1 port map( A1 => n6804, A2 => n13741, B1 => n6806, B2 => 
                           n13738, C1 => n137, C2 => n13735, ZN => n5486);
   U4169 : AOI221_X1 port map( B1 => n13693, B2 => n8890, C1 => n13690, C2 => 
                           n8858, A => n5494, ZN => n5493);
   U4170 : OAI222_X1 port map( A1 => n6798, A2 => n13687, B1 => n6800, B2 => 
                           n13684, C1 => n5, C2 => n13681, ZN => n5494);
   U4171 : AOI221_X1 port map( B1 => n13855, B2 => n8127, C1 => n13852, C2 => 
                           n8095, A => n5507, ZN => n5506);
   U4172 : OAI222_X1 port map( A1 => n6840, A2 => n13849, B1 => n6842, B2 => 
                           n13846, C1 => n408, C2 => n13843, ZN => n5507);
   U4173 : AOI221_X1 port map( B1 => n13801, B2 => n8317, C1 => n13798, C2 => 
                           n8285, A => n5515, ZN => n5514);
   U4174 : OAI222_X1 port map( A1 => n6834, A2 => n13795, B1 => n6836, B2 => 
                           n13792, C1 => n232, C2 => n13789, ZN => n5515);
   U4175 : AOI221_X1 port map( B1 => n13747, B2 => n8635, C1 => n13744, C2 => 
                           n8603, A => n5523, ZN => n5522);
   U4176 : OAI222_X1 port map( A1 => n6828, A2 => n13741, B1 => n6830, B2 => 
                           n13738, C1 => n136, C2 => n13735, ZN => n5523);
   U4177 : AOI221_X1 port map( B1 => n13693, B2 => n8889, C1 => n13690, C2 => 
                           n8857, A => n5531, ZN => n5530);
   U4178 : OAI222_X1 port map( A1 => n6822, A2 => n13687, B1 => n6824, B2 => 
                           n13684, C1 => n4, C2 => n13681, ZN => n5531);
   U4179 : AOI221_X1 port map( B1 => n13855, B2 => n8126, C1 => n13852, C2 => 
                           n8094, A => n5544, ZN => n5543);
   U4180 : OAI222_X1 port map( A1 => n6864, A2 => n13849, B1 => n6866, B2 => 
                           n13846, C1 => n407, C2 => n13843, ZN => n5544);
   U4181 : AOI221_X1 port map( B1 => n13801, B2 => n8316, C1 => n13798, C2 => 
                           n8284, A => n5552, ZN => n5551);
   U4182 : OAI222_X1 port map( A1 => n6858, A2 => n13795, B1 => n6860, B2 => 
                           n13792, C1 => n231, C2 => n13789, ZN => n5552);
   U4183 : AOI221_X1 port map( B1 => n13747, B2 => n8634, C1 => n13744, C2 => 
                           n8602, A => n5560, ZN => n5559);
   U4184 : OAI222_X1 port map( A1 => n6852, A2 => n13741, B1 => n6854, B2 => 
                           n13738, C1 => n135, C2 => n13735, ZN => n5560);
   U4185 : AOI221_X1 port map( B1 => n13693, B2 => n8888, C1 => n13690, C2 => 
                           n8856, A => n5568, ZN => n5567);
   U4186 : OAI222_X1 port map( A1 => n6846, A2 => n13687, B1 => n6848, B2 => 
                           n13684, C1 => n3, C2 => n13681, ZN => n5568);
   U4187 : AOI221_X1 port map( B1 => n13855, B2 => n8125, C1 => n13852, C2 => 
                           n8093, A => n5581, ZN => n5580);
   U4188 : OAI222_X1 port map( A1 => n6888, A2 => n13849, B1 => n6890, B2 => 
                           n13846, C1 => n406, C2 => n13843, ZN => n5581);
   U4189 : AOI221_X1 port map( B1 => n13801, B2 => n8315, C1 => n13798, C2 => 
                           n8283, A => n5589, ZN => n5588);
   U4190 : OAI222_X1 port map( A1 => n6882, A2 => n13795, B1 => n6884, B2 => 
                           n13792, C1 => n230, C2 => n13789, ZN => n5589);
   U4191 : AOI221_X1 port map( B1 => n13747, B2 => n8633, C1 => n13744, C2 => 
                           n8601, A => n5597, ZN => n5596);
   U4192 : OAI222_X1 port map( A1 => n6876, A2 => n13741, B1 => n6878, B2 => 
                           n13738, C1 => n134, C2 => n13735, ZN => n5597);
   U4193 : AOI221_X1 port map( B1 => n13693, B2 => n8887, C1 => n13690, C2 => 
                           n8855, A => n5605, ZN => n5604);
   U4194 : OAI222_X1 port map( A1 => n6870, A2 => n13687, B1 => n6872, B2 => 
                           n13684, C1 => n2, C2 => n13681, ZN => n5605);
   U4195 : AOI221_X1 port map( B1 => n14020, B2 => n8300, C1 => n14017, C2 => 
                           n8268, A => n4823, ZN => n4822);
   U4196 : OAI222_X1 port map( A1 => n2361, A2 => n14014, B1 => n7244, B2 => 
                           n14010, C1 => n2375, C2 => n14008, ZN => n4823);
   U4197 : AOI221_X1 port map( B1 => n13966, B2 => n8618, C1 => n13963, C2 => 
                           n8586, A => n4831, ZN => n4830);
   U4198 : OAI222_X1 port map( A1 => n2077, A2 => n13960, B1 => n7238, B2 => 
                           n13956, C1 => n2091, C2 => n13954, ZN => n4831);
   U4199 : AOI221_X1 port map( B1 => n8290, B2 => n14021, C1 => n8258, C2 => 
                           n14016, A => n5204, ZN => n5203);
   U4200 : OAI222_X1 port map( A1 => n14013, A2 => n2351, B1 => n7484, B2 => 
                           n14010, C1 => n14007, C2 => n2365, ZN => n5204);
   U4201 : AOI221_X1 port map( B1 => n8862, B2 => n13925, C1 => n8830, C2 => 
                           n13920, A => n5224, ZN => n5223);
   U4202 : OAI222_X1 port map( A1 => n7470, A2 => n13917, B1 => n7472, B2 => 
                           n13914, C1 => n7471, C2 => n13911, ZN => n5224);
   U4203 : AOI221_X1 port map( B1 => n14073, B2 => n8111, C1 => n14070, C2 => 
                           n8079, A => n4778, ZN => n4777);
   U4204 : OAI222_X1 port map( A1 => n2480, A2 => n14067, B1 => n2418, B2 => 
                           n14064, C1 => n2482, C2 => n14061, ZN => n4778);
   U4205 : AOI221_X1 port map( B1 => n14020, B2 => n8301, C1 => n14017, C2 => 
                           n8269, A => n4786, ZN => n4785);
   U4206 : OAI222_X1 port map( A1 => n2362, A2 => n14014, B1 => n2390, B2 => 
                           n14010, C1 => n2376, C2 => n14008, ZN => n4786);
   U4207 : AOI221_X1 port map( B1 => n13966, B2 => n8619, C1 => n13963, C2 => 
                           n8587, A => n4794, ZN => n4793);
   U4208 : OAI222_X1 port map( A1 => n2078, A2 => n13960, B1 => n2106, B2 => 
                           n13956, C1 => n2092, C2 => n13954, ZN => n4794);
   U4209 : AOI221_X1 port map( B1 => n13924, B2 => n8873, C1 => n13921, C2 => 
                           n8841, A => n4802, ZN => n4801);
   U4210 : OAI222_X1 port map( A1 => n2506, A2 => n13917, B1 => n1929, B2 => 
                           n13914, C1 => n1915, C2 => n13911, ZN => n4802);
   U4211 : AOI221_X1 port map( B1 => n13924, B2 => n8872, C1 => n13921, C2 => 
                           n8840, A => n4839, ZN => n4838);
   U4212 : OAI222_X1 port map( A1 => n2505, A2 => n13917, B1 => n1928, B2 => 
                           n13914, C1 => n1914, C2 => n13911, ZN => n4839);
   U4213 : AOI221_X1 port map( B1 => n14020, B2 => n8299, C1 => n14017, C2 => 
                           n8267, A => n4860, ZN => n4859);
   U4214 : OAI222_X1 port map( A1 => n2360, A2 => n14014, B1 => n7268, B2 => 
                           n14010, C1 => n2374, C2 => n14008, ZN => n4860);
   U4215 : AOI221_X1 port map( B1 => n13966, B2 => n8617, C1 => n13963, C2 => 
                           n8585, A => n4868, ZN => n4867);
   U4216 : OAI222_X1 port map( A1 => n2076, A2 => n13960, B1 => n7262, B2 => 
                           n13956, C1 => n2090, C2 => n13954, ZN => n4868);
   U4217 : AOI221_X1 port map( B1 => n13924, B2 => n8871, C1 => n13921, C2 => 
                           n8839, A => n4876, ZN => n4875);
   U4218 : OAI222_X1 port map( A1 => n7254, A2 => n13917, B1 => n7256, B2 => 
                           n13914, C1 => n7255, C2 => n13911, ZN => n4876);
   U4219 : AOI221_X1 port map( B1 => n14020, B2 => n8298, C1 => n14017, C2 => 
                           n8266, A => n4897, ZN => n4896);
   U4220 : OAI222_X1 port map( A1 => n2359, A2 => n14014, B1 => n7292, B2 => 
                           n14010, C1 => n2373, C2 => n14008, ZN => n4897);
   U4221 : AOI221_X1 port map( B1 => n13966, B2 => n8616, C1 => n13963, C2 => 
                           n8584, A => n4905, ZN => n4904);
   U4222 : OAI222_X1 port map( A1 => n2075, A2 => n13960, B1 => n7286, B2 => 
                           n13956, C1 => n2089, C2 => n13954, ZN => n4905);
   U4223 : AOI221_X1 port map( B1 => n13924, B2 => n8870, C1 => n13921, C2 => 
                           n8838, A => n4913, ZN => n4912);
   U4224 : OAI222_X1 port map( A1 => n7278, A2 => n13917, B1 => n7280, B2 => 
                           n13914, C1 => n7279, C2 => n13911, ZN => n4913);
   U4225 : AOI221_X1 port map( B1 => n14019, B2 => n8316, C1 => n14016, C2 => 
                           n8284, A => n4231, ZN => n4230);
   U4226 : OAI222_X1 port map( A1 => n6858, A2 => n14013, B1 => n6860, B2 => 
                           n14012, C1 => n231, C2 => n14007, ZN => n4231);
   U4227 : AOI221_X1 port map( B1 => n13965, B2 => n8634, C1 => n13962, C2 => 
                           n8602, A => n4239, ZN => n4238);
   U4228 : OAI222_X1 port map( A1 => n6852, A2 => n13959, B1 => n6854, B2 => 
                           n13958, C1 => n135, C2 => n13953, ZN => n4239);
   U4229 : AOI221_X1 port map( B1 => n14020, B2 => n8297, C1 => n14018, C2 => 
                           n8265, A => n4934, ZN => n4933);
   U4230 : OAI222_X1 port map( A1 => n2358, A2 => n14015, B1 => n7316, B2 => 
                           n14010, C1 => n2372, C2 => n14009, ZN => n4934);
   U4231 : AOI221_X1 port map( B1 => n13924, B2 => n8869, C1 => n13922, C2 => 
                           n8837, A => n4950, ZN => n4949);
   U4232 : OAI222_X1 port map( A1 => n7302, A2 => n13917, B1 => n7304, B2 => 
                           n13914, C1 => n7303, C2 => n13911, ZN => n4950);
   U4233 : AOI221_X1 port map( B1 => n13853, B2 => n8111, C1 => n13850, C2 => 
                           n8079, A => n6099, ZN => n6098);
   U4234 : OAI222_X1 port map( A1 => n2480, A2 => n13847, B1 => n2418, B2 => 
                           n13844, C1 => n2482, C2 => n13841, ZN => n6099);
   U4235 : AOI221_X1 port map( B1 => n13745, B2 => n8619, C1 => n13742, C2 => 
                           n8587, A => n6115, ZN => n6114);
   U4236 : OAI222_X1 port map( A1 => n2078, A2 => n13739, B1 => n2106, B2 => 
                           n13736, C1 => n2092, C2 => n13733, ZN => n6115);
   U4237 : AOI221_X1 port map( B1 => n13691, B2 => n8873, C1 => n13688, C2 => 
                           n8841, A => n6123, ZN => n6122);
   U4238 : OAI222_X1 port map( A1 => n2506, A2 => n13685, B1 => n1929, B2 => 
                           n13682, C1 => n1915, C2 => n13679, ZN => n6123);
   U4239 : AOI221_X1 port map( B1 => n13745, B2 => n8618, C1 => n13742, C2 => 
                           n8586, A => n6152, ZN => n6151);
   U4240 : OAI222_X1 port map( A1 => n2077, A2 => n13739, B1 => n7238, B2 => 
                           n13736, C1 => n2091, C2 => n13733, ZN => n6152);
   U4241 : AOI221_X1 port map( B1 => n13691, B2 => n8872, C1 => n13688, C2 => 
                           n8840, A => n6160, ZN => n6159);
   U4242 : OAI222_X1 port map( A1 => n2505, A2 => n13685, B1 => n1928, B2 => 
                           n13682, C1 => n1914, C2 => n13679, ZN => n6160);
   U4243 : AOI221_X1 port map( B1 => n13745, B2 => n8617, C1 => n13742, C2 => 
                           n8585, A => n6189, ZN => n6188);
   U4244 : OAI222_X1 port map( A1 => n2076, A2 => n13739, B1 => n7262, B2 => 
                           n13736, C1 => n2090, C2 => n13733, ZN => n6189);
   U4245 : AOI221_X1 port map( B1 => n13691, B2 => n8871, C1 => n13688, C2 => 
                           n8839, A => n6197, ZN => n6196);
   U4246 : OAI222_X1 port map( A1 => n7254, A2 => n13685, B1 => n7256, B2 => 
                           n13682, C1 => n7255, C2 => n13679, ZN => n6197);
   U4247 : AOI221_X1 port map( B1 => n13745, B2 => n8616, C1 => n13742, C2 => 
                           n8584, A => n6226, ZN => n6225);
   U4248 : OAI222_X1 port map( A1 => n2075, A2 => n13739, B1 => n7286, B2 => 
                           n13736, C1 => n2089, C2 => n13733, ZN => n6226);
   U4249 : AOI221_X1 port map( B1 => n13691, B2 => n8870, C1 => n13688, C2 => 
                           n8838, A => n6234, ZN => n6233);
   U4250 : OAI222_X1 port map( A1 => n7278, A2 => n13685, B1 => n7280, B2 => 
                           n13682, C1 => n7279, C2 => n13679, ZN => n6234);
   U4251 : AOI221_X1 port map( B1 => n13745, B2 => n8615, C1 => n13742, C2 => 
                           n8583, A => n6263, ZN => n6262);
   U4252 : OAI222_X1 port map( A1 => n2074, A2 => n13739, B1 => n7310, B2 => 
                           n13736, C1 => n2088, C2 => n13733, ZN => n6263);
   U4253 : AOI221_X1 port map( B1 => n13691, B2 => n8869, C1 => n13688, C2 => 
                           n8837, A => n6271, ZN => n6270);
   U4254 : OAI222_X1 port map( A1 => n7302, A2 => n13685, B1 => n7304, B2 => 
                           n13682, C1 => n7303, C2 => n13679, ZN => n6271);
   U4255 : AOI221_X1 port map( B1 => n13745, B2 => n8614, C1 => n13742, C2 => 
                           n8582, A => n6300, ZN => n6299);
   U4256 : OAI222_X1 port map( A1 => n2073, A2 => n13739, B1 => n7334, B2 => 
                           n13736, C1 => n2087, C2 => n13733, ZN => n6300);
   U4257 : AOI221_X1 port map( B1 => n13691, B2 => n8868, C1 => n13688, C2 => 
                           n8836, A => n6308, ZN => n6307);
   U4258 : OAI222_X1 port map( A1 => n7326, A2 => n13685, B1 => n7328, B2 => 
                           n13682, C1 => n7327, C2 => n13679, ZN => n6308);
   U4259 : AOI221_X1 port map( B1 => n13745, B2 => n8613, C1 => n13742, C2 => 
                           n8581, A => n6337, ZN => n6336);
   U4260 : OAI222_X1 port map( A1 => n2072, A2 => n13739, B1 => n7358, B2 => 
                           n13736, C1 => n2086, C2 => n13733, ZN => n6337);
   U4261 : AOI221_X1 port map( B1 => n13691, B2 => n8867, C1 => n13688, C2 => 
                           n8835, A => n6345, ZN => n6344);
   U4262 : OAI222_X1 port map( A1 => n7350, A2 => n13685, B1 => n7352, B2 => 
                           n13682, C1 => n7351, C2 => n13679, ZN => n6345);
   U4263 : AOI221_X1 port map( B1 => n13745, B2 => n8612, C1 => n13742, C2 => 
                           n8580, A => n6374, ZN => n6373);
   U4264 : OAI222_X1 port map( A1 => n2071, A2 => n13739, B1 => n7382, B2 => 
                           n13736, C1 => n2085, C2 => n13733, ZN => n6374);
   U4265 : AOI221_X1 port map( B1 => n13691, B2 => n8866, C1 => n13688, C2 => 
                           n8834, A => n6382, ZN => n6381);
   U4266 : OAI222_X1 port map( A1 => n7374, A2 => n13685, B1 => n7376, B2 => 
                           n13682, C1 => n7375, C2 => n13679, ZN => n6382);
   U4267 : AOI221_X1 port map( B1 => n13745, B2 => n8611, C1 => n13742, C2 => 
                           n8579, A => n6411, ZN => n6410);
   U4268 : OAI222_X1 port map( A1 => n2070, A2 => n13739, B1 => n7406, B2 => 
                           n13736, C1 => n2084, C2 => n13733, ZN => n6411);
   U4269 : AOI221_X1 port map( B1 => n13691, B2 => n8865, C1 => n13688, C2 => 
                           n8833, A => n6419, ZN => n6418);
   U4270 : OAI222_X1 port map( A1 => n7398, A2 => n13685, B1 => n7400, B2 => 
                           n13682, C1 => n7399, C2 => n13679, ZN => n6419);
   U4271 : AOI221_X1 port map( B1 => n13745, B2 => n8610, C1 => n13742, C2 => 
                           n8578, A => n6448, ZN => n6447);
   U4272 : OAI222_X1 port map( A1 => n2069, A2 => n13739, B1 => n7430, B2 => 
                           n13736, C1 => n2083, C2 => n13733, ZN => n6448);
   U4273 : AOI221_X1 port map( B1 => n13691, B2 => n8864, C1 => n13688, C2 => 
                           n8832, A => n6456, ZN => n6455);
   U4274 : OAI222_X1 port map( A1 => n7422, A2 => n13685, B1 => n7424, B2 => 
                           n13682, C1 => n7423, C2 => n13679, ZN => n6456);
   U4275 : AOI221_X1 port map( B1 => n13745, B2 => n8609, C1 => n13742, C2 => 
                           n8577, A => n6485, ZN => n6484);
   U4276 : OAI222_X1 port map( A1 => n2068, A2 => n13739, B1 => n7454, B2 => 
                           n13736, C1 => n2082, C2 => n13733, ZN => n6485);
   U4277 : AOI221_X1 port map( B1 => n13691, B2 => n8863, C1 => n13688, C2 => 
                           n8831, A => n6493, ZN => n6492);
   U4278 : OAI222_X1 port map( A1 => n7446, A2 => n13685, B1 => n7448, B2 => 
                           n13682, C1 => n7447, C2 => n13679, ZN => n6493);
   U4279 : AOI221_X1 port map( B1 => n13966, B2 => n8621, C1 => n13963, C2 => 
                           n8589, A => n4720, ZN => n4719);
   U4280 : OAI222_X1 port map( A1 => n2080, A2 => n13960, B1 => n7166, B2 => 
                           n13957, C1 => n2094, C2 => n13954, ZN => n4720);
   U4281 : AOI221_X1 port map( B1 => n13924, B2 => n8875, C1 => n13921, C2 => 
                           n8843, A => n4728, ZN => n4727);
   U4282 : OAI222_X1 port map( A1 => n7158, A2 => n13918, B1 => n7160, B2 => 
                           n13915, C1 => n7159, C2 => n13912, ZN => n4728);
   U4283 : AOI221_X1 port map( B1 => n13966, B2 => n8620, C1 => n13963, C2 => 
                           n8588, A => n4757, ZN => n4756);
   U4284 : OAI222_X1 port map( A1 => n2079, A2 => n13960, B1 => n7190, B2 => 
                           n13957, C1 => n2093, C2 => n13954, ZN => n4757);
   U4285 : AOI221_X1 port map( B1 => n13924, B2 => n8874, C1 => n13921, C2 => 
                           n8842, A => n4765, ZN => n4764);
   U4286 : OAI222_X1 port map( A1 => n7182, A2 => n13918, B1 => n7184, B2 => 
                           n13915, C1 => n7183, C2 => n13912, ZN => n4765);
   U4287 : AOI221_X1 port map( B1 => n13800, B2 => n8303, C1 => n13797, C2 => 
                           n8271, A => n6033, ZN => n6032);
   U4288 : OAI222_X1 port map( A1 => n2364, A2 => n13794, B1 => n7172, B2 => 
                           n13791, C1 => n2378, C2 => n13788, ZN => n6033);
   U4289 : AOI221_X1 port map( B1 => n13746, B2 => n8621, C1 => n13743, C2 => 
                           n8589, A => n6041, ZN => n6040);
   U4290 : OAI222_X1 port map( A1 => n2080, A2 => n13740, B1 => n7166, B2 => 
                           n13737, C1 => n2094, C2 => n13734, ZN => n6041);
   U4291 : AOI221_X1 port map( B1 => n13692, B2 => n8875, C1 => n13689, C2 => 
                           n8843, A => n6049, ZN => n6048);
   U4292 : OAI222_X1 port map( A1 => n7158, A2 => n13686, B1 => n7160, B2 => 
                           n13683, C1 => n7159, C2 => n13680, ZN => n6049);
   U4293 : AOI221_X1 port map( B1 => n13800, B2 => n8302, C1 => n13797, C2 => 
                           n8270, A => n6070, ZN => n6069);
   U4294 : OAI222_X1 port map( A1 => n2363, A2 => n13794, B1 => n7196, B2 => 
                           n13791, C1 => n2377, C2 => n13788, ZN => n6070);
   U4295 : AOI221_X1 port map( B1 => n13746, B2 => n8620, C1 => n13743, C2 => 
                           n8588, A => n6078, ZN => n6077);
   U4296 : OAI222_X1 port map( A1 => n2079, A2 => n13740, B1 => n7190, B2 => 
                           n13737, C1 => n2093, C2 => n13734, ZN => n6078);
   U4297 : AOI221_X1 port map( B1 => n13692, B2 => n8874, C1 => n13689, C2 => 
                           n8842, A => n6086, ZN => n6085);
   U4298 : OAI222_X1 port map( A1 => n7182, A2 => n13686, B1 => n7184, B2 => 
                           n13683, C1 => n7183, C2 => n13680, ZN => n6086);
   U4299 : AOI221_X1 port map( B1 => n13799, B2 => n8290, C1 => n13796, C2 => 
                           n8258, A => n6525, ZN => n6524);
   U4300 : OAI222_X1 port map( A1 => n2351, A2 => n13793, B1 => n7484, B2 => 
                           n13790, C1 => n2365, C2 => n13787, ZN => n6525);
   U4301 : AOI221_X1 port map( B1 => n13745, B2 => n8608, C1 => n13742, C2 => 
                           n8576, A => n6535, ZN => n6534);
   U4302 : OAI222_X1 port map( A1 => n2067, A2 => n13739, B1 => n7478, B2 => 
                           n13736, C1 => n2081, C2 => n13733, ZN => n6535);
   U4303 : AOI221_X1 port map( B1 => n13691, B2 => n8862, C1 => n13688, C2 => 
                           n8830, A => n6545, ZN => n6544);
   U4304 : OAI222_X1 port map( A1 => n7470, A2 => n13685, B1 => n7472, B2 => 
                           n13682, C1 => n7471, C2 => n13679, ZN => n6545);
   U4305 : AOI221_X1 port map( B1 => n14021, B2 => n8296, C1 => n14018, C2 => 
                           n8264, A => n4971, ZN => n4970);
   U4306 : OAI222_X1 port map( A1 => n2357, A2 => n14015, B1 => n7340, B2 => 
                           n14010, C1 => n2371, C2 => n14009, ZN => n4971);
   U4307 : AOI221_X1 port map( B1 => n13925, B2 => n8868, C1 => n13922, C2 => 
                           n8836, A => n4987, ZN => n4986);
   U4308 : OAI222_X1 port map( A1 => n7326, A2 => n13917, B1 => n7328, B2 => 
                           n13914, C1 => n7327, C2 => n13911, ZN => n4987);
   U4309 : AOI221_X1 port map( B1 => n14021, B2 => n8295, C1 => n14018, C2 => 
                           n8263, A => n5008, ZN => n5007);
   U4310 : OAI222_X1 port map( A1 => n2356, A2 => n14015, B1 => n7364, B2 => 
                           n14010, C1 => n2370, C2 => n14009, ZN => n5008);
   U4311 : AOI221_X1 port map( B1 => n13925, B2 => n8867, C1 => n13922, C2 => 
                           n8835, A => n5024, ZN => n5023);
   U4312 : OAI222_X1 port map( A1 => n7350, A2 => n13917, B1 => n7352, B2 => 
                           n13914, C1 => n7351, C2 => n13911, ZN => n5024);
   U4313 : AOI221_X1 port map( B1 => n14021, B2 => n8294, C1 => n14018, C2 => 
                           n8262, A => n5045, ZN => n5044);
   U4314 : OAI222_X1 port map( A1 => n2355, A2 => n14015, B1 => n7388, B2 => 
                           n14010, C1 => n2369, C2 => n14009, ZN => n5045);
   U4315 : AOI221_X1 port map( B1 => n13925, B2 => n8866, C1 => n13922, C2 => 
                           n8834, A => n5061, ZN => n5060);
   U4316 : OAI222_X1 port map( A1 => n7374, A2 => n13917, B1 => n7376, B2 => 
                           n13914, C1 => n7375, C2 => n13911, ZN => n5061);
   U4317 : AOI221_X1 port map( B1 => n13925, B2 => n8865, C1 => n13922, C2 => 
                           n8833, A => n5098, ZN => n5097);
   U4318 : OAI222_X1 port map( A1 => n7398, A2 => n13917, B1 => n7400, B2 => 
                           n13914, C1 => n7399, C2 => n13911, ZN => n5098);
   U4319 : AOI221_X1 port map( B1 => n13925, B2 => n8864, C1 => n13922, C2 => 
                           n8832, A => n5135, ZN => n5134);
   U4320 : OAI222_X1 port map( A1 => n7422, A2 => n13917, B1 => n7424, B2 => 
                           n13914, C1 => n7423, C2 => n13911, ZN => n5135);
   U4321 : AOI221_X1 port map( B1 => n14021, B2 => n8291, C1 => n14016, C2 => 
                           n8259, A => n5156, ZN => n5155);
   U4322 : OAI222_X1 port map( A1 => n2352, A2 => n14013, B1 => n7460, B2 => 
                           n14010, C1 => n2366, C2 => n14007, ZN => n5156);
   U4323 : AOI221_X1 port map( B1 => n13967, B2 => n8609, C1 => n13962, C2 => 
                           n8577, A => n5164, ZN => n5163);
   U4324 : OAI222_X1 port map( A1 => n2068, A2 => n13959, B1 => n7454, B2 => 
                           n13956, C1 => n2082, C2 => n13953, ZN => n5164);
   U4325 : AOI221_X1 port map( B1 => n14021, B2 => n8293, C1 => n14018, C2 => 
                           n8261, A => n5082, ZN => n5081);
   U4326 : OAI222_X1 port map( A1 => n2354, A2 => n14015, B1 => n7412, B2 => 
                           n14010, C1 => n2368, C2 => n14009, ZN => n5082);
   U4327 : AOI221_X1 port map( B1 => n14021, B2 => n8292, C1 => n14018, C2 => 
                           n8260, A => n5119, ZN => n5118);
   U4328 : OAI222_X1 port map( A1 => n2353, A2 => n14015, B1 => n7436, B2 => 
                           n14010, C1 => n2367, C2 => n14009, ZN => n5119);
   U4329 : AOI221_X1 port map( B1 => n13925, B2 => n8863, C1 => n13920, C2 => 
                           n8831, A => n5172, ZN => n5171);
   U4330 : OAI222_X1 port map( A1 => n7446, A2 => n13917, B1 => n7448, B2 => 
                           n13914, C1 => n7447, C2 => n13911, ZN => n5172);
   U4331 : AOI221_X1 port map( B1 => n8321, B2 => n14021, C1 => n8289, C2 => 
                           n14016, A => n3994, ZN => n3991);
   U4332 : OAI222_X1 port map( A1 => n14013, A2 => n1782, B1 => n6740, B2 => 
                           n14012, C1 => n14007, C2 => n1783, ZN => n3994);
   U4333 : AOI221_X1 port map( B1 => n13747, B2 => n8639, C1 => n13744, C2 => 
                           n8607, A => n5341, ZN => n5338);
   U4334 : OAI222_X1 port map( A1 => n1741, A2 => n13741, B1 => n6734, B2 => 
                           n13738, C1 => n1742, C2 => n13735, ZN => n5341);
   U4335 : AOI221_X1 port map( B1 => n14075, B2 => n8130, C1 => n14072, C2 => 
                           n8098, A => n4073, ZN => n4072);
   U4336 : OAI222_X1 port map( A1 => n6768, A2 => n14069, B1 => n6770, B2 => 
                           n14066, C1 => n411, C2 => n14063, ZN => n4073);
   U4337 : AOI221_X1 port map( B1 => n14019, B2 => n8320, C1 => n14016, C2 => 
                           n8288, A => n4081, ZN => n4080);
   U4338 : OAI222_X1 port map( A1 => n6762, A2 => n14013, B1 => n6764, B2 => 
                           n14012, C1 => n235, C2 => n14007, ZN => n4081);
   U4339 : AOI221_X1 port map( B1 => n13965, B2 => n8638, C1 => n13962, C2 => 
                           n8606, A => n4089, ZN => n4088);
   U4340 : OAI222_X1 port map( A1 => n6756, A2 => n13959, B1 => n6758, B2 => 
                           n13958, C1 => n139, C2 => n13953, ZN => n4089);
   U4341 : AOI221_X1 port map( B1 => n13923, B2 => n8892, C1 => n13920, C2 => 
                           n8860, A => n4099, ZN => n4098);
   U4342 : OAI222_X1 port map( A1 => n6750, A2 => n13919, B1 => n6752, B2 => 
                           n13916, C1 => n7, C2 => n13913, ZN => n4099);
   U4343 : AOI221_X1 port map( B1 => n14075, B2 => n8129, C1 => n14072, C2 => 
                           n8097, A => n4112, ZN => n4111);
   U4344 : OAI222_X1 port map( A1 => n6792, A2 => n14069, B1 => n6794, B2 => 
                           n14066, C1 => n410, C2 => n14063, ZN => n4112);
   U4345 : AOI221_X1 port map( B1 => n14019, B2 => n8319, C1 => n14016, C2 => 
                           n8287, A => n4120, ZN => n4119);
   U4346 : OAI222_X1 port map( A1 => n6786, A2 => n14013, B1 => n6788, B2 => 
                           n14012, C1 => n234, C2 => n14007, ZN => n4120);
   U4347 : AOI221_X1 port map( B1 => n13965, B2 => n8637, C1 => n13962, C2 => 
                           n8605, A => n4128, ZN => n4127);
   U4348 : OAI222_X1 port map( A1 => n132, A2 => n13959, B1 => n6782, B2 => 
                           n13958, C1 => n138, C2 => n13953, ZN => n4128);
   U4349 : AOI221_X1 port map( B1 => n13923, B2 => n8891, C1 => n13920, C2 => 
                           n8859, A => n4136, ZN => n4135);
   U4350 : OAI222_X1 port map( A1 => n6774, A2 => n13919, B1 => n6776, B2 => 
                           n13916, C1 => n6, C2 => n13913, ZN => n4136);
   U4351 : AOI221_X1 port map( B1 => n13855, B2 => n8129, C1 => n13852, C2 => 
                           n8097, A => n5433, ZN => n5432);
   U4352 : OAI222_X1 port map( A1 => n6792, A2 => n13849, B1 => n6794, B2 => 
                           n13846, C1 => n410, C2 => n13843, ZN => n5433);
   U4353 : AOI221_X1 port map( B1 => n13801, B2 => n8319, C1 => n13798, C2 => 
                           n8287, A => n5441, ZN => n5440);
   U4354 : OAI222_X1 port map( A1 => n6786, A2 => n13795, B1 => n6788, B2 => 
                           n13792, C1 => n234, C2 => n13789, ZN => n5441);
   U4355 : AOI221_X1 port map( B1 => n13747, B2 => n8637, C1 => n13744, C2 => 
                           n8605, A => n5449, ZN => n5448);
   U4356 : OAI222_X1 port map( A1 => n132, A2 => n13741, B1 => n6782, B2 => 
                           n13738, C1 => n138, C2 => n13735, ZN => n5449);
   U4357 : AOI221_X1 port map( B1 => n13693, B2 => n8891, C1 => n13690, C2 => 
                           n8859, A => n5457, ZN => n5456);
   U4358 : OAI222_X1 port map( A1 => n6774, A2 => n13687, B1 => n6776, B2 => 
                           n13684, C1 => n6, C2 => n13681, ZN => n5457);
   U4359 : AOI221_X1 port map( B1 => n14019, B2 => n8318, C1 => n14016, C2 => 
                           n8286, A => n4157, ZN => n4156);
   U4360 : OAI222_X1 port map( A1 => n6810, A2 => n14013, B1 => n6812, B2 => 
                           n14012, C1 => n233, C2 => n14007, ZN => n4157);
   U4361 : AOI221_X1 port map( B1 => n13965, B2 => n8636, C1 => n13962, C2 => 
                           n8604, A => n4165, ZN => n4164);
   U4362 : OAI222_X1 port map( A1 => n6804, A2 => n13959, B1 => n6806, B2 => 
                           n13958, C1 => n137, C2 => n13953, ZN => n4165);
   U4363 : AOI221_X1 port map( B1 => n13923, B2 => n8888, C1 => n13920, C2 => 
                           n8856, A => n4247, ZN => n4246);
   U4364 : OAI222_X1 port map( A1 => n6846, A2 => n13919, B1 => n6848, B2 => 
                           n13916, C1 => n3, C2 => n13913, ZN => n4247);
   U4365 : AOI221_X1 port map( B1 => n14075, B2 => n8124, C1 => n14072, C2 => 
                           n8092, A => n4297, ZN => n4296);
   U4366 : OAI222_X1 port map( A1 => n6912, A2 => n14069, B1 => n6914, B2 => 
                           n14066, C1 => n405, C2 => n14063, ZN => n4297);
   U4367 : AOI221_X1 port map( B1 => n14019, B2 => n8314, C1 => n14016, C2 => 
                           n8282, A => n4305, ZN => n4304);
   U4368 : OAI222_X1 port map( A1 => n6906, A2 => n14013, B1 => n6908, B2 => 
                           n14012, C1 => n229, C2 => n14007, ZN => n4305);
   U4369 : AOI221_X1 port map( B1 => n13965, B2 => n8632, C1 => n13962, C2 => 
                           n8600, A => n4313, ZN => n4312);
   U4370 : OAI222_X1 port map( A1 => n6900, A2 => n13959, B1 => n6902, B2 => 
                           n13958, C1 => n133, C2 => n13953, ZN => n4313);
   U4371 : AOI221_X1 port map( B1 => n13923, B2 => n8886, C1 => n13920, C2 => 
                           n8854, A => n4321, ZN => n4320);
   U4372 : OAI222_X1 port map( A1 => n6894, A2 => n13919, B1 => n6896, B2 => 
                           n13916, C1 => n1, C2 => n13913, ZN => n4321);
   U4373 : AOI221_X1 port map( B1 => n13747, B2 => n8632, C1 => n13744, C2 => 
                           n8600, A => n5634, ZN => n5633);
   U4374 : OAI222_X1 port map( A1 => n6900, A2 => n13741, B1 => n6902, B2 => 
                           n13738, C1 => n133, C2 => n13735, ZN => n5634);
   U4375 : AOI221_X1 port map( B1 => n13693, B2 => n8886, C1 => n13690, C2 => 
                           n8854, A => n5642, ZN => n5641);
   U4376 : OAI222_X1 port map( A1 => n6894, A2 => n13687, B1 => n6896, B2 => 
                           n13684, C1 => n1, C2 => n13681, ZN => n5642);
   U4377 : AOI221_X1 port map( B1 => n14074, B2 => n8123, C1 => n14071, C2 => 
                           n8091, A => n4334, ZN => n4333);
   U4378 : OAI222_X1 port map( A1 => n6936, A2 => n14068, B1 => n6938, B2 => 
                           n14065, C1 => n1706, C2 => n14062, ZN => n4334);
   U4379 : AOI221_X1 port map( B1 => n13966, B2 => n8631, C1 => n13963, C2 => 
                           n8599, A => n4350, ZN => n4349);
   U4380 : OAI222_X1 port map( A1 => n6924, A2 => n13960, B1 => n6926, B2 => 
                           n13957, C1 => n1303, C2 => n13954, ZN => n4350);
   U4381 : AOI221_X1 port map( B1 => n13924, B2 => n8885, C1 => n13921, C2 => 
                           n8853, A => n4358, ZN => n4357);
   U4382 : OAI222_X1 port map( A1 => n6918, A2 => n13918, B1 => n6920, B2 => 
                           n13915, C1 => n637, C2 => n13912, ZN => n4358);
   U4383 : AOI221_X1 port map( B1 => n13800, B2 => n8313, C1 => n13797, C2 => 
                           n8281, A => n5663, ZN => n5662);
   U4384 : OAI222_X1 port map( A1 => n6930, A2 => n13794, B1 => n6932, B2 => 
                           n13791, C1 => n1574, C2 => n13788, ZN => n5663);
   U4385 : AOI221_X1 port map( B1 => n13746, B2 => n8631, C1 => n13743, C2 => 
                           n8599, A => n5671, ZN => n5670);
   U4386 : OAI222_X1 port map( A1 => n6924, A2 => n13740, B1 => n6926, B2 => 
                           n13737, C1 => n1303, C2 => n13734, ZN => n5671);
   U4387 : AOI221_X1 port map( B1 => n13692, B2 => n8885, C1 => n13689, C2 => 
                           n8853, A => n5679, ZN => n5678);
   U4388 : OAI222_X1 port map( A1 => n6918, A2 => n13686, B1 => n6920, B2 => 
                           n13683, C1 => n637, C2 => n13680, ZN => n5679);
   U4389 : AOI221_X1 port map( B1 => n14074, B2 => n8122, C1 => n14071, C2 => 
                           n8090, A => n4371, ZN => n4370);
   U4390 : OAI222_X1 port map( A1 => n6960, A2 => n14068, B1 => n6962, B2 => 
                           n14065, C1 => n1705, C2 => n14062, ZN => n4371);
   U4391 : AOI221_X1 port map( B1 => n14019, B2 => n8312, C1 => n14016, C2 => 
                           n8280, A => n4379, ZN => n4378);
   U4392 : OAI222_X1 port map( A1 => n6954, A2 => n14013, B1 => n6956, B2 => 
                           n14011, C1 => n1573, C2 => n14007, ZN => n4379);
   U4393 : AOI221_X1 port map( B1 => n13965, B2 => n8630, C1 => n13962, C2 => 
                           n8598, A => n4387, ZN => n4386);
   U4394 : OAI222_X1 port map( A1 => n6948, A2 => n13959, B1 => n6950, B2 => 
                           n13957, C1 => n1302, C2 => n13953, ZN => n4387);
   U4395 : AOI221_X1 port map( B1 => n13923, B2 => n8884, C1 => n13920, C2 => 
                           n8852, A => n4395, ZN => n4394);
   U4396 : OAI222_X1 port map( A1 => n6942, A2 => n13918, B1 => n6944, B2 => 
                           n13915, C1 => n636, C2 => n13912, ZN => n4395);
   U4397 : AOI221_X1 port map( B1 => n13800, B2 => n8312, C1 => n13797, C2 => 
                           n8280, A => n5700, ZN => n5699);
   U4398 : OAI222_X1 port map( A1 => n6954, A2 => n13794, B1 => n6956, B2 => 
                           n13791, C1 => n1573, C2 => n13788, ZN => n5700);
   U4399 : AOI221_X1 port map( B1 => n13746, B2 => n8630, C1 => n13743, C2 => 
                           n8598, A => n5708, ZN => n5707);
   U4400 : OAI222_X1 port map( A1 => n6948, A2 => n13740, B1 => n6950, B2 => 
                           n13737, C1 => n1302, C2 => n13734, ZN => n5708);
   U4401 : AOI221_X1 port map( B1 => n13692, B2 => n8884, C1 => n13689, C2 => 
                           n8852, A => n5716, ZN => n5715);
   U4402 : OAI222_X1 port map( A1 => n6942, A2 => n13686, B1 => n6944, B2 => 
                           n13683, C1 => n636, C2 => n13680, ZN => n5716);
   U4403 : AOI221_X1 port map( B1 => n14074, B2 => n8121, C1 => n14071, C2 => 
                           n8089, A => n4408, ZN => n4407);
   U4404 : OAI222_X1 port map( A1 => n6984, A2 => n14068, B1 => n6986, B2 => 
                           n14065, C1 => n1704, C2 => n14062, ZN => n4408);
   U4405 : AOI221_X1 port map( B1 => n14019, B2 => n8311, C1 => n14016, C2 => 
                           n8279, A => n4416, ZN => n4415);
   U4406 : OAI222_X1 port map( A1 => n6978, A2 => n14013, B1 => n6980, B2 => 
                           n14011, C1 => n1572, C2 => n14007, ZN => n4416);
   U4407 : AOI221_X1 port map( B1 => n13965, B2 => n8629, C1 => n13962, C2 => 
                           n8597, A => n4424, ZN => n4423);
   U4408 : OAI222_X1 port map( A1 => n6972, A2 => n13959, B1 => n6974, B2 => 
                           n13957, C1 => n1301, C2 => n13953, ZN => n4424);
   U4409 : AOI221_X1 port map( B1 => n13923, B2 => n8883, C1 => n13920, C2 => 
                           n8851, A => n4432, ZN => n4431);
   U4410 : OAI222_X1 port map( A1 => n6966, A2 => n13918, B1 => n6968, B2 => 
                           n13915, C1 => n635, C2 => n13912, ZN => n4432);
   U4411 : AOI221_X1 port map( B1 => n13800, B2 => n8311, C1 => n13797, C2 => 
                           n8279, A => n5737, ZN => n5736);
   U4412 : OAI222_X1 port map( A1 => n6978, A2 => n13794, B1 => n6980, B2 => 
                           n13791, C1 => n1572, C2 => n13788, ZN => n5737);
   U4413 : AOI221_X1 port map( B1 => n13746, B2 => n8629, C1 => n13743, C2 => 
                           n8597, A => n5745, ZN => n5744);
   U4414 : OAI222_X1 port map( A1 => n6972, A2 => n13740, B1 => n6974, B2 => 
                           n13737, C1 => n1301, C2 => n13734, ZN => n5745);
   U4415 : AOI221_X1 port map( B1 => n13692, B2 => n8883, C1 => n13689, C2 => 
                           n8851, A => n5753, ZN => n5752);
   U4416 : OAI222_X1 port map( A1 => n6966, A2 => n13686, B1 => n6968, B2 => 
                           n13683, C1 => n635, C2 => n13680, ZN => n5753);
   U4417 : AOI221_X1 port map( B1 => n14074, B2 => n8120, C1 => n14071, C2 => 
                           n8088, A => n4445, ZN => n4444);
   U4418 : OAI222_X1 port map( A1 => n7008, A2 => n14068, B1 => n7010, B2 => 
                           n14065, C1 => n1703, C2 => n14062, ZN => n4445);
   U4419 : AOI221_X1 port map( B1 => n14019, B2 => n8310, C1 => n14016, C2 => 
                           n8278, A => n4453, ZN => n4452);
   U4420 : OAI222_X1 port map( A1 => n7002, A2 => n14013, B1 => n7004, B2 => 
                           n14011, C1 => n1571, C2 => n14007, ZN => n4453);
   U4421 : AOI221_X1 port map( B1 => n13965, B2 => n8628, C1 => n13962, C2 => 
                           n8596, A => n4461, ZN => n4460);
   U4422 : OAI222_X1 port map( A1 => n6996, A2 => n13959, B1 => n6998, B2 => 
                           n13957, C1 => n1300, C2 => n13953, ZN => n4461);
   U4423 : AOI221_X1 port map( B1 => n13923, B2 => n8882, C1 => n13920, C2 => 
                           n8850, A => n4469, ZN => n4468);
   U4424 : OAI222_X1 port map( A1 => n6990, A2 => n13918, B1 => n6992, B2 => 
                           n13915, C1 => n634, C2 => n13912, ZN => n4469);
   U4425 : AOI221_X1 port map( B1 => n13800, B2 => n8310, C1 => n13797, C2 => 
                           n8278, A => n5774, ZN => n5773);
   U4426 : OAI222_X1 port map( A1 => n7002, A2 => n13794, B1 => n7004, B2 => 
                           n13791, C1 => n1571, C2 => n13788, ZN => n5774);
   U4427 : AOI221_X1 port map( B1 => n13746, B2 => n8628, C1 => n13743, C2 => 
                           n8596, A => n5782, ZN => n5781);
   U4428 : OAI222_X1 port map( A1 => n6996, A2 => n13740, B1 => n6998, B2 => 
                           n13737, C1 => n1300, C2 => n13734, ZN => n5782);
   U4429 : AOI221_X1 port map( B1 => n13692, B2 => n8882, C1 => n13689, C2 => 
                           n8850, A => n5790, ZN => n5789);
   U4430 : OAI222_X1 port map( A1 => n6990, A2 => n13686, B1 => n6992, B2 => 
                           n13683, C1 => n634, C2 => n13680, ZN => n5790);
   U4431 : AOI221_X1 port map( B1 => n13965, B2 => n8627, C1 => n13963, C2 => 
                           n8595, A => n4498, ZN => n4497);
   U4432 : OAI222_X1 port map( A1 => n7020, A2 => n13960, B1 => n7022, B2 => 
                           n13957, C1 => n1299, C2 => n13954, ZN => n4498);
   U4433 : AOI221_X1 port map( B1 => n13923, B2 => n8881, C1 => n13921, C2 => 
                           n8849, A => n4506, ZN => n4505);
   U4434 : OAI222_X1 port map( A1 => n7014, A2 => n13918, B1 => n7016, B2 => 
                           n13915, C1 => n633, C2 => n13912, ZN => n4506);
   U4435 : AOI221_X1 port map( B1 => n13800, B2 => n8309, C1 => n13797, C2 => 
                           n8277, A => n5811, ZN => n5810);
   U4436 : OAI222_X1 port map( A1 => n1564, A2 => n13794, B1 => n7028, B2 => 
                           n13791, C1 => n1570, C2 => n13788, ZN => n5811);
   U4437 : AOI221_X1 port map( B1 => n13746, B2 => n8627, C1 => n13743, C2 => 
                           n8595, A => n5819, ZN => n5818);
   U4438 : OAI222_X1 port map( A1 => n7020, A2 => n13740, B1 => n7022, B2 => 
                           n13737, C1 => n1299, C2 => n13734, ZN => n5819);
   U4439 : AOI221_X1 port map( B1 => n13692, B2 => n8881, C1 => n13689, C2 => 
                           n8849, A => n5827, ZN => n5826);
   U4440 : OAI222_X1 port map( A1 => n7014, A2 => n13686, B1 => n7016, B2 => 
                           n13683, C1 => n633, C2 => n13680, ZN => n5827);
   U4441 : AOI221_X1 port map( B1 => n14074, B2 => n8118, C1 => n14071, C2 => 
                           n8086, A => n4519, ZN => n4518);
   U4442 : OAI222_X1 port map( A1 => n1695, A2 => n14068, B1 => n7058, B2 => 
                           n14065, C1 => n1701, C2 => n14062, ZN => n4519);
   U4443 : AOI221_X1 port map( B1 => n13965, B2 => n8626, C1 => n13963, C2 => 
                           n8594, A => n4535, ZN => n4534);
   U4444 : OAI222_X1 port map( A1 => n1293, A2 => n13960, B1 => n7046, B2 => 
                           n13957, C1 => n1298, C2 => n13954, ZN => n4535);
   U4445 : AOI221_X1 port map( B1 => n13923, B2 => n8880, C1 => n13921, C2 => 
                           n8848, A => n4543, ZN => n4542);
   U4446 : OAI222_X1 port map( A1 => n7038, A2 => n13918, B1 => n7040, B2 => 
                           n13915, C1 => n632, C2 => n13912, ZN => n4543);
   U4447 : AOI221_X1 port map( B1 => n13800, B2 => n8308, C1 => n13797, C2 => 
                           n8276, A => n5848, ZN => n5847);
   U4448 : OAI222_X1 port map( A1 => n1563, A2 => n13794, B1 => n7052, B2 => 
                           n13791, C1 => n1569, C2 => n13788, ZN => n5848);
   U4449 : AOI221_X1 port map( B1 => n13746, B2 => n8626, C1 => n13743, C2 => 
                           n8594, A => n5856, ZN => n5855);
   U4450 : OAI222_X1 port map( A1 => n1293, A2 => n13740, B1 => n7046, B2 => 
                           n13737, C1 => n1298, C2 => n13734, ZN => n5856);
   U4451 : AOI221_X1 port map( B1 => n13692, B2 => n8880, C1 => n13689, C2 => 
                           n8848, A => n5864, ZN => n5863);
   U4452 : OAI222_X1 port map( A1 => n7038, A2 => n13686, B1 => n7040, B2 => 
                           n13683, C1 => n632, C2 => n13680, ZN => n5864);
   U4453 : AOI221_X1 port map( B1 => n14074, B2 => n8117, C1 => n14071, C2 => 
                           n8085, A => n4556, ZN => n4555);
   U4454 : OAI222_X1 port map( A1 => n1694, A2 => n14068, B1 => n7082, B2 => 
                           n14065, C1 => n1700, C2 => n14062, ZN => n4556);
   U4455 : AOI221_X1 port map( B1 => n13966, B2 => n8625, C1 => n13963, C2 => 
                           n8593, A => n4572, ZN => n4571);
   U4456 : OAI222_X1 port map( A1 => n1292, A2 => n13960, B1 => n7070, B2 => 
                           n13957, C1 => n1297, C2 => n13954, ZN => n4572);
   U4457 : AOI221_X1 port map( B1 => n13924, B2 => n8879, C1 => n13921, C2 => 
                           n8847, A => n4580, ZN => n4579);
   U4458 : OAI222_X1 port map( A1 => n7062, A2 => n13918, B1 => n7064, B2 => 
                           n13915, C1 => n631, C2 => n13912, ZN => n4580);
   U4459 : AOI221_X1 port map( B1 => n13800, B2 => n8307, C1 => n13797, C2 => 
                           n8275, A => n5885, ZN => n5884);
   U4460 : OAI222_X1 port map( A1 => n1562, A2 => n13794, B1 => n7076, B2 => 
                           n13791, C1 => n1568, C2 => n13788, ZN => n5885);
   U4461 : AOI221_X1 port map( B1 => n13746, B2 => n8625, C1 => n13743, C2 => 
                           n8593, A => n5893, ZN => n5892);
   U4462 : OAI222_X1 port map( A1 => n1292, A2 => n13740, B1 => n7070, B2 => 
                           n13737, C1 => n1297, C2 => n13734, ZN => n5893);
   U4463 : AOI221_X1 port map( B1 => n13692, B2 => n8879, C1 => n13689, C2 => 
                           n8847, A => n5901, ZN => n5900);
   U4464 : OAI222_X1 port map( A1 => n7062, A2 => n13686, B1 => n7064, B2 => 
                           n13683, C1 => n631, C2 => n13680, ZN => n5901);
   U4465 : AOI221_X1 port map( B1 => n14074, B2 => n8116, C1 => n14071, C2 => 
                           n8084, A => n4593, ZN => n4592);
   U4466 : OAI222_X1 port map( A1 => n1693, A2 => n14068, B1 => n7106, B2 => 
                           n14065, C1 => n1699, C2 => n14062, ZN => n4593);
   U4467 : AOI221_X1 port map( B1 => n13966, B2 => n8624, C1 => n13963, C2 => 
                           n8592, A => n4609, ZN => n4608);
   U4468 : OAI222_X1 port map( A1 => n1291, A2 => n13960, B1 => n7094, B2 => 
                           n13957, C1 => n1296, C2 => n13954, ZN => n4609);
   U4469 : AOI221_X1 port map( B1 => n13924, B2 => n8878, C1 => n13921, C2 => 
                           n8846, A => n4617, ZN => n4616);
   U4470 : OAI222_X1 port map( A1 => n7086, A2 => n13918, B1 => n7088, B2 => 
                           n13915, C1 => n630, C2 => n13912, ZN => n4617);
   U4471 : AOI221_X1 port map( B1 => n13800, B2 => n8306, C1 => n13797, C2 => 
                           n8274, A => n5922, ZN => n5921);
   U4472 : OAI222_X1 port map( A1 => n1561, A2 => n13794, B1 => n7100, B2 => 
                           n13791, C1 => n1567, C2 => n13788, ZN => n5922);
   U4473 : AOI221_X1 port map( B1 => n13746, B2 => n8624, C1 => n13743, C2 => 
                           n8592, A => n5930, ZN => n5929);
   U4474 : OAI222_X1 port map( A1 => n1291, A2 => n13740, B1 => n7094, B2 => 
                           n13737, C1 => n1296, C2 => n13734, ZN => n5930);
   U4475 : AOI221_X1 port map( B1 => n13692, B2 => n8878, C1 => n13689, C2 => 
                           n8846, A => n5938, ZN => n5937);
   U4476 : OAI222_X1 port map( A1 => n7086, A2 => n13686, B1 => n7088, B2 => 
                           n13683, C1 => n630, C2 => n13680, ZN => n5938);
   U4477 : AOI221_X1 port map( B1 => n14074, B2 => n8115, C1 => n14071, C2 => 
                           n8083, A => n4630, ZN => n4629);
   U4478 : OAI222_X1 port map( A1 => n1692, A2 => n14068, B1 => n7130, B2 => 
                           n14065, C1 => n1698, C2 => n14062, ZN => n4630);
   U4479 : AOI221_X1 port map( B1 => n13966, B2 => n8623, C1 => n13963, C2 => 
                           n8591, A => n4646, ZN => n4645);
   U4480 : OAI222_X1 port map( A1 => n1290, A2 => n13960, B1 => n7118, B2 => 
                           n13957, C1 => n1295, C2 => n13954, ZN => n4646);
   U4481 : AOI221_X1 port map( B1 => n13924, B2 => n8877, C1 => n13921, C2 => 
                           n8845, A => n4654, ZN => n4653);
   U4482 : OAI222_X1 port map( A1 => n7110, A2 => n13918, B1 => n7112, B2 => 
                           n13915, C1 => n629, C2 => n13912, ZN => n4654);
   U4483 : AOI221_X1 port map( B1 => n13800, B2 => n8305, C1 => n13797, C2 => 
                           n8273, A => n5959, ZN => n5958);
   U4484 : OAI222_X1 port map( A1 => n1560, A2 => n13794, B1 => n7124, B2 => 
                           n13791, C1 => n1566, C2 => n13788, ZN => n5959);
   U4485 : AOI221_X1 port map( B1 => n13746, B2 => n8623, C1 => n13743, C2 => 
                           n8591, A => n5967, ZN => n5966);
   U4486 : OAI222_X1 port map( A1 => n1290, A2 => n13740, B1 => n7118, B2 => 
                           n13737, C1 => n1295, C2 => n13734, ZN => n5967);
   U4487 : AOI221_X1 port map( B1 => n13692, B2 => n8877, C1 => n13689, C2 => 
                           n8845, A => n5975, ZN => n5974);
   U4488 : OAI222_X1 port map( A1 => n7110, A2 => n13686, B1 => n7112, B2 => 
                           n13683, C1 => n629, C2 => n13680, ZN => n5975);
   U4489 : AOI221_X1 port map( B1 => n14074, B2 => n8114, C1 => n14071, C2 => 
                           n8082, A => n4667, ZN => n4666);
   U4490 : OAI222_X1 port map( A1 => n7152, A2 => n14068, B1 => n7154, B2 => 
                           n14065, C1 => n1697, C2 => n14062, ZN => n4667);
   U4491 : AOI221_X1 port map( B1 => n13966, B2 => n8622, C1 => n13963, C2 => 
                           n8590, A => n4683, ZN => n4682);
   U4492 : OAI222_X1 port map( A1 => n1289, A2 => n13960, B1 => n7142, B2 => 
                           n13957, C1 => n1294, C2 => n13954, ZN => n4683);
   U4493 : AOI221_X1 port map( B1 => n13924, B2 => n8876, C1 => n13921, C2 => 
                           n8844, A => n4691, ZN => n4690);
   U4494 : OAI222_X1 port map( A1 => n7134, A2 => n13918, B1 => n7136, B2 => 
                           n13915, C1 => n628, C2 => n13912, ZN => n4691);
   U4495 : AOI221_X1 port map( B1 => n13800, B2 => n8304, C1 => n13797, C2 => 
                           n8272, A => n5996, ZN => n5995);
   U4496 : OAI222_X1 port map( A1 => n7146, A2 => n13794, B1 => n7148, B2 => 
                           n13791, C1 => n1565, C2 => n13788, ZN => n5996);
   U4497 : AOI221_X1 port map( B1 => n13746, B2 => n8622, C1 => n13743, C2 => 
                           n8590, A => n6004, ZN => n6003);
   U4498 : OAI222_X1 port map( A1 => n1289, A2 => n13740, B1 => n7142, B2 => 
                           n13737, C1 => n1294, C2 => n13734, ZN => n6004);
   U4499 : AOI221_X1 port map( B1 => n13692, B2 => n8876, C1 => n13689, C2 => 
                           n8844, A => n6012, ZN => n6011);
   U4500 : OAI222_X1 port map( A1 => n7134, A2 => n13686, B1 => n7136, B2 => 
                           n13683, C1 => n628, C2 => n13680, ZN => n6012);
   U4501 : AOI221_X1 port map( B1 => n14270, B2 => n1740, C1 => n7469, C2 => 
                           n14267, A => n6568, ZN => n6567);
   U4502 : OAI222_X1 port map( A1 => n14264, A2 => n115, B1 => n14261, B2 => 
                           n131, C1 => n14258, C2 => n107, ZN => n6568);
   U4503 : AOI221_X1 port map( B1 => n14216, B2 => n1766, C1 => n830, C2 => 
                           n14213, A => n6581, ZN => n6580);
   U4504 : OAI222_X1 port map( A1 => n14210, A2 => n228, B1 => n7812, B2 => 
                           n14207, C1 => n14204, C2 => n220, ZN => n6581);
   U4505 : AOI221_X1 port map( B1 => n14271, B2 => n1739, C1 => n7491, C2 => 
                           n14268, A => n2789, ZN => n2786);
   U4506 : OAI222_X1 port map( A1 => n14266, A2 => n114, B1 => n14263, B2 => 
                           n130, C1 => n14260, C2 => n106, ZN => n2789);
   U4507 : AOI221_X1 port map( B1 => n14217, B2 => n1765, C1 => n14214, C2 => 
                           n1773, A => n2815, ZN => n2812);
   U4508 : OAI222_X1 port map( A1 => n14212, A2 => n227, B1 => n7808, B2 => 
                           n14209, C1 => n14206, C2 => n219, ZN => n2815);
   U4509 : AOI221_X1 port map( B1 => n14216, B2 => n1764, C1 => n14213, C2 => 
                           n1772, A => n2895, ZN => n2894);
   U4510 : OAI222_X1 port map( A1 => n14212, A2 => n226, B1 => n7804, B2 => 
                           n14209, C1 => n14206, C2 => n218, ZN => n2895);
   U4511 : AOI221_X1 port map( B1 => n14075, B2 => n8128, C1 => n14072, C2 => 
                           n8096, A => n4149, ZN => n4148);
   U4512 : OAI222_X1 port map( A1 => n6816, A2 => n14069, B1 => n6818, B2 => 
                           n14066, C1 => n409, C2 => n14063, ZN => n4149);
   U4513 : AOI221_X1 port map( B1 => n13923, B2 => n8890, C1 => n13920, C2 => 
                           n8858, A => n4173, ZN => n4172);
   U4514 : OAI222_X1 port map( A1 => n6798, A2 => n13919, B1 => n6800, B2 => 
                           n13916, C1 => n5, C2 => n13913, ZN => n4173);
   U4515 : AOI221_X1 port map( B1 => n14075, B2 => n8127, C1 => n14072, C2 => 
                           n8095, A => n4186, ZN => n4185);
   U4516 : OAI222_X1 port map( A1 => n6840, A2 => n14069, B1 => n6842, B2 => 
                           n14066, C1 => n408, C2 => n14063, ZN => n4186);
   U4517 : AOI221_X1 port map( B1 => n14019, B2 => n8317, C1 => n14016, C2 => 
                           n8285, A => n4194, ZN => n4193);
   U4518 : OAI222_X1 port map( A1 => n6834, A2 => n14013, B1 => n6836, B2 => 
                           n14012, C1 => n232, C2 => n14007, ZN => n4194);
   U4519 : AOI221_X1 port map( B1 => n13965, B2 => n8635, C1 => n13962, C2 => 
                           n8603, A => n4202, ZN => n4201);
   U4520 : OAI222_X1 port map( A1 => n6828, A2 => n13959, B1 => n6830, B2 => 
                           n13958, C1 => n136, C2 => n13953, ZN => n4202);
   U4521 : AOI221_X1 port map( B1 => n14075, B2 => n8126, C1 => n14072, C2 => 
                           n8094, A => n4223, ZN => n4222);
   U4522 : OAI222_X1 port map( A1 => n6864, A2 => n14069, B1 => n6866, B2 => 
                           n14066, C1 => n407, C2 => n14063, ZN => n4223);
   U4523 : AOI221_X1 port map( B1 => n14270, B2 => n1738, C1 => n7492, C2 => 
                           n14267, A => n2887, ZN => n2886);
   U4524 : OAI222_X1 port map( A1 => n14266, A2 => n113, B1 => n14263, B2 => 
                           n129, C1 => n14260, C2 => n105, ZN => n2887);
   U4525 : AOI221_X1 port map( B1 => n14270, B2 => n1737, C1 => n7493, C2 => 
                           n14267, A => n2924, ZN => n2923);
   U4526 : OAI222_X1 port map( A1 => n14266, A2 => n112, B1 => n14263, B2 => 
                           n128, C1 => n14260, C2 => n104, ZN => n2924);
   U4527 : AOI221_X1 port map( B1 => n14216, B2 => n1763, C1 => n14213, C2 => 
                           n1771, A => n2932, ZN => n2931);
   U4528 : OAI222_X1 port map( A1 => n14212, A2 => n225, B1 => n7800, B2 => 
                           n14209, C1 => n14206, C2 => n217, ZN => n2932);
   U4529 : AOI221_X1 port map( B1 => n13923, B2 => n8889, C1 => n13920, C2 => 
                           n8857, A => n4210, ZN => n4209);
   U4530 : OAI222_X1 port map( A1 => n6822, A2 => n13919, B1 => n6824, B2 => 
                           n13916, C1 => n4, C2 => n13913, ZN => n4210);
   U4531 : AOI221_X1 port map( B1 => n14270, B2 => n1736, C1 => n7494, C2 => 
                           n14267, A => n2961, ZN => n2960);
   U4532 : OAI222_X1 port map( A1 => n14266, A2 => n111, B1 => n14263, B2 => 
                           n127, C1 => n14260, C2 => n103, ZN => n2961);
   U4533 : AOI221_X1 port map( B1 => n14216, B2 => n1762, C1 => n14213, C2 => 
                           n1770, A => n2969, ZN => n2968);
   U4534 : OAI222_X1 port map( A1 => n14212, A2 => n224, B1 => n7796, B2 => 
                           n14209, C1 => n14206, C2 => n216, ZN => n2969);
   U4535 : AOI221_X1 port map( B1 => n14270, B2 => n1735, C1 => n7495, C2 => 
                           n14267, A => n2998, ZN => n2997);
   U4536 : OAI222_X1 port map( A1 => n14266, A2 => n110, B1 => n14263, B2 => 
                           n126, C1 => n14260, C2 => n102, ZN => n2998);
   U4537 : AOI221_X1 port map( B1 => n14216, B2 => n1761, C1 => n14213, C2 => 
                           n1769, A => n3006, ZN => n3005);
   U4538 : OAI222_X1 port map( A1 => n14212, A2 => n223, B1 => n7792, B2 => 
                           n14209, C1 => n14206, C2 => n215, ZN => n3006);
   U4539 : AOI221_X1 port map( B1 => n14270, B2 => n1734, C1 => n7497, C2 => 
                           n14267, A => n3035, ZN => n3034);
   U4540 : OAI222_X1 port map( A1 => n14266, A2 => n109, B1 => n14263, B2 => 
                           n125, C1 => n14260, C2 => n101, ZN => n3035);
   U4541 : AOI221_X1 port map( B1 => n14216, B2 => n1760, C1 => n14213, C2 => 
                           n1768, A => n3043, ZN => n3042);
   U4542 : OAI222_X1 port map( A1 => n14212, A2 => n222, B1 => n7788, B2 => 
                           n14209, C1 => n14206, C2 => n214, ZN => n3043);
   U4543 : AOI221_X1 port map( B1 => n14270, B2 => n1733, C1 => n7499, C2 => 
                           n14267, A => n3072, ZN => n3071);
   U4544 : OAI222_X1 port map( A1 => n14266, A2 => n108, B1 => n14263, B2 => 
                           n124, C1 => n14260, C2 => n100, ZN => n3072);
   U4545 : AOI221_X1 port map( B1 => n14216, B2 => n1759, C1 => n14213, C2 => 
                           n1767, A => n3080, ZN => n3079);
   U4546 : OAI222_X1 port map( A1 => n14212, A2 => n221, B1 => n7784, B2 => 
                           n14209, C1 => n14206, C2 => n213, ZN => n3080);
   U4547 : AOI221_X1 port map( B1 => n14270, B2 => n2066, C1 => n7500, C2 => 
                           n14267, A => n3109, ZN => n3108);
   U4548 : OAI222_X1 port map( A1 => n14266, A2 => n1240, B1 => n14263, B2 => 
                           n1288, C1 => n14260, C2 => n1216, ZN => n3109);
   U4549 : AOI221_X1 port map( B1 => n14216, B2 => n2303, C1 => n14213, C2 => 
                           n2326, A => n3117, ZN => n3116);
   U4550 : OAI222_X1 port map( A1 => n14212, A2 => n1559, B1 => n7780, B2 => 
                           n14209, C1 => n14206, C2 => n1535, ZN => n3117);
   U4551 : AOI221_X1 port map( B1 => n14270, B2 => n2065, C1 => n7501, C2 => 
                           n14267, A => n3146, ZN => n3145);
   U4552 : OAI222_X1 port map( A1 => n14265, A2 => n1239, B1 => n14262, B2 => 
                           n1287, C1 => n14259, C2 => n1215, ZN => n3146);
   U4553 : AOI221_X1 port map( B1 => n14216, B2 => n2302, C1 => n14213, C2 => 
                           n2325, A => n3154, ZN => n3153);
   U4554 : OAI222_X1 port map( A1 => n14211, A2 => n1558, B1 => n7776, B2 => 
                           n14208, C1 => n14205, C2 => n1534, ZN => n3154);
   U4555 : AOI221_X1 port map( B1 => n14270, B2 => n2064, C1 => n7503, C2 => 
                           n14267, A => n3183, ZN => n3182);
   U4556 : OAI222_X1 port map( A1 => n14265, A2 => n1238, B1 => n14262, B2 => 
                           n1286, C1 => n14259, C2 => n1214, ZN => n3183);
   U4557 : AOI221_X1 port map( B1 => n14216, B2 => n2301, C1 => n14213, C2 => 
                           n2324, A => n3191, ZN => n3190);
   U4558 : OAI222_X1 port map( A1 => n14211, A2 => n1557, B1 => n7772, B2 => 
                           n14208, C1 => n14205, C2 => n1533, ZN => n3191);
   U4559 : AOI221_X1 port map( B1 => n14270, B2 => n2063, C1 => n7505, C2 => 
                           n14267, A => n3220, ZN => n3219);
   U4560 : OAI222_X1 port map( A1 => n14265, A2 => n1237, B1 => n14262, B2 => 
                           n1285, C1 => n14259, C2 => n1213, ZN => n3220);
   U4561 : AOI221_X1 port map( B1 => n14216, B2 => n2300, C1 => n14214, C2 => 
                           n2323, A => n3228, ZN => n3227);
   U4562 : OAI222_X1 port map( A1 => n14211, A2 => n1556, B1 => n7768, B2 => 
                           n14208, C1 => n14205, C2 => n1532, ZN => n3228);
   U4563 : AOI221_X1 port map( B1 => n14074, B2 => n8119, C1 => n14071, C2 => 
                           n8087, A => n4482, ZN => n4481);
   U4564 : OAI222_X1 port map( A1 => n1696, A2 => n14068, B1 => n7034, B2 => 
                           n14065, C1 => n1702, C2 => n14062, ZN => n4482);
   U4565 : AOI221_X1 port map( B1 => n14270, B2 => n2062, C1 => n7506, C2 => 
                           n14267, A => n3257, ZN => n3256);
   U4566 : OAI222_X1 port map( A1 => n14265, A2 => n1236, B1 => n14262, B2 => 
                           n1284, C1 => n14259, C2 => n1212, ZN => n3257);
   U4567 : AOI221_X1 port map( B1 => n14216, B2 => n2299, C1 => n14214, C2 => 
                           n2322, A => n3265, ZN => n3264);
   U4568 : OAI222_X1 port map( A1 => n14211, A2 => n1555, B1 => n7764, B2 => 
                           n14208, C1 => n14205, C2 => n1531, ZN => n3265);
   U4569 : AOI221_X1 port map( B1 => n14271, B2 => n2061, C1 => n7507, C2 => 
                           n14268, A => n3294, ZN => n3293);
   U4570 : OAI222_X1 port map( A1 => n14265, A2 => n1235, B1 => n14262, B2 => 
                           n1283, C1 => n14259, C2 => n1211, ZN => n3294);
   U4571 : AOI221_X1 port map( B1 => n14217, B2 => n2298, C1 => n14214, C2 => 
                           n2321, A => n3302, ZN => n3301);
   U4572 : OAI222_X1 port map( A1 => n14211, A2 => n1554, B1 => n7760, B2 => 
                           n14208, C1 => n14205, C2 => n1530, ZN => n3302);
   U4573 : AOI221_X1 port map( B1 => n14271, B2 => n2060, C1 => n7509, C2 => 
                           n14268, A => n3333, ZN => n3332);
   U4574 : OAI222_X1 port map( A1 => n14265, A2 => n1234, B1 => n14262, B2 => 
                           n1282, C1 => n14259, C2 => n1210, ZN => n3333);
   U4575 : AOI221_X1 port map( B1 => n14217, B2 => n2297, C1 => n14214, C2 => 
                           n2320, A => n3341, ZN => n3340);
   U4576 : OAI222_X1 port map( A1 => n14211, A2 => n1553, B1 => n7756, B2 => 
                           n14208, C1 => n14205, C2 => n1529, ZN => n3341);
   U4577 : AOI221_X1 port map( B1 => n14271, B2 => n2059, C1 => n7511, C2 => 
                           n14268, A => n3370, ZN => n3369);
   U4578 : OAI222_X1 port map( A1 => n14265, A2 => n1233, B1 => n14262, B2 => 
                           n1281, C1 => n14259, C2 => n1209, ZN => n3370);
   U4579 : AOI221_X1 port map( B1 => n14217, B2 => n2296, C1 => n14214, C2 => 
                           n2319, A => n3378, ZN => n3377);
   U4580 : OAI222_X1 port map( A1 => n14211, A2 => n1552, B1 => n7752, B2 => 
                           n14208, C1 => n14205, C2 => n1528, ZN => n3378);
   U4581 : AOI221_X1 port map( B1 => n14271, B2 => n2058, C1 => n7512, C2 => 
                           n14268, A => n3407, ZN => n3406);
   U4582 : OAI222_X1 port map( A1 => n14265, A2 => n1232, B1 => n14262, B2 => 
                           n1280, C1 => n14259, C2 => n1208, ZN => n3407);
   U4583 : AOI221_X1 port map( B1 => n14217, B2 => n2295, C1 => n14214, C2 => 
                           n2318, A => n3415, ZN => n3414);
   U4584 : OAI222_X1 port map( A1 => n14211, A2 => n1551, B1 => n7748, B2 => 
                           n14208, C1 => n14205, C2 => n1527, ZN => n3415);
   U4585 : AOI221_X1 port map( B1 => n14271, B2 => n2057, C1 => n7513, C2 => 
                           n14268, A => n3444, ZN => n3443);
   U4586 : OAI222_X1 port map( A1 => n14265, A2 => n1231, B1 => n14262, B2 => 
                           n1279, C1 => n14259, C2 => n1207, ZN => n3444);
   U4587 : AOI221_X1 port map( B1 => n14217, B2 => n2294, C1 => n14214, C2 => 
                           n2317, A => n3452, ZN => n3451);
   U4588 : OAI222_X1 port map( A1 => n14211, A2 => n1550, B1 => n7744, B2 => 
                           n14208, C1 => n14205, C2 => n1526, ZN => n3452);
   U4589 : AOI221_X1 port map( B1 => n14271, B2 => n2056, C1 => n7515, C2 => 
                           n14268, A => n3481, ZN => n3480);
   U4590 : OAI222_X1 port map( A1 => n14265, A2 => n1230, B1 => n14262, B2 => 
                           n1278, C1 => n14259, C2 => n1206, ZN => n3481);
   U4591 : AOI221_X1 port map( B1 => n14217, B2 => n2293, C1 => n14214, C2 => 
                           n2316, A => n3489, ZN => n3488);
   U4592 : OAI222_X1 port map( A1 => n14211, A2 => n1549, B1 => n7740, B2 => 
                           n14208, C1 => n14205, C2 => n1525, ZN => n3489);
   U4593 : AOI221_X1 port map( B1 => n14271, B2 => n2055, C1 => n7517, C2 => 
                           n14268, A => n3518, ZN => n3517);
   U4594 : OAI222_X1 port map( A1 => n14265, A2 => n1229, B1 => n14262, B2 => 
                           n1277, C1 => n14259, C2 => n1205, ZN => n3518);
   U4595 : AOI221_X1 port map( B1 => n14217, B2 => n2292, C1 => n14214, C2 => 
                           n2315, A => n3526, ZN => n3525);
   U4596 : OAI222_X1 port map( A1 => n14211, A2 => n1548, B1 => n7736, B2 => 
                           n14208, C1 => n14205, C2 => n1524, ZN => n3526);
   U4597 : AOI221_X1 port map( B1 => n14163, B2 => n825, C1 => n14160, C2 => 
                           n1659, A => n3534, ZN => n3533);
   U4598 : OAI222_X1 port map( A1 => n2468, A2 => n14157, B1 => n1680, B2 => 
                           n14154, C1 => n2447, C2 => n14151, ZN => n3534);
   U4599 : AOI221_X1 port map( B1 => n791, B2 => n14272, C1 => n14269, C2 => 
                           n1252, A => n3555, ZN => n3554);
   U4600 : OAI222_X1 port map( A1 => n14265, A2 => n1228, B1 => n14262, B2 => 
                           n1276, C1 => n14259, C2 => n1204, ZN => n3555);
   U4601 : AOI221_X1 port map( B1 => n777, B2 => n14218, C1 => n774, C2 => 
                           n14213, A => n3563, ZN => n3562);
   U4602 : OAI222_X1 port map( A1 => n14211, A2 => n1547, B1 => n7732, B2 => 
                           n14208, C1 => n14205, C2 => n1523, ZN => n3563);
   U4603 : AOI221_X1 port map( B1 => n727, B2 => n14272, C1 => n7519, C2 => 
                           n14268, A => n3592, ZN => n3591);
   U4604 : OAI222_X1 port map( A1 => n14264, A2 => n1227, B1 => n14261, B2 => 
                           n1275, C1 => n14258, C2 => n1203, ZN => n3592);
   U4605 : AOI221_X1 port map( B1 => n14217, B2 => n2290, C1 => n14214, C2 => 
                           n2313, A => n3600, ZN => n3599);
   U4606 : OAI222_X1 port map( A1 => n14210, A2 => n1546, B1 => n7728, B2 => 
                           n14207, C1 => n14204, C2 => n1522, ZN => n3600);
   U4607 : AOI221_X1 port map( B1 => n14271, B2 => n2052, C1 => n7521, C2 => 
                           n14268, A => n3629, ZN => n3628);
   U4608 : OAI222_X1 port map( A1 => n14264, A2 => n1226, B1 => n14261, B2 => 
                           n1274, C1 => n14258, C2 => n1202, ZN => n3629);
   U4609 : AOI221_X1 port map( B1 => n14217, B2 => n2289, C1 => n14214, C2 => 
                           n2312, A => n3637, ZN => n3636);
   U4610 : OAI222_X1 port map( A1 => n14210, A2 => n1545, B1 => n7724, B2 => 
                           n14207, C1 => n14204, C2 => n1521, ZN => n3637);
   U4611 : AOI221_X1 port map( B1 => n14271, B2 => n2051, C1 => n7523, C2 => 
                           n14268, A => n3666, ZN => n3665);
   U4612 : OAI222_X1 port map( A1 => n14264, A2 => n1225, B1 => n14261, B2 => 
                           n1273, C1 => n14258, C2 => n1201, ZN => n3666);
   U4613 : AOI221_X1 port map( B1 => n14217, B2 => n2288, C1 => n14214, C2 => 
                           n2311, A => n3674, ZN => n3673);
   U4614 : OAI222_X1 port map( A1 => n14210, A2 => n1544, B1 => n7720, B2 => 
                           n14207, C1 => n14204, C2 => n1520, ZN => n3674);
   U4615 : AOI221_X1 port map( B1 => n14271, B2 => n2050, C1 => n7524, C2 => 
                           n14268, A => n3703, ZN => n3702);
   U4616 : OAI222_X1 port map( A1 => n14264, A2 => n1224, B1 => n14261, B2 => 
                           n1272, C1 => n14258, C2 => n1200, ZN => n3703);
   U4618 : AOI221_X1 port map( B1 => n14217, B2 => n2287, C1 => n14215, C2 => 
                           n2310, A => n3711, ZN => n3710);
   U4619 : OAI222_X1 port map( A1 => n14210, A2 => n1543, B1 => n7716, B2 => 
                           n14207, C1 => n14204, C2 => n1519, ZN => n3711);
   U4620 : AOI221_X1 port map( B1 => n14271, B2 => n2049, C1 => n7525, C2 => 
                           n14269, A => n3740, ZN => n3739);
   U4621 : OAI222_X1 port map( A1 => n14264, A2 => n1223, B1 => n14261, B2 => 
                           n1271, C1 => n14258, C2 => n1199, ZN => n3740);
   U4622 : AOI221_X1 port map( B1 => n14218, B2 => n2286, C1 => n14215, C2 => 
                           n2309, A => n3748, ZN => n3747);
   U4623 : OAI222_X1 port map( A1 => n14210, A2 => n1542, B1 => n7712, B2 => 
                           n14207, C1 => n14204, C2 => n1518, ZN => n3748);
   U4624 : AOI221_X1 port map( B1 => n14272, B2 => n2048, C1 => n7527, C2 => 
                           n14269, A => n3777, ZN => n3776);
   U4625 : OAI222_X1 port map( A1 => n14264, A2 => n1222, B1 => n14261, B2 => 
                           n1270, C1 => n14258, C2 => n1198, ZN => n3777);
   U4626 : AOI221_X1 port map( B1 => n14218, B2 => n2285, C1 => n14215, C2 => 
                           n2308, A => n3785, ZN => n3784);
   U4627 : OAI222_X1 port map( A1 => n14210, A2 => n1541, B1 => n7708, B2 => 
                           n14207, C1 => n14204, C2 => n1517, ZN => n3785);
   U4628 : AOI221_X1 port map( B1 => n14272, B2 => n2047, C1 => n7529, C2 => 
                           n14269, A => n3814, ZN => n3813);
   U4629 : OAI222_X1 port map( A1 => n14264, A2 => n1221, B1 => n14261, B2 => 
                           n1269, C1 => n14258, C2 => n1197, ZN => n3814);
   U4630 : AOI221_X1 port map( B1 => n14218, B2 => n2284, C1 => n14215, C2 => 
                           n2307, A => n3822, ZN => n3821);
   U4631 : OAI222_X1 port map( A1 => n14210, A2 => n1540, B1 => n7704, B2 => 
                           n14207, C1 => n14204, C2 => n1516, ZN => n3822);
   U4632 : AOI221_X1 port map( B1 => n14272, B2 => n2046, C1 => n7530, C2 => 
                           n14269, A => n3851, ZN => n3850);
   U4633 : OAI222_X1 port map( A1 => n14264, A2 => n1220, B1 => n14261, B2 => 
                           n1268, C1 => n14258, C2 => n1196, ZN => n3851);
   U4634 : AOI221_X1 port map( B1 => n14218, B2 => n2283, C1 => n14215, C2 => 
                           n2306, A => n3859, ZN => n3858);
   U4635 : OAI222_X1 port map( A1 => n14210, A2 => n1539, B1 => n7700, B2 => 
                           n14207, C1 => n14204, C2 => n1515, ZN => n3859);
   U4636 : AOI221_X1 port map( B1 => n14272, B2 => n2045, C1 => n7531, C2 => 
                           n14269, A => n3888, ZN => n3887);
   U4637 : OAI222_X1 port map( A1 => n14264, A2 => n1219, B1 => n14261, B2 => 
                           n1267, C1 => n14258, C2 => n1195, ZN => n3888);
   U4638 : AOI221_X1 port map( B1 => n14218, B2 => n2282, C1 => n14215, C2 => 
                           n2305, A => n3896, ZN => n3895);
   U4639 : OAI222_X1 port map( A1 => n14210, A2 => n1538, B1 => n7696, B2 => 
                           n14207, C1 => n14204, C2 => n1514, ZN => n3896);
   U4640 : AOI221_X1 port map( B1 => n14272, B2 => n2044, C1 => n7533, C2 => 
                           n14269, A => n3925, ZN => n3924);
   U4641 : OAI222_X1 port map( A1 => n14264, A2 => n1218, B1 => n14261, B2 => 
                           n1266, C1 => n14258, C2 => n1194, ZN => n3925);
   U4642 : AOI221_X1 port map( B1 => n14218, B2 => n2281, C1 => n14213, C2 => 
                           n2304, A => n3933, ZN => n3932);
   U4643 : OAI222_X1 port map( A1 => n14210, A2 => n1537, B1 => n7692, B2 => 
                           n14207, C1 => n14204, C2 => n1513, ZN => n3933);
   U4644 : AOI221_X1 port map( B1 => n14272, B2 => n2043, C1 => n7535, C2 => 
                           n14269, A => n5247, ZN => n5246);
   U4645 : OAI222_X1 port map( A1 => n14264, A2 => n1217, B1 => n14261, B2 => 
                           n1265, C1 => n14258, C2 => n1193, ZN => n5247);
   U4646 : AOI221_X1 port map( B1 => n14218, B2 => n2280, C1 => n831, C2 => 
                           n14213, A => n5255, ZN => n5254);
   U4647 : OAI222_X1 port map( A1 => n14210, A2 => n1536, B1 => n7688, B2 => 
                           n14207, C1 => n14204, C2 => n1512, ZN => n5255);
   U4648 : OAI222_X1 port map( A1 => n2590, A2 => n14085, B1 => n5176, B2 => 
                           n14082, C1 => n14078, C2 => n2181, ZN => n9135);
   U4649 : NOR4_X1 port map( A1 => n5177, A2 => n5178, A3 => n5179, A4 => n5180
                           , ZN => n5176);
   U4650 : NAND4_X1 port map( A1 => n5220, A2 => n5221, A3 => n5222, A4 => 
                           n5223, ZN => n5177);
   U4651 : NAND4_X1 port map( A1 => n5210, A2 => n5211, A3 => n5212, A4 => 
                           n5213, ZN => n5178);
   U4652 : OAI222_X1 port map( A1 => n2600, A2 => n14085, B1 => n4806, B2 => 
                           n14082, C1 => n14077, C2 => n2171, ZN => n9145);
   U4653 : NOR4_X1 port map( A1 => n4807, A2 => n4808, A3 => n4809, A4 => n4810
                           , ZN => n4806);
   U4654 : NAND4_X1 port map( A1 => n4835, A2 => n4836, A3 => n4837, A4 => 
                           n4838, ZN => n4807);
   U4655 : NAND4_X1 port map( A1 => n4827, A2 => n4828, A3 => n4829, A4 => 
                           n4830, ZN => n4808);
   U4656 : OAI222_X1 port map( A1 => n2599, A2 => n14085, B1 => n4843, B2 => 
                           n14082, C1 => n14077, C2 => n2172, ZN => n9144);
   U4657 : NOR4_X1 port map( A1 => n4844, A2 => n4845, A3 => n4846, A4 => n4847
                           , ZN => n4843);
   U4658 : NAND4_X1 port map( A1 => n4872, A2 => n4873, A3 => n4874, A4 => 
                           n4875, ZN => n4844);
   U4659 : NAND4_X1 port map( A1 => n4864, A2 => n4865, A3 => n4866, A4 => 
                           n4867, ZN => n4845);
   U4660 : OAI222_X1 port map( A1 => n2598, A2 => n14085, B1 => n4880, B2 => 
                           n14082, C1 => n14077, C2 => n2173, ZN => n9143);
   U4661 : NOR4_X1 port map( A1 => n4881, A2 => n4882, A3 => n4883, A4 => n4884
                           , ZN => n4880);
   U4662 : NAND4_X1 port map( A1 => n4909, A2 => n4910, A3 => n4911, A4 => 
                           n4912, ZN => n4881);
   U4663 : NAND4_X1 port map( A1 => n4901, A2 => n4902, A3 => n4903, A4 => 
                           n4904, ZN => n4882);
   U4664 : OAI222_X1 port map( A1 => n2597, A2 => n14085, B1 => n4917, B2 => 
                           n14082, C1 => n14078, C2 => n2174, ZN => n9142);
   U4665 : NOR4_X1 port map( A1 => n4918, A2 => n4919, A3 => n4920, A4 => n4921
                           , ZN => n4917);
   U4666 : NAND4_X1 port map( A1 => n4946, A2 => n4947, A3 => n4948, A4 => 
                           n4949, ZN => n4918);
   U4667 : NAND4_X1 port map( A1 => n4938, A2 => n4939, A3 => n4940, A4 => 
                           n4941, ZN => n4919);
   U4668 : OAI222_X1 port map( A1 => n2596, A2 => n14085, B1 => n4954, B2 => 
                           n14082, C1 => n14078, C2 => n2175, ZN => n9141);
   U4669 : NOR4_X1 port map( A1 => n4955, A2 => n4956, A3 => n4957, A4 => n4958
                           , ZN => n4954);
   U4670 : NAND4_X1 port map( A1 => n4983, A2 => n4984, A3 => n4985, A4 => 
                           n4986, ZN => n4955);
   U4671 : NAND4_X1 port map( A1 => n4975, A2 => n4976, A3 => n4977, A4 => 
                           n4978, ZN => n4956);
   U4672 : OAI222_X1 port map( A1 => n2595, A2 => n14085, B1 => n4991, B2 => 
                           n14082, C1 => n14078, C2 => n2176, ZN => n9140);
   U4673 : NOR4_X1 port map( A1 => n4992, A2 => n4993, A3 => n4994, A4 => n4995
                           , ZN => n4991);
   U4674 : NAND4_X1 port map( A1 => n5020, A2 => n5021, A3 => n5022, A4 => 
                           n5023, ZN => n4992);
   U4675 : NAND4_X1 port map( A1 => n5012, A2 => n5013, A3 => n5014, A4 => 
                           n5015, ZN => n4993);
   U4676 : OAI222_X1 port map( A1 => n2594, A2 => n14085, B1 => n5028, B2 => 
                           n14082, C1 => n14078, C2 => n2177, ZN => n9139);
   U4677 : NOR4_X1 port map( A1 => n5029, A2 => n5030, A3 => n5031, A4 => n5032
                           , ZN => n5028);
   U4678 : NAND4_X1 port map( A1 => n5057, A2 => n5058, A3 => n5059, A4 => 
                           n5060, ZN => n5029);
   U4679 : NAND4_X1 port map( A1 => n5049, A2 => n5050, A3 => n5051, A4 => 
                           n5052, ZN => n5030);
   U4680 : OAI222_X1 port map( A1 => n2593, A2 => n14085, B1 => n5065, B2 => 
                           n14082, C1 => n14078, C2 => n2178, ZN => n9138);
   U4681 : NOR4_X1 port map( A1 => n5066, A2 => n5067, A3 => n5068, A4 => n5069
                           , ZN => n5065);
   U4682 : NAND4_X1 port map( A1 => n5094, A2 => n5095, A3 => n5096, A4 => 
                           n5097, ZN => n5066);
   U4683 : NAND4_X1 port map( A1 => n5086, A2 => n5087, A3 => n5088, A4 => 
                           n5089, ZN => n5067);
   U4684 : OAI222_X1 port map( A1 => n2592, A2 => n14085, B1 => n5102, B2 => 
                           n14082, C1 => n14078, C2 => n2179, ZN => n9137);
   U4685 : NOR4_X1 port map( A1 => n5103, A2 => n5104, A3 => n5105, A4 => n5106
                           , ZN => n5102);
   U4686 : NAND4_X1 port map( A1 => n5131, A2 => n5132, A3 => n5133, A4 => 
                           n5134, ZN => n5103);
   U4687 : NAND4_X1 port map( A1 => n5123, A2 => n5124, A3 => n5125, A4 => 
                           n5126, ZN => n5104);
   U4688 : OAI222_X1 port map( A1 => n2591, A2 => n14085, B1 => n5139, B2 => 
                           n14082, C1 => n14078, C2 => n2180, ZN => n9136);
   U4689 : NOR4_X1 port map( A1 => n5140, A2 => n5141, A3 => n5142, A4 => n5143
                           , ZN => n5139);
   U4690 : NAND4_X1 port map( A1 => n5168, A2 => n5169, A3 => n5170, A4 => 
                           n5171, ZN => n5140);
   U4691 : NAND4_X1 port map( A1 => n5160, A2 => n5161, A3 => n5162, A4 => 
                           n5163, ZN => n5141);
   U4692 : OAI222_X1 port map( A1 => n2614, A2 => n14086, B1 => n4288, B2 => 
                           n14084, C1 => n14076, C2 => n2157, ZN => n9159);
   U4693 : NOR4_X1 port map( A1 => n4289, A2 => n4290, A3 => n4291, A4 => n4292
                           , ZN => n4288);
   U4694 : NAND4_X1 port map( A1 => n4317, A2 => n4318, A3 => n4319, A4 => 
                           n4320, ZN => n4289);
   U4695 : NAND4_X1 port map( A1 => n4309, A2 => n4310, A3 => n4311, A4 => 
                           n4312, ZN => n4290);
   U4696 : AOI221_X1 port map( B1 => n8482, B2 => n13952, C1 => n8450, C2 => 
                           n13947, A => n5216, ZN => n5212);
   U4697 : OAI22_X1 port map( A1 => n13946, A2 => n1376, B1 => n13943, B2 => 
                           n1352, ZN => n5216);
   U4698 : AOI221_X1 port map( B1 => n8513, B2 => n13952, C1 => n8481, C2 => 
                           n13947, A => n4026, ZN => n4016);
   U4699 : OAI22_X1 port map( A1 => n13946, A2 => n171, B1 => n13943, B2 => 
                           n163, ZN => n4026);
   U4700 : AOI221_X1 port map( B1 => n8002, B2 => n14736, C1 => n7970, C2 => 
                           n14733, A => n2865, ZN => n2861);
   U4701 : OAI22_X1 port map( A1 => n315, A2 => n14115, B1 => n14354, B2 => 
                           n323, ZN => n2865);
   U4702 : AOI221_X1 port map( B1 => n8001, B2 => n14736, C1 => n7969, C2 => 
                           n14733, A => n2912, ZN => n2909);
   U4703 : OAI22_X1 port map( A1 => n314, A2 => n14116, B1 => n14354, B2 => 
                           n322, ZN => n2912);
   U4704 : AOI221_X1 port map( B1 => n8000, B2 => n14736, C1 => n7968, C2 => 
                           n14733, A => n2949, ZN => n2946);
   U4705 : OAI22_X1 port map( A1 => n313, A2 => n14115, B1 => n14354, B2 => 
                           n321, ZN => n2949);
   U4706 : AOI221_X1 port map( B1 => n7999, B2 => n14736, C1 => n7967, C2 => 
                           n14733, A => n2986, ZN => n2983);
   U4707 : OAI22_X1 port map( A1 => n312, A2 => n14116, B1 => n14354, B2 => 
                           n320, ZN => n2986);
   U4708 : AOI221_X1 port map( B1 => n7998, B2 => n14736, C1 => n7966, C2 => 
                           n14733, A => n3023, ZN => n3020);
   U4709 : OAI22_X1 port map( A1 => n311, A2 => n14115, B1 => n14354, B2 => 
                           n319, ZN => n3023);
   U4710 : AOI221_X1 port map( B1 => n7997, B2 => n14736, C1 => n7965, C2 => 
                           n14733, A => n3060, ZN => n3057);
   U4712 : OAI22_X1 port map( A1 => n310, A2 => n14116, B1 => n14354, B2 => 
                           n318, ZN => n3060);
   U4713 : AOI221_X1 port map( B1 => n7996, B2 => n14736, C1 => n7964, C2 => 
                           n14733, A => n3097, ZN => n3094);
   U4714 : OAI22_X1 port map( A1 => n309, A2 => n14115, B1 => n14354, B2 => 
                           n317, ZN => n3097);
   U4715 : AOI221_X1 port map( B1 => n8003, B2 => n14734, C1 => n7971, C2 => 
                           n14731, A => n6600, ZN => n6597);
   U4716 : OAI22_X1 port map( A1 => n316, A2 => n14115, B1 => n14354, B2 => 
                           n324, ZN => n6600);
   U4717 : AOI221_X1 port map( B1 => n7982, B2 => n14734, C1 => n7950, C2 => 
                           n14731, A => n3617, ZN => n3614);
   U4718 : OAI22_X1 port map( A1 => n924, A2 => n14115, B1 => n14355, B2 => 
                           n518, ZN => n3617);
   U4719 : AOI221_X1 port map( B1 => n7981, B2 => n14734, C1 => n7949, C2 => 
                           n14731, A => n3654, ZN => n3651);
   U4720 : OAI22_X1 port map( A1 => n922, A2 => n14115, B1 => n14355, B2 => 
                           n517, ZN => n3654);
   U4721 : AOI221_X1 port map( B1 => n7980, B2 => n14734, C1 => n7948, C2 => 
                           n14731, A => n3691, ZN => n3688);
   U4722 : OAI22_X1 port map( A1 => n918, A2 => n14115, B1 => n14355, B2 => 
                           n516, ZN => n3691);
   U4723 : AOI221_X1 port map( B1 => n7979, B2 => n14734, C1 => n7947, C2 => 
                           n14731, A => n3728, ZN => n3725);
   U4724 : OAI22_X1 port map( A1 => n916, A2 => n14115, B1 => n14355, B2 => 
                           n515, ZN => n3728);
   U4725 : AOI221_X1 port map( B1 => n7978, B2 => n14734, C1 => n7946, C2 => 
                           n14731, A => n3765, ZN => n3762);
   U4726 : OAI22_X1 port map( A1 => n912, A2 => n14115, B1 => n14355, B2 => 
                           n514, ZN => n3765);
   U4727 : AOI221_X1 port map( B1 => n7977, B2 => n14734, C1 => n7945, C2 => 
                           n14731, A => n3802, ZN => n3799);
   U4728 : OAI22_X1 port map( A1 => n910, A2 => n14115, B1 => n14354, B2 => 
                           n513, ZN => n3802);
   U4729 : AOI221_X1 port map( B1 => n7976, B2 => n14734, C1 => n7944, C2 => 
                           n14731, A => n3839, ZN => n3836);
   U4730 : OAI22_X1 port map( A1 => n906, A2 => n14115, B1 => n14355, B2 => 
                           n512, ZN => n3839);
   U4731 : AOI221_X1 port map( B1 => n7975, B2 => n14734, C1 => n7943, C2 => 
                           n14731, A => n3876, ZN => n3873);
   U4732 : OAI22_X1 port map( A1 => n904, A2 => n14115, B1 => n14354, B2 => 
                           n511, ZN => n3876);
   U4733 : AOI221_X1 port map( B1 => n7974, B2 => n14734, C1 => n7942, C2 => 
                           n14731, A => n3913, ZN => n3910);
   U4734 : OAI22_X1 port map( A1 => n900, A2 => n14115, B1 => n14355, B2 => 
                           n510, ZN => n3913);
   U4735 : AOI221_X1 port map( B1 => n7973, B2 => n14734, C1 => n7941, C2 => 
                           n14731, A => n3950, ZN => n3947);
   U4736 : OAI22_X1 port map( A1 => n898, A2 => n14115, B1 => n14354, B2 => 
                           n509, ZN => n3950);
   U4737 : AOI221_X1 port map( B1 => n7972, B2 => n14734, C1 => n7940, C2 => 
                           n14731, A => n5272, ZN => n5269);
   U4738 : OAI22_X1 port map( A1 => n819, A2 => n14115, B1 => n14355, B2 => 
                           n508, ZN => n5272);
   U4739 : AOI221_X1 port map( B1 => n13950, B2 => n8507, C1 => n13947, C2 => 
                           n8475, A => n4277, ZN => n4274);
   U4740 : OAI22_X1 port map( A1 => n165, A2 => n13944, B1 => n157, B2 => 
                           n13941, ZN => n4277);
   U4741 : AOI221_X1 port map( B1 => n13908, B2 => n8824, C1 => n13905, C2 => 
                           n8793, A => n4285, ZN => n4282);
   U4742 : OAI22_X1 port map( A1 => n34, A2 => n13902, B1 => n26, B2 => n13899,
                           ZN => n4285);
   U4743 : AOI221_X1 port map( B1 => n13732, B2 => n8512, C1 => n13729, C2 => 
                           n8480, A => n5413, ZN => n5410);
   U4744 : OAI22_X1 port map( A1 => n170, A2 => n13726, B1 => n162, B2 => 
                           n13723, ZN => n5413);
   U4745 : AOI221_X1 port map( B1 => n13678, B2 => n8829, C1 => n13675, C2 => 
                           n8798, A => n5421, ZN => n5418);
   U4746 : OAI22_X1 port map( A1 => n39, A2 => n13672, B1 => n31, B2 => n13669,
                           ZN => n5421);
   U4747 : AOI221_X1 port map( B1 => n13732, B2 => n8510, C1 => n13729, C2 => 
                           n8478, A => n5487, ZN => n5484);
   U4748 : OAI22_X1 port map( A1 => n168, A2 => n13726, B1 => n160, B2 => 
                           n13723, ZN => n5487);
   U4749 : AOI221_X1 port map( B1 => n13678, B2 => n8827, C1 => n13675, C2 => 
                           n8796, A => n5495, ZN => n5492);
   U4750 : OAI22_X1 port map( A1 => n37, A2 => n13672, B1 => n29, B2 => n13669,
                           ZN => n5495);
   U4751 : AOI221_X1 port map( B1 => n13732, B2 => n8509, C1 => n13729, C2 => 
                           n8477, A => n5524, ZN => n5521);
   U4752 : OAI22_X1 port map( A1 => n167, A2 => n13726, B1 => n159, B2 => 
                           n13723, ZN => n5524);
   U4753 : AOI221_X1 port map( B1 => n13678, B2 => n8826, C1 => n13675, C2 => 
                           n8795, A => n5532, ZN => n5529);
   U4754 : OAI22_X1 port map( A1 => n36, A2 => n13672, B1 => n28, B2 => n13669,
                           ZN => n5532);
   U4755 : AOI221_X1 port map( B1 => n13732, B2 => n8508, C1 => n13729, C2 => 
                           n8476, A => n5561, ZN => n5558);
   U4756 : OAI22_X1 port map( A1 => n166, A2 => n13726, B1 => n158, B2 => 
                           n13723, ZN => n5561);
   U4757 : AOI221_X1 port map( B1 => n13678, B2 => n8825, C1 => n13675, C2 => 
                           n8794, A => n5569, ZN => n5566);
   U4758 : OAI22_X1 port map( A1 => n35, A2 => n13672, B1 => n27, B2 => n13669,
                           ZN => n5569);
   U4759 : AOI221_X1 port map( B1 => n13732, B2 => n8507, C1 => n13729, C2 => 
                           n8475, A => n5598, ZN => n5595);
   U4760 : OAI22_X1 port map( A1 => n165, A2 => n13726, B1 => n157, B2 => 
                           n13723, ZN => n5598);
   U4761 : AOI221_X1 port map( B1 => n13678, B2 => n8824, C1 => n13675, C2 => 
                           n8793, A => n5606, ZN => n5603);
   U4762 : OAI22_X1 port map( A1 => n34, A2 => n13672, B1 => n26, B2 => n13669,
                           ZN => n5606);
   U4763 : AOI221_X1 port map( B1 => n13951, B2 => n8493, C1 => n13948, C2 => 
                           n8461, A => n4795, ZN => n4792);
   U4764 : OAI22_X1 port map( A1 => n1387, A2 => n13945, B1 => n1363, B2 => 
                           n13942, ZN => n4795);
   U4765 : AOI221_X1 port map( B1 => n13909, B2 => n8810, C1 => n13906, C2 => 
                           n8779, A => n4803, ZN => n4800);
   U4766 : OAI22_X1 port map( A1 => n721, A2 => n13903, B1 => n795, B2 => 
                           n13900, ZN => n4803);
   U4767 : AOI221_X1 port map( B1 => n13951, B2 => n8492, C1 => n13948, C2 => 
                           n8460, A => n4832, ZN => n4829);
   U4768 : OAI22_X1 port map( A1 => n1386, A2 => n13945, B1 => n1362, B2 => 
                           n13942, ZN => n4832);
   U4769 : AOI221_X1 port map( B1 => n13909, B2 => n8809, C1 => n13906, C2 => 
                           n8778, A => n4840, ZN => n4837);
   U4770 : OAI22_X1 port map( A1 => n720, A2 => n13903, B1 => n731, B2 => 
                           n13900, ZN => n4840);
   U4771 : AOI221_X1 port map( B1 => n13951, B2 => n8491, C1 => n13948, C2 => 
                           n8459, A => n4869, ZN => n4866);
   U4772 : OAI22_X1 port map( A1 => n1385, A2 => n13945, B1 => n1361, B2 => 
                           n13942, ZN => n4869);
   U4773 : AOI221_X1 port map( B1 => n13909, B2 => n8808, C1 => n13906, C2 => 
                           n8777, A => n4877, ZN => n4874);
   U4774 : OAI22_X1 port map( A1 => n719, A2 => n13903, B1 => n695, B2 => 
                           n13900, ZN => n4877);
   U4775 : AOI221_X1 port map( B1 => n13951, B2 => n8490, C1 => n13948, C2 => 
                           n8458, A => n4906, ZN => n4903);
   U4776 : OAI22_X1 port map( A1 => n1384, A2 => n13945, B1 => n1360, B2 => 
                           n13942, ZN => n4906);
   U4777 : AOI221_X1 port map( B1 => n13909, B2 => n8807, C1 => n13906, C2 => 
                           n8776, A => n4914, ZN => n4911);
   U4778 : OAI22_X1 port map( A1 => n718, A2 => n13903, B1 => n694, B2 => 
                           n13900, ZN => n4914);
   U4779 : AOI221_X1 port map( B1 => n13951, B2 => n8489, C1 => n13949, C2 => 
                           n8457, A => n4943, ZN => n4940);
   U4780 : OAI22_X1 port map( A1 => n1383, A2 => n13945, B1 => n1359, B2 => 
                           n13942, ZN => n4943);
   U4781 : AOI221_X1 port map( B1 => n13909, B2 => n8806, C1 => n13907, C2 => 
                           n8775, A => n4951, ZN => n4948);
   U4782 : OAI22_X1 port map( A1 => n717, A2 => n13903, B1 => n693, B2 => 
                           n13900, ZN => n4951);
   U4783 : AOI221_X1 port map( B1 => n13730, B2 => n8493, C1 => n13727, C2 => 
                           n8461, A => n6116, ZN => n6113);
   U4784 : OAI22_X1 port map( A1 => n1387, A2 => n13724, B1 => n1363, B2 => 
                           n13721, ZN => n6116);
   U4785 : AOI221_X1 port map( B1 => n13676, B2 => n8810, C1 => n13673, C2 => 
                           n8779, A => n6124, ZN => n6121);
   U4786 : OAI22_X1 port map( A1 => n721, A2 => n13670, B1 => n795, B2 => 
                           n13667, ZN => n6124);
   U4787 : AOI221_X1 port map( B1 => n13730, B2 => n8492, C1 => n13727, C2 => 
                           n8460, A => n6153, ZN => n6150);
   U4788 : OAI22_X1 port map( A1 => n1386, A2 => n13724, B1 => n1362, B2 => 
                           n13721, ZN => n6153);
   U4789 : AOI221_X1 port map( B1 => n13676, B2 => n8809, C1 => n13673, C2 => 
                           n8778, A => n6161, ZN => n6158);
   U4790 : OAI22_X1 port map( A1 => n720, A2 => n13670, B1 => n731, B2 => 
                           n13667, ZN => n6161);
   U4791 : AOI221_X1 port map( B1 => n13730, B2 => n8491, C1 => n13727, C2 => 
                           n8459, A => n6190, ZN => n6187);
   U4792 : OAI22_X1 port map( A1 => n1385, A2 => n13724, B1 => n1361, B2 => 
                           n13721, ZN => n6190);
   U4793 : AOI221_X1 port map( B1 => n13676, B2 => n8808, C1 => n13673, C2 => 
                           n8777, A => n6198, ZN => n6195);
   U4794 : OAI22_X1 port map( A1 => n719, A2 => n13670, B1 => n695, B2 => 
                           n13667, ZN => n6198);
   U4795 : AOI221_X1 port map( B1 => n13730, B2 => n8490, C1 => n13727, C2 => 
                           n8458, A => n6227, ZN => n6224);
   U4796 : OAI22_X1 port map( A1 => n1384, A2 => n13724, B1 => n1360, B2 => 
                           n13721, ZN => n6227);
   U4797 : AOI221_X1 port map( B1 => n13676, B2 => n8807, C1 => n13673, C2 => 
                           n8776, A => n6235, ZN => n6232);
   U4798 : OAI22_X1 port map( A1 => n718, A2 => n13670, B1 => n694, B2 => 
                           n13667, ZN => n6235);
   U4799 : AOI221_X1 port map( B1 => n13730, B2 => n8489, C1 => n13727, C2 => 
                           n8457, A => n6264, ZN => n6261);
   U4800 : OAI22_X1 port map( A1 => n1383, A2 => n13724, B1 => n1359, B2 => 
                           n13721, ZN => n6264);
   U4801 : AOI221_X1 port map( B1 => n13676, B2 => n8806, C1 => n13673, C2 => 
                           n8775, A => n6272, ZN => n6269);
   U4802 : OAI22_X1 port map( A1 => n717, A2 => n13670, B1 => n693, B2 => 
                           n13667, ZN => n6272);
   U4803 : AOI221_X1 port map( B1 => n13730, B2 => n8488, C1 => n13727, C2 => 
                           n8456, A => n6301, ZN => n6298);
   U4804 : OAI22_X1 port map( A1 => n1382, A2 => n13724, B1 => n1358, B2 => 
                           n13721, ZN => n6301);
   U4805 : AOI221_X1 port map( B1 => n13676, B2 => n8805, C1 => n13673, C2 => 
                           n8774, A => n6309, ZN => n6306);
   U4806 : OAI22_X1 port map( A1 => n716, A2 => n13670, B1 => n692, B2 => 
                           n13667, ZN => n6309);
   U4807 : AOI221_X1 port map( B1 => n13730, B2 => n8487, C1 => n13727, C2 => 
                           n8455, A => n6338, ZN => n6335);
   U4808 : OAI22_X1 port map( A1 => n1381, A2 => n13724, B1 => n1357, B2 => 
                           n13721, ZN => n6338);
   U4809 : AOI221_X1 port map( B1 => n13676, B2 => n8804, C1 => n13673, C2 => 
                           n8773, A => n6346, ZN => n6343);
   U4810 : OAI22_X1 port map( A1 => n715, A2 => n13670, B1 => n691, B2 => 
                           n13667, ZN => n6346);
   U4811 : AOI221_X1 port map( B1 => n13730, B2 => n8486, C1 => n13727, C2 => 
                           n8454, A => n6375, ZN => n6372);
   U4812 : OAI22_X1 port map( A1 => n1380, A2 => n13724, B1 => n1356, B2 => 
                           n13721, ZN => n6375);
   U4813 : AOI221_X1 port map( B1 => n13676, B2 => n8803, C1 => n13673, C2 => 
                           n8772, A => n6383, ZN => n6380);
   U4814 : OAI22_X1 port map( A1 => n714, A2 => n13670, B1 => n690, B2 => 
                           n13667, ZN => n6383);
   U4815 : AOI221_X1 port map( B1 => n13730, B2 => n8485, C1 => n13727, C2 => 
                           n8453, A => n6412, ZN => n6409);
   U4816 : OAI22_X1 port map( A1 => n1379, A2 => n13724, B1 => n1355, B2 => 
                           n13721, ZN => n6412);
   U4817 : AOI221_X1 port map( B1 => n13676, B2 => n8802, C1 => n13673, C2 => 
                           n8771, A => n6420, ZN => n6417);
   U4818 : OAI22_X1 port map( A1 => n713, A2 => n13670, B1 => n689, B2 => 
                           n13667, ZN => n6420);
   U4819 : AOI221_X1 port map( B1 => n13730, B2 => n8484, C1 => n13727, C2 => 
                           n8452, A => n6449, ZN => n6446);
   U4820 : OAI22_X1 port map( A1 => n1378, A2 => n13724, B1 => n1354, B2 => 
                           n13721, ZN => n6449);
   U4821 : AOI221_X1 port map( B1 => n13676, B2 => n8801, C1 => n13673, C2 => 
                           n8770, A => n6457, ZN => n6454);
   U4822 : OAI22_X1 port map( A1 => n712, A2 => n13670, B1 => n688, B2 => 
                           n13667, ZN => n6457);
   U4823 : AOI221_X1 port map( B1 => n13730, B2 => n8483, C1 => n13727, C2 => 
                           n8451, A => n6486, ZN => n6483);
   U4824 : OAI22_X1 port map( A1 => n1377, A2 => n13724, B1 => n1353, B2 => 
                           n13721, ZN => n6486);
   U4825 : AOI221_X1 port map( B1 => n13676, B2 => n8800, C1 => n13673, C2 => 
                           n8769, A => n6494, ZN => n6491);
   U4826 : OAI22_X1 port map( A1 => n711, A2 => n13670, B1 => n687, B2 => 
                           n13667, ZN => n6494);
   U4827 : AOI221_X1 port map( B1 => n13951, B2 => n8495, C1 => n13948, C2 => 
                           n8463, A => n4721, ZN => n4718);
   U4828 : OAI22_X1 port map( A1 => n1389, A2 => n13945, B1 => n1365, B2 => 
                           n13942, ZN => n4721);
   U4829 : AOI221_X1 port map( B1 => n13909, B2 => n8812, C1 => n13906, C2 => 
                           n8781, A => n4729, ZN => n4726);
   U4830 : OAI22_X1 port map( A1 => n723, A2 => n13903, B1 => n699, B2 => 
                           n13900, ZN => n4729);
   U4831 : AOI221_X1 port map( B1 => n13951, B2 => n8494, C1 => n13948, C2 => 
                           n8462, A => n4758, ZN => n4755);
   U4832 : OAI22_X1 port map( A1 => n1388, A2 => n13945, B1 => n1364, B2 => 
                           n13942, ZN => n4758);
   U4833 : AOI221_X1 port map( B1 => n13909, B2 => n8811, C1 => n13906, C2 => 
                           n8780, A => n4766, ZN => n4763);
   U4834 : OAI22_X1 port map( A1 => n722, A2 => n13903, B1 => n698, B2 => 
                           n13900, ZN => n4766);
   U4835 : AOI221_X1 port map( B1 => n13731, B2 => n8495, C1 => n13728, C2 => 
                           n8463, A => n6042, ZN => n6039);
   U4836 : OAI22_X1 port map( A1 => n1389, A2 => n13725, B1 => n1365, B2 => 
                           n13722, ZN => n6042);
   U4837 : AOI221_X1 port map( B1 => n13677, B2 => n8812, C1 => n13674, C2 => 
                           n8781, A => n6050, ZN => n6047);
   U4838 : OAI22_X1 port map( A1 => n723, A2 => n13671, B1 => n699, B2 => 
                           n13668, ZN => n6050);
   U4839 : AOI221_X1 port map( B1 => n13731, B2 => n8494, C1 => n13728, C2 => 
                           n8462, A => n6079, ZN => n6076);
   U4840 : OAI22_X1 port map( A1 => n1388, A2 => n13725, B1 => n1364, B2 => 
                           n13722, ZN => n6079);
   U4841 : AOI221_X1 port map( B1 => n13677, B2 => n8811, C1 => n13674, C2 => 
                           n8780, A => n6087, ZN => n6084);
   U4842 : OAI22_X1 port map( A1 => n722, A2 => n13671, B1 => n698, B2 => 
                           n13668, ZN => n6087);
   U4843 : AOI221_X1 port map( B1 => n13730, B2 => n8482, C1 => n13727, C2 => 
                           n8450, A => n6537, ZN => n6533);
   U4844 : OAI22_X1 port map( A1 => n1376, A2 => n13724, B1 => n1352, B2 => 
                           n13721, ZN => n6537);
   U4845 : AOI221_X1 port map( B1 => n13676, B2 => n8799, C1 => n13673, C2 => 
                           n8768, A => n6546, ZN => n6543);
   U4846 : OAI22_X1 port map( A1 => n710, A2 => n13670, B1 => n686, B2 => 
                           n13667, ZN => n6546);
   U4847 : AOI221_X1 port map( B1 => n13952, B2 => n8488, C1 => n13949, C2 => 
                           n8456, A => n4980, ZN => n4977);
   U4848 : OAI22_X1 port map( A1 => n1382, A2 => n13946, B1 => n1358, B2 => 
                           n13943, ZN => n4980);
   U4849 : AOI221_X1 port map( B1 => n13910, B2 => n8805, C1 => n13907, C2 => 
                           n8774, A => n4988, ZN => n4985);
   U4850 : OAI22_X1 port map( A1 => n716, A2 => n13904, B1 => n692, B2 => 
                           n13901, ZN => n4988);
   U4851 : AOI221_X1 port map( B1 => n13952, B2 => n8487, C1 => n13949, C2 => 
                           n8455, A => n5017, ZN => n5014);
   U4852 : OAI22_X1 port map( A1 => n1381, A2 => n13946, B1 => n1357, B2 => 
                           n13943, ZN => n5017);
   U4853 : AOI221_X1 port map( B1 => n13910, B2 => n8804, C1 => n13907, C2 => 
                           n8773, A => n5025, ZN => n5022);
   U4854 : OAI22_X1 port map( A1 => n715, A2 => n13904, B1 => n691, B2 => 
                           n13901, ZN => n5025);
   U4855 : AOI221_X1 port map( B1 => n13952, B2 => n8486, C1 => n13949, C2 => 
                           n8454, A => n5054, ZN => n5051);
   U4856 : OAI22_X1 port map( A1 => n1380, A2 => n13946, B1 => n1356, B2 => 
                           n13943, ZN => n5054);
   U4857 : AOI221_X1 port map( B1 => n13910, B2 => n8803, C1 => n13907, C2 => 
                           n8772, A => n5062, ZN => n5059);
   U4858 : OAI22_X1 port map( A1 => n714, A2 => n13904, B1 => n690, B2 => 
                           n13901, ZN => n5062);
   U4859 : AOI221_X1 port map( B1 => n13952, B2 => n8485, C1 => n13949, C2 => 
                           n8453, A => n5091, ZN => n5088);
   U4860 : OAI22_X1 port map( A1 => n1379, A2 => n13946, B1 => n1355, B2 => 
                           n13943, ZN => n5091);
   U4861 : AOI221_X1 port map( B1 => n13910, B2 => n8802, C1 => n13907, C2 => 
                           n8771, A => n5099, ZN => n5096);
   U4862 : OAI22_X1 port map( A1 => n713, A2 => n13904, B1 => n689, B2 => 
                           n13901, ZN => n5099);
   U4863 : AOI221_X1 port map( B1 => n13952, B2 => n8484, C1 => n13949, C2 => 
                           n8452, A => n5128, ZN => n5125);
   U4864 : OAI22_X1 port map( A1 => n1378, A2 => n13946, B1 => n1354, B2 => 
                           n13943, ZN => n5128);
   U4865 : AOI221_X1 port map( B1 => n13910, B2 => n8801, C1 => n13907, C2 => 
                           n8770, A => n5136, ZN => n5133);
   U4866 : OAI22_X1 port map( A1 => n712, A2 => n13904, B1 => n688, B2 => 
                           n13901, ZN => n5136);
   U4867 : AOI221_X1 port map( B1 => n13952, B2 => n8483, C1 => n13947, C2 => 
                           n8451, A => n5165, ZN => n5162);
   U4868 : OAI22_X1 port map( A1 => n1377, A2 => n13946, B1 => n1353, B2 => 
                           n13943, ZN => n5165);
   U4869 : AOI221_X1 port map( B1 => n13910, B2 => n8800, C1 => n13905, C2 => 
                           n8769, A => n5173, ZN => n5170);
   U4870 : OAI22_X1 port map( A1 => n711, A2 => n13904, B1 => n687, B2 => 
                           n13901, ZN => n5173);
   U4871 : AOI221_X1 port map( B1 => n13732, B2 => n8513, C1 => n13729, C2 => 
                           n8481, A => n5347, ZN => n5337);
   U4872 : OAI22_X1 port map( A1 => n171, A2 => n13726, B1 => n163, B2 => 
                           n13723, ZN => n5347);
   U4873 : AOI221_X1 port map( B1 => n13678, B2 => n8894, C1 => n13675, C2 => 
                           n8895, A => n5373, ZN => n5363);
   U4874 : OAI22_X1 port map( A1 => n40, A2 => n13672, B1 => n32, B2 => n13669,
                           ZN => n5373);
   U4875 : AOI221_X1 port map( B1 => n13950, B2 => n8512, C1 => n13947, C2 => 
                           n8480, A => n4090, ZN => n4087);
   U4876 : OAI22_X1 port map( A1 => n170, A2 => n13944, B1 => n162, B2 => 
                           n13941, ZN => n4090);
   U4877 : AOI221_X1 port map( B1 => n13908, B2 => n8829, C1 => n13905, C2 => 
                           n8798, A => n4100, ZN => n4097);
   U4878 : OAI22_X1 port map( A1 => n39, A2 => n13902, B1 => n31, B2 => n13899,
                           ZN => n4100);
   U4879 : AOI221_X1 port map( B1 => n13950, B2 => n8511, C1 => n13947, C2 => 
                           n8479, A => n4129, ZN => n4126);
   U4880 : OAI22_X1 port map( A1 => n169, A2 => n13944, B1 => n161, B2 => 
                           n13941, ZN => n4129);
   U4881 : AOI221_X1 port map( B1 => n13908, B2 => n8828, C1 => n13905, C2 => 
                           n8797, A => n4137, ZN => n4134);
   U4882 : OAI22_X1 port map( A1 => n38, A2 => n13902, B1 => n30, B2 => n13899,
                           ZN => n4137);
   U4883 : AOI221_X1 port map( B1 => n13732, B2 => n8511, C1 => n13729, C2 => 
                           n8479, A => n5450, ZN => n5447);
   U4884 : OAI22_X1 port map( A1 => n169, A2 => n13726, B1 => n161, B2 => 
                           n13723, ZN => n5450);
   U4885 : AOI221_X1 port map( B1 => n13678, B2 => n8828, C1 => n13675, C2 => 
                           n8797, A => n5458, ZN => n5455);
   U4886 : OAI22_X1 port map( A1 => n38, A2 => n13672, B1 => n30, B2 => n13669,
                           ZN => n5458);
   U4887 : AOI221_X1 port map( B1 => n13950, B2 => n8510, C1 => n13947, C2 => 
                           n8478, A => n4166, ZN => n4163);
   U4888 : OAI22_X1 port map( A1 => n168, A2 => n13944, B1 => n160, B2 => 
                           n13941, ZN => n4166);
   U4889 : AOI221_X1 port map( B1 => n13908, B2 => n8827, C1 => n13905, C2 => 
                           n8796, A => n4174, ZN => n4171);
   U4890 : OAI22_X1 port map( A1 => n37, A2 => n13902, B1 => n29, B2 => n13899,
                           ZN => n4174);
   U4891 : AOI221_X1 port map( B1 => n13950, B2 => n8509, C1 => n13947, C2 => 
                           n8477, A => n4203, ZN => n4200);
   U4892 : OAI22_X1 port map( A1 => n167, A2 => n13944, B1 => n159, B2 => 
                           n13941, ZN => n4203);
   U4893 : AOI221_X1 port map( B1 => n13908, B2 => n8826, C1 => n13905, C2 => 
                           n8795, A => n4211, ZN => n4208);
   U4894 : OAI22_X1 port map( A1 => n36, A2 => n13902, B1 => n28, B2 => n13899,
                           ZN => n4211);
   U4895 : AOI221_X1 port map( B1 => n13950, B2 => n8508, C1 => n13947, C2 => 
                           n8476, A => n4240, ZN => n4237);
   U4896 : OAI22_X1 port map( A1 => n166, A2 => n13944, B1 => n158, B2 => 
                           n13941, ZN => n4240);
   U4897 : AOI221_X1 port map( B1 => n13908, B2 => n8825, C1 => n13905, C2 => 
                           n8794, A => n4248, ZN => n4245);
   U4898 : OAI22_X1 port map( A1 => n35, A2 => n13902, B1 => n27, B2 => n13899,
                           ZN => n4248);
   U4899 : AOI221_X1 port map( B1 => n13950, B2 => n8506, C1 => n13947, C2 => 
                           n8474, A => n4314, ZN => n4311);
   U4900 : OAI22_X1 port map( A1 => n164, A2 => n13944, B1 => n156, B2 => 
                           n13941, ZN => n4314);
   U4901 : AOI221_X1 port map( B1 => n13908, B2 => n8823, C1 => n13905, C2 => 
                           n8792, A => n4322, ZN => n4319);
   U4902 : OAI22_X1 port map( A1 => n33, A2 => n13902, B1 => n25, B2 => n13899,
                           ZN => n4322);
   U4903 : AOI221_X1 port map( B1 => n13732, B2 => n8506, C1 => n13729, C2 => 
                           n8474, A => n5635, ZN => n5632);
   U4904 : OAI22_X1 port map( A1 => n164, A2 => n13726, B1 => n156, B2 => 
                           n13723, ZN => n5635);
   U4905 : AOI221_X1 port map( B1 => n13678, B2 => n8823, C1 => n13675, C2 => 
                           n8792, A => n5643, ZN => n5640);
   U4906 : OAI22_X1 port map( A1 => n33, A2 => n13672, B1 => n25, B2 => n13669,
                           ZN => n5643);
   U4907 : AOI221_X1 port map( B1 => n13951, B2 => n8505, C1 => n13948, C2 => 
                           n8473, A => n4351, ZN => n4348);
   U4908 : OAI22_X1 port map( A1 => n1399, A2 => n13945, B1 => n1375, B2 => 
                           n13942, ZN => n4351);
   U4909 : AOI221_X1 port map( B1 => n13909, B2 => n8822, C1 => n13906, C2 => 
                           n8791, A => n4359, ZN => n4356);
   U4910 : OAI22_X1 port map( A1 => n738, A2 => n13903, B1 => n709, B2 => 
                           n13900, ZN => n4359);
   U4911 : AOI221_X1 port map( B1 => n13731, B2 => n8505, C1 => n13728, C2 => 
                           n8473, A => n5672, ZN => n5669);
   U4912 : OAI22_X1 port map( A1 => n1399, A2 => n13725, B1 => n1375, B2 => 
                           n13722, ZN => n5672);
   U4913 : AOI221_X1 port map( B1 => n13677, B2 => n8822, C1 => n13674, C2 => 
                           n8791, A => n5680, ZN => n5677);
   U4914 : OAI22_X1 port map( A1 => n738, A2 => n13671, B1 => n709, B2 => 
                           n13668, ZN => n5680);
   U4915 : AOI221_X1 port map( B1 => n7995, B2 => n14735, C1 => n7963, C2 => 
                           n14732, A => n3134, ZN => n3131);
   U4916 : OAI22_X1 port map( A1 => n964, A2 => n14116, B1 => n14354, B2 => 
                           n531, ZN => n3134);
   U4917 : AOI221_X1 port map( B1 => n13950, B2 => n8504, C1 => n13947, C2 => 
                           n8472, A => n4388, ZN => n4385);
   U4918 : OAI22_X1 port map( A1 => n1398, A2 => n13944, B1 => n1374, B2 => 
                           n13941, ZN => n4388);
   U4919 : AOI221_X1 port map( B1 => n13908, B2 => n8821, C1 => n13905, C2 => 
                           n8790, A => n4396, ZN => n4393);
   U4920 : OAI22_X1 port map( A1 => n737, A2 => n13902, B1 => n708, B2 => 
                           n13899, ZN => n4396);
   U4921 : AOI221_X1 port map( B1 => n13731, B2 => n8504, C1 => n13728, C2 => 
                           n8472, A => n5709, ZN => n5706);
   U4922 : OAI22_X1 port map( A1 => n1398, A2 => n13725, B1 => n1374, B2 => 
                           n13722, ZN => n5709);
   U4923 : AOI221_X1 port map( B1 => n13677, B2 => n8821, C1 => n13674, C2 => 
                           n8790, A => n5717, ZN => n5714);
   U4924 : OAI22_X1 port map( A1 => n737, A2 => n13671, B1 => n708, B2 => 
                           n13668, ZN => n5717);
   U4925 : AOI221_X1 port map( B1 => n7994, B2 => n14735, C1 => n7962, C2 => 
                           n14732, A => n3171, ZN => n3168);
   U4926 : OAI22_X1 port map( A1 => n960, A2 => n14116, B1 => n14354, B2 => 
                           n530, ZN => n3171);
   U4927 : AOI221_X1 port map( B1 => n13950, B2 => n8503, C1 => n13947, C2 => 
                           n8471, A => n4425, ZN => n4422);
   U4928 : OAI22_X1 port map( A1 => n1397, A2 => n13944, B1 => n1373, B2 => 
                           n13941, ZN => n4425);
   U4929 : AOI221_X1 port map( B1 => n13908, B2 => n8820, C1 => n13905, C2 => 
                           n8789, A => n4433, ZN => n4430);
   U4930 : OAI22_X1 port map( A1 => n733, A2 => n13902, B1 => n707, B2 => 
                           n13899, ZN => n4433);
   U4931 : AOI221_X1 port map( B1 => n13731, B2 => n8503, C1 => n13728, C2 => 
                           n8471, A => n5746, ZN => n5743);
   U4932 : OAI22_X1 port map( A1 => n1397, A2 => n13725, B1 => n1373, B2 => 
                           n13722, ZN => n5746);
   U4933 : AOI221_X1 port map( B1 => n13677, B2 => n8820, C1 => n13674, C2 => 
                           n8789, A => n5754, ZN => n5751);
   U4934 : OAI22_X1 port map( A1 => n733, A2 => n13671, B1 => n707, B2 => 
                           n13668, ZN => n5754);
   U4935 : AOI221_X1 port map( B1 => n7993, B2 => n14735, C1 => n7961, C2 => 
                           n14732, A => n3208, ZN => n3205);
   U4936 : OAI22_X1 port map( A1 => n958, A2 => n14116, B1 => n14354, B2 => 
                           n529, ZN => n3208);
   U4937 : AOI221_X1 port map( B1 => n13950, B2 => n8502, C1 => n13947, C2 => 
                           n8470, A => n4462, ZN => n4459);
   U4938 : OAI22_X1 port map( A1 => n1396, A2 => n13944, B1 => n1372, B2 => 
                           n13941, ZN => n4462);
   U4939 : AOI221_X1 port map( B1 => n13908, B2 => n8819, C1 => n13905, C2 => 
                           n8788, A => n4470, ZN => n4467);
   U4940 : OAI22_X1 port map( A1 => n732, A2 => n13902, B1 => n706, B2 => 
                           n13899, ZN => n4470);
   U4941 : AOI221_X1 port map( B1 => n13731, B2 => n8502, C1 => n13728, C2 => 
                           n8470, A => n5783, ZN => n5780);
   U4942 : OAI22_X1 port map( A1 => n1396, A2 => n13725, B1 => n1372, B2 => 
                           n13722, ZN => n5783);
   U4943 : AOI221_X1 port map( B1 => n13677, B2 => n8819, C1 => n13674, C2 => 
                           n8788, A => n5791, ZN => n5788);
   U4944 : OAI22_X1 port map( A1 => n732, A2 => n13671, B1 => n706, B2 => 
                           n13668, ZN => n5791);
   U4945 : AOI221_X1 port map( B1 => n7992, B2 => n14735, C1 => n7960, C2 => 
                           n14732, A => n3245, ZN => n3242);
   U4946 : OAI22_X1 port map( A1 => n954, A2 => n14116, B1 => n14354, B2 => 
                           n528, ZN => n3245);
   U4947 : AOI221_X1 port map( B1 => n13950, B2 => n8501, C1 => n13948, C2 => 
                           n8469, A => n4499, ZN => n4496);
   U4948 : OAI22_X1 port map( A1 => n1395, A2 => n13944, B1 => n1371, B2 => 
                           n13941, ZN => n4499);
   U4949 : AOI221_X1 port map( B1 => n13908, B2 => n8818, C1 => n13906, C2 => 
                           n8787, A => n4507, ZN => n4504);
   U4950 : OAI22_X1 port map( A1 => n730, A2 => n13902, B1 => n705, B2 => 
                           n13899, ZN => n4507);
   U4951 : AOI221_X1 port map( B1 => n13731, B2 => n8501, C1 => n13728, C2 => 
                           n8469, A => n5820, ZN => n5817);
   U4952 : OAI22_X1 port map( A1 => n1395, A2 => n13725, B1 => n1371, B2 => 
                           n13722, ZN => n5820);
   U4953 : AOI221_X1 port map( B1 => n13677, B2 => n8818, C1 => n13674, C2 => 
                           n8787, A => n5828, ZN => n5825);
   U4954 : OAI22_X1 port map( A1 => n730, A2 => n13671, B1 => n705, B2 => 
                           n13668, ZN => n5828);
   U4955 : AOI221_X1 port map( B1 => n7991, B2 => n14735, C1 => n7959, C2 => 
                           n14732, A => n3282, ZN => n3279);
   U4956 : OAI22_X1 port map( A1 => n952, A2 => n14116, B1 => n14355, B2 => 
                           n527, ZN => n3282);
   U4957 : AOI221_X1 port map( B1 => n13950, B2 => n8500, C1 => n13948, C2 => 
                           n8468, A => n4536, ZN => n4533);
   U4958 : OAI22_X1 port map( A1 => n1394, A2 => n13944, B1 => n1370, B2 => 
                           n13941, ZN => n4536);
   U4959 : AOI221_X1 port map( B1 => n13908, B2 => n8817, C1 => n13906, C2 => 
                           n8786, A => n4544, ZN => n4541);
   U4960 : OAI22_X1 port map( A1 => n729, A2 => n13902, B1 => n704, B2 => 
                           n13899, ZN => n4544);
   U4961 : AOI221_X1 port map( B1 => n13731, B2 => n8500, C1 => n13728, C2 => 
                           n8468, A => n5857, ZN => n5854);
   U4962 : OAI22_X1 port map( A1 => n1394, A2 => n13725, B1 => n1370, B2 => 
                           n13722, ZN => n5857);
   U4963 : AOI221_X1 port map( B1 => n13677, B2 => n8817, C1 => n13674, C2 => 
                           n8786, A => n5865, ZN => n5862);
   U4964 : OAI22_X1 port map( A1 => n729, A2 => n13671, B1 => n704, B2 => 
                           n13668, ZN => n5865);
   U4965 : AOI221_X1 port map( B1 => n7990, B2 => n14735, C1 => n7958, C2 => 
                           n14732, A => n3321, ZN => n3318);
   U4966 : OAI22_X1 port map( A1 => n948, A2 => n14116, B1 => n14355, B2 => 
                           n526, ZN => n3321);
   U4967 : AOI221_X1 port map( B1 => n13951, B2 => n8499, C1 => n13948, C2 => 
                           n8467, A => n4573, ZN => n4570);
   U4968 : OAI22_X1 port map( A1 => n1393, A2 => n13945, B1 => n1369, B2 => 
                           n13942, ZN => n4573);
   U4969 : AOI221_X1 port map( B1 => n13909, B2 => n8816, C1 => n13906, C2 => 
                           n8785, A => n4581, ZN => n4578);
   U4970 : OAI22_X1 port map( A1 => n728, A2 => n13903, B1 => n703, B2 => 
                           n13900, ZN => n4581);
   U4971 : AOI221_X1 port map( B1 => n13731, B2 => n8499, C1 => n13728, C2 => 
                           n8467, A => n5894, ZN => n5891);
   U4972 : OAI22_X1 port map( A1 => n1393, A2 => n13725, B1 => n1369, B2 => 
                           n13722, ZN => n5894);
   U4973 : AOI221_X1 port map( B1 => n13677, B2 => n8816, C1 => n13674, C2 => 
                           n8785, A => n5902, ZN => n5899);
   U4974 : OAI22_X1 port map( A1 => n728, A2 => n13671, B1 => n703, B2 => 
                           n13668, ZN => n5902);
   U4975 : AOI221_X1 port map( B1 => n7989, B2 => n14735, C1 => n7957, C2 => 
                           n14732, A => n3358, ZN => n3355);
   U4976 : OAI22_X1 port map( A1 => n946, A2 => n14116, B1 => n14355, B2 => 
                           n525, ZN => n3358);
   U4977 : AOI221_X1 port map( B1 => n13951, B2 => n8498, C1 => n13948, C2 => 
                           n8466, A => n4610, ZN => n4607);
   U4978 : OAI22_X1 port map( A1 => n1392, A2 => n13945, B1 => n1368, B2 => 
                           n13942, ZN => n4610);
   U4979 : AOI221_X1 port map( B1 => n13909, B2 => n8815, C1 => n13906, C2 => 
                           n8784, A => n4618, ZN => n4615);
   U4980 : OAI22_X1 port map( A1 => n726, A2 => n13903, B1 => n702, B2 => 
                           n13900, ZN => n4618);
   U4981 : AOI221_X1 port map( B1 => n13731, B2 => n8498, C1 => n13728, C2 => 
                           n8466, A => n5931, ZN => n5928);
   U4982 : OAI22_X1 port map( A1 => n1392, A2 => n13725, B1 => n1368, B2 => 
                           n13722, ZN => n5931);
   U4983 : AOI221_X1 port map( B1 => n13677, B2 => n8815, C1 => n13674, C2 => 
                           n8784, A => n5939, ZN => n5936);
   U4984 : OAI22_X1 port map( A1 => n726, A2 => n13671, B1 => n702, B2 => 
                           n13668, ZN => n5939);
   U4985 : AOI221_X1 port map( B1 => n7988, B2 => n14735, C1 => n7956, C2 => 
                           n14732, A => n3395, ZN => n3392);
   U4986 : OAI22_X1 port map( A1 => n942, A2 => n14116, B1 => n14355, B2 => 
                           n524, ZN => n3395);
   U4987 : AOI221_X1 port map( B1 => n13951, B2 => n8497, C1 => n13948, C2 => 
                           n8465, A => n4647, ZN => n4644);
   U4988 : OAI22_X1 port map( A1 => n1391, A2 => n13945, B1 => n1367, B2 => 
                           n13942, ZN => n4647);
   U4989 : AOI221_X1 port map( B1 => n13909, B2 => n8814, C1 => n13906, C2 => 
                           n8783, A => n4655, ZN => n4652);
   U4990 : OAI22_X1 port map( A1 => n725, A2 => n13903, B1 => n701, B2 => 
                           n13900, ZN => n4655);
   U4991 : AOI221_X1 port map( B1 => n13731, B2 => n8497, C1 => n13728, C2 => 
                           n8465, A => n5968, ZN => n5965);
   U4992 : OAI22_X1 port map( A1 => n1391, A2 => n13725, B1 => n1367, B2 => 
                           n13722, ZN => n5968);
   U4993 : AOI221_X1 port map( B1 => n13677, B2 => n8814, C1 => n13674, C2 => 
                           n8783, A => n5976, ZN => n5973);
   U4994 : OAI22_X1 port map( A1 => n725, A2 => n13671, B1 => n701, B2 => 
                           n13668, ZN => n5976);
   U4995 : AOI221_X1 port map( B1 => n7987, B2 => n14735, C1 => n7955, C2 => 
                           n14732, A => n3432, ZN => n3429);
   U4996 : OAI22_X1 port map( A1 => n940, A2 => n14116, B1 => n14355, B2 => 
                           n523, ZN => n3432);
   U4997 : AOI221_X1 port map( B1 => n13951, B2 => n8496, C1 => n13948, C2 => 
                           n8464, A => n4684, ZN => n4681);
   U4998 : OAI22_X1 port map( A1 => n1390, A2 => n13945, B1 => n1366, B2 => 
                           n13942, ZN => n4684);
   U4999 : AOI221_X1 port map( B1 => n13909, B2 => n8813, C1 => n13906, C2 => 
                           n8782, A => n4692, ZN => n4689);
   U5000 : OAI22_X1 port map( A1 => n724, A2 => n13903, B1 => n700, B2 => 
                           n13900, ZN => n4692);
   U5001 : AOI221_X1 port map( B1 => n13731, B2 => n8496, C1 => n13728, C2 => 
                           n8464, A => n6005, ZN => n6002);
   U5002 : OAI22_X1 port map( A1 => n1390, A2 => n13725, B1 => n1366, B2 => 
                           n13722, ZN => n6005);
   U5003 : AOI221_X1 port map( B1 => n13677, B2 => n8813, C1 => n13674, C2 => 
                           n8782, A => n6013, ZN => n6010);
   U5004 : OAI22_X1 port map( A1 => n724, A2 => n13671, B1 => n700, B2 => 
                           n13668, ZN => n6013);
   U5005 : AOI221_X1 port map( B1 => n7986, B2 => n14735, C1 => n7954, C2 => 
                           n14732, A => n3469, ZN => n3466);
   U5006 : OAI22_X1 port map( A1 => n936, A2 => n14116, B1 => n14355, B2 => 
                           n522, ZN => n3469);
   U5007 : AOI221_X1 port map( B1 => n7985, B2 => n14735, C1 => n7953, C2 => 
                           n14732, A => n3506, ZN => n3503);
   U5008 : OAI22_X1 port map( A1 => n934, A2 => n14116, B1 => n14355, B2 => 
                           n521, ZN => n3506);
   U5009 : AOI221_X1 port map( B1 => n7329, B2 => n13221, C1 => n13223, C2 => 
                           n7325, A => n3543, ZN => n3540);
   U5010 : OAI22_X1 port map( A1 => n805, A2 => n2761, B1 => n806, B2 => n2757,
                           ZN => n3543);
   U5011 : AOI221_X1 port map( B1 => n7983, B2 => n14735, C1 => n7951, C2 => 
                           n14732, A => n3580, ZN => n3577);
   U5012 : OAI22_X1 port map( A1 => n928, A2 => n14116, B1 => n14355, B2 => 
                           n519, ZN => n3580);
   U5013 : OAI222_X1 port map( A1 => n7437, A2 => n13229, B1 => n14715, B2 => 
                           n13228, C1 => n14761, C2 => n13232, ZN => n10031);
   U5014 : OAI222_X1 port map( A1 => n7461, A2 => n13229, B1 => n14703, B2 => 
                           n13228, C1 => n14755, C2 => n13232, ZN => n10030);
   U5015 : OAI222_X1 port map( A1 => n7438, A2 => n14717, B1 => n14715, B2 => 
                           n14709, C1 => n14761, C2 => n14704, ZN => n9999);
   U5016 : OAI222_X1 port map( A1 => n7462, A2 => n14716, B1 => n14707, B2 => 
                           n14703, C1 => n14755, C2 => n14704, ZN => n9998);
   U5017 : OAI222_X1 port map( A1 => n6742, A2 => n14716, B1 => n14707, B2 => 
                           n14682, C1 => n14935, C2 => n14704, ZN => n10028);
   U5018 : OAI222_X1 port map( A1 => n6766, A2 => n14716, B1 => n14707, B2 => 
                           n14676, C1 => n14929, C2 => n14704, ZN => n10027);
   U5019 : OAI222_X1 port map( A1 => n6790, A2 => n14716, B1 => n14707, B2 => 
                           n14670, C1 => n14923, C2 => n14704, ZN => n10026);
   U5020 : OAI222_X1 port map( A1 => n6814, A2 => n14716, B1 => n14707, B2 => 
                           n14664, C1 => n14917, C2 => n14704, ZN => n10025);
   U5021 : OAI222_X1 port map( A1 => n6838, A2 => n14716, B1 => n14708, B2 => 
                           n14658, C1 => n14911, C2 => n14704, ZN => n10024);
   U5022 : OAI222_X1 port map( A1 => n6862, A2 => n14716, B1 => n14707, B2 => 
                           n14652, C1 => n14905, C2 => n14704, ZN => n10023);
   U5023 : OAI222_X1 port map( A1 => n6886, A2 => n14716, B1 => n14707, B2 => 
                           n14646, C1 => n14899, C2 => n14704, ZN => n10022);
   U5024 : OAI222_X1 port map( A1 => n6910, A2 => n14716, B1 => n14707, B2 => 
                           n14640, C1 => n14893, C2 => n14704, ZN => n10021);
   U5025 : OAI222_X1 port map( A1 => n6934, A2 => n14716, B1 => n14707, B2 => 
                           n14634, C1 => n14887, C2 => n14704, ZN => n10020);
   U5026 : OAI222_X1 port map( A1 => n6958, A2 => n14717, B1 => n14707, B2 => 
                           n14628, C1 => n14881, C2 => n14705, ZN => n10019);
   U5027 : OAI222_X1 port map( A1 => n6982, A2 => n14717, B1 => n14708, B2 => 
                           n14622, C1 => n14875, C2 => n14705, ZN => n10018);
   U5028 : OAI222_X1 port map( A1 => n7006, A2 => n14717, B1 => n14708, B2 => 
                           n14616, C1 => n14869, C2 => n14705, ZN => n10017);
   U5029 : OAI222_X1 port map( A1 => n7030, A2 => n14717, B1 => n14708, B2 => 
                           n14610, C1 => n14863, C2 => n14705, ZN => n10016);
   U5030 : OAI222_X1 port map( A1 => n7054, A2 => n14717, B1 => n14708, B2 => 
                           n14604, C1 => n14857, C2 => n14705, ZN => n10015);
   U5031 : OAI222_X1 port map( A1 => n7078, A2 => n14717, B1 => n14708, B2 => 
                           n14598, C1 => n14851, C2 => n14705, ZN => n10014);
   U5032 : OAI222_X1 port map( A1 => n7102, A2 => n14717, B1 => n14708, B2 => 
                           n14592, C1 => n14845, C2 => n14705, ZN => n10013);
   U5033 : OAI222_X1 port map( A1 => n7126, A2 => n14717, B1 => n14708, B2 => 
                           n14586, C1 => n14839, C2 => n14705, ZN => n10012);
   U5034 : OAI222_X1 port map( A1 => n7150, A2 => n14717, B1 => n14708, B2 => 
                           n14580, C1 => n14833, C2 => n14705, ZN => n10011);
   U5035 : OAI222_X1 port map( A1 => n7174, A2 => n14717, B1 => n14708, B2 => 
                           n14574, C1 => n14827, C2 => n14705, ZN => n10010);
   U5036 : OAI222_X1 port map( A1 => n7486, A2 => n14716, B1 => n14707, B2 => 
                           n14697, C1 => n14749, C2 => n14704, ZN => n9997);
   U5037 : OAI222_X1 port map( A1 => n7246, A2 => n14717, B1 => n14709, B2 => 
                           n14556, C1 => n14809, C2 => n14706, ZN => n10007);
   U5038 : OAI222_X1 port map( A1 => n7270, A2 => n14717, B1 => n14709, B2 => 
                           n14550, C1 => n14803, C2 => n14706, ZN => n10006);
   U5039 : OAI222_X1 port map( A1 => n7294, A2 => n14718, B1 => n14709, B2 => 
                           n14544, C1 => n14797, C2 => n14706, ZN => n10005);
   U5040 : OAI222_X1 port map( A1 => n7318, A2 => n14718, B1 => n14709, B2 => 
                           n14538, C1 => n14791, C2 => n14706, ZN => n10004);
   U5041 : OAI222_X1 port map( A1 => n7342, A2 => n14718, B1 => n14709, B2 => 
                           n14532, C1 => n14785, C2 => n14706, ZN => n10003);
   U5042 : OAI222_X1 port map( A1 => n7366, A2 => n14718, B1 => n14709, B2 => 
                           n14526, C1 => n14779, C2 => n14706, ZN => n10002);
   U5043 : OAI222_X1 port map( A1 => n7390, A2 => n14718, B1 => n14709, B2 => 
                           n14520, C1 => n14773, C2 => n14706, ZN => n10001);
   U5044 : OAI222_X1 port map( A1 => n6918, A2 => n13638, B1 => n14887, B2 => 
                           n13635, C1 => n14630, C2 => n13633, ZN => n11492);
   U5045 : OAI222_X1 port map( A1 => n6726, A2 => n13639, B1 => n14935, B2 => 
                           n13636, C1 => n14678, C2 => n13633, ZN => n11500);
   U5046 : OAI222_X1 port map( A1 => n6750, A2 => n13639, B1 => n14929, B2 => 
                           n13636, C1 => n14672, C2 => n13633, ZN => n11499);
   U5047 : OAI222_X1 port map( A1 => n6774, A2 => n13639, B1 => n14923, B2 => 
                           n13636, C1 => n14666, C2 => n13633, ZN => n11498);
   U5048 : OAI222_X1 port map( A1 => n6798, A2 => n13639, B1 => n14917, B2 => 
                           n13636, C1 => n14660, C2 => n13633, ZN => n11497);
   U5049 : OAI222_X1 port map( A1 => n6822, A2 => n13639, B1 => n14911, B2 => 
                           n13636, C1 => n14654, C2 => n13633, ZN => n11496);
   U5050 : OAI222_X1 port map( A1 => n6846, A2 => n13639, B1 => n14905, B2 => 
                           n13636, C1 => n14648, C2 => n13633, ZN => n11495);
   U5051 : OAI222_X1 port map( A1 => n6870, A2 => n13639, B1 => n14899, B2 => 
                           n13636, C1 => n14642, C2 => n13633, ZN => n11494);
   U5052 : OAI222_X1 port map( A1 => n6894, A2 => n13639, B1 => n14893, B2 => 
                           n13636, C1 => n14636, C2 => n13633, ZN => n11493);
   U5053 : OAI222_X1 port map( A1 => n14887, A2 => n14453, B1 => n6936, B2 => 
                           n14450, C1 => n14629, C2 => n14448, ZN => n9764);
   U5054 : OAI222_X1 port map( A1 => n14887, A2 => n14480, B1 => n7782, B2 => 
                           n14476, C1 => n14629, C2 => n14475, ZN => n9860);
   U5055 : OAI222_X1 port map( A1 => n14887, A2 => n14489, B1 => n7783, B2 => 
                           n14485, C1 => n14629, C2 => n14484, ZN => n9892);
   U5056 : OAI222_X1 port map( A1 => n14887, A2 => n14435, B1 => n6938, B2 => 
                           n14431, C1 => n14629, C2 => n14430, ZN => n9700);
   U5057 : OAI222_X1 port map( A1 => n14892, A2 => n13296, B1 => n6932, B2 => 
                           n13293, C1 => n14634, C2 => n13291, ZN => n10276);
   U5058 : OAI222_X1 port map( A1 => n14892, A2 => n13314, B1 => n6930, B2 => 
                           n13311, C1 => n14634, C2 => n13309, ZN => n10340);
   U5059 : OAI222_X1 port map( A1 => n14892, A2 => n13341, B1 => n7780, B2 => 
                           n13338, C1 => n14633, C2 => n13336, ZN => n10436);
   U5060 : OAI222_X1 port map( A1 => n14891, A2 => n13350, B1 => n7781, B2 => 
                           n13347, C1 => n14633, C2 => n13345, ZN => n10468);
   U5061 : OAI222_X1 port map( A1 => n14891, A2 => n13377, B1 => n6929, B2 => 
                           n13374, C1 => n14633, C2 => n13372, ZN => n10564);
   U5062 : OAI222_X1 port map( A1 => n14890, A2 => n13458, B1 => n6926, B2 => 
                           n13455, C1 => n14632, C2 => n13453, ZN => n10852);
   U5063 : OAI222_X1 port map( A1 => n14890, A2 => n13476, B1 => n6924, B2 => 
                           n13473, C1 => n14632, C2 => n13471, ZN => n10916);
   U5064 : OAI222_X1 port map( A1 => n14890, A2 => n13539, B1 => n6923, B2 => 
                           n13536, C1 => n14631, C2 => n13534, ZN => n11140);
   U5065 : OAI222_X1 port map( A1 => n14889, A2 => n13620, B1 => n6920, B2 => 
                           n13617, C1 => n14631, C2 => n13615, ZN => n11428);
   U5066 : OAI222_X1 port map( A1 => n14889, A2 => n14316, B1 => n7636, B2 => 
                           n14312, C1 => n14630, C2 => n14311, ZN => n9284);
   U5067 : OAI222_X1 port map( A1 => n14888, A2 => n14399, B1 => n7634, B2 => 
                           n14395, C1 => n14630, C2 => n14394, ZN => n9572);
   U5068 : OAI222_X1 port map( A1 => n14935, A2 => n14436, B1 => n6746, B2 => 
                           n14432, C1 => n14677, C2 => n14430, ZN => n9708);
   U5069 : OAI222_X1 port map( A1 => n14929, A2 => n14436, B1 => n6770, B2 => 
                           n14431, C1 => n14671, C2 => n14430, ZN => n9707);
   U5070 : OAI222_X1 port map( A1 => n14923, A2 => n14436, B1 => n6794, B2 => 
                           n14431, C1 => n14665, C2 => n14430, ZN => n9706);
   U5071 : OAI222_X1 port map( A1 => n14917, A2 => n14436, B1 => n6818, B2 => 
                           n14431, C1 => n14659, C2 => n14430, ZN => n9705);
   U5072 : OAI222_X1 port map( A1 => n14911, A2 => n14436, B1 => n6842, B2 => 
                           n14431, C1 => n14653, C2 => n14430, ZN => n9704);
   U5073 : OAI222_X1 port map( A1 => n14905, A2 => n14436, B1 => n6866, B2 => 
                           n14431, C1 => n14647, C2 => n14430, ZN => n9703);
   U5074 : OAI222_X1 port map( A1 => n14899, A2 => n14436, B1 => n6890, B2 => 
                           n14431, C1 => n14641, C2 => n14430, ZN => n9702);
   U5075 : OAI222_X1 port map( A1 => n14893, A2 => n14436, B1 => n6914, B2 => 
                           n14431, C1 => n14635, C2 => n14430, ZN => n9701);
   U5076 : OAI222_X1 port map( A1 => n14935, A2 => n14445, B1 => n6745, B2 => 
                           n14441, C1 => n14677, C2 => n14439, ZN => n9740);
   U5077 : OAI222_X1 port map( A1 => n14935, A2 => n14454, B1 => n6744, B2 => 
                           n14450, C1 => n14677, C2 => n14448, ZN => n9772);
   U5078 : OAI222_X1 port map( A1 => n14929, A2 => n14454, B1 => n6768, B2 => 
                           n14449, C1 => n14671, C2 => n14448, ZN => n9771);
   U5079 : OAI222_X1 port map( A1 => n14923, A2 => n14454, B1 => n6792, B2 => 
                           n14450, C1 => n14665, C2 => n14448, ZN => n9770);
   U5080 : OAI222_X1 port map( A1 => n14917, A2 => n14454, B1 => n6816, B2 => 
                           n14450, C1 => n14659, C2 => n14448, ZN => n9769);
   U5081 : OAI222_X1 port map( A1 => n14911, A2 => n14454, B1 => n6840, B2 => 
                           n14449, C1 => n14653, C2 => n14448, ZN => n9768);
   U5082 : OAI222_X1 port map( A1 => n14905, A2 => n14454, B1 => n6864, B2 => 
                           n14449, C1 => n14647, C2 => n14448, ZN => n9767);
   U5083 : OAI222_X1 port map( A1 => n14899, A2 => n14454, B1 => n6888, B2 => 
                           n14450, C1 => n14641, C2 => n14448, ZN => n9766);
   U5084 : OAI222_X1 port map( A1 => n14893, A2 => n14454, B1 => n6912, B2 => 
                           n14449, C1 => n14635, C2 => n14448, ZN => n9765);
   U5085 : OAI222_X1 port map( A1 => n14935, A2 => n14481, B1 => n7814, B2 => 
                           n14477, C1 => n14677, C2 => n14475, ZN => n9868);
   U5086 : OAI222_X1 port map( A1 => n14929, A2 => n14481, B1 => n7810, B2 => 
                           n14476, C1 => n14671, C2 => n14475, ZN => n9867);
   U5087 : OAI222_X1 port map( A1 => n14923, A2 => n14481, B1 => n7806, B2 => 
                           n14476, C1 => n14665, C2 => n14475, ZN => n9866);
   U5088 : OAI222_X1 port map( A1 => n14917, A2 => n14481, B1 => n7802, B2 => 
                           n14476, C1 => n14659, C2 => n14475, ZN => n9865);
   U5089 : OAI222_X1 port map( A1 => n14911, A2 => n14481, B1 => n7798, B2 => 
                           n14476, C1 => n14653, C2 => n14475, ZN => n9864);
   U5090 : OAI222_X1 port map( A1 => n14905, A2 => n14481, B1 => n7794, B2 => 
                           n14476, C1 => n14647, C2 => n14475, ZN => n9863);
   U5091 : OAI222_X1 port map( A1 => n14899, A2 => n14481, B1 => n7790, B2 => 
                           n14476, C1 => n14641, C2 => n14475, ZN => n9862);
   U5092 : OAI222_X1 port map( A1 => n14893, A2 => n14481, B1 => n7786, B2 => 
                           n14476, C1 => n14635, C2 => n14475, ZN => n9861);
   U5093 : OAI222_X1 port map( A1 => n14935, A2 => n14490, B1 => n7815, B2 => 
                           n14486, C1 => n14677, C2 => n14484, ZN => n9900);
   U5094 : OAI222_X1 port map( A1 => n14929, A2 => n14490, B1 => n7811, B2 => 
                           n14485, C1 => n14671, C2 => n14484, ZN => n9899);
   U5095 : OAI222_X1 port map( A1 => n14923, A2 => n14490, B1 => n7807, B2 => 
                           n14485, C1 => n14665, C2 => n14484, ZN => n9898);
   U5096 : OAI222_X1 port map( A1 => n14917, A2 => n14490, B1 => n7803, B2 => 
                           n14485, C1 => n14659, C2 => n14484, ZN => n9897);
   U5097 : OAI222_X1 port map( A1 => n14911, A2 => n14490, B1 => n7799, B2 => 
                           n14485, C1 => n14653, C2 => n14484, ZN => n9896);
   U5098 : OAI222_X1 port map( A1 => n14905, A2 => n14490, B1 => n7795, B2 => 
                           n14485, C1 => n14647, C2 => n14484, ZN => n9895);
   U5099 : OAI222_X1 port map( A1 => n14899, A2 => n14490, B1 => n7791, B2 => 
                           n14485, C1 => n14641, C2 => n14484, ZN => n9894);
   U5100 : OAI222_X1 port map( A1 => n14893, A2 => n14490, B1 => n7787, B2 => 
                           n14485, C1 => n14635, C2 => n14484, ZN => n9893);
   U5101 : OAI222_X1 port map( A1 => n14937, A2 => n14317, B1 => n7684, B2 => 
                           n14313, C1 => n14678, C2 => n14311, ZN => n9292);
   U5102 : OAI222_X1 port map( A1 => n14931, A2 => n14317, B1 => n7678, B2 => 
                           n14312, C1 => n14672, C2 => n14311, ZN => n9291);
   U5103 : OAI222_X1 port map( A1 => n14925, A2 => n14317, B1 => n7672, B2 => 
                           n14312, C1 => n14666, C2 => n14311, ZN => n9290);
   U5104 : OAI222_X1 port map( A1 => n14919, A2 => n14317, B1 => n7666, B2 => 
                           n14312, C1 => n14660, C2 => n14311, ZN => n9289);
   U5105 : OAI222_X1 port map( A1 => n14913, A2 => n14317, B1 => n7660, B2 => 
                           n14312, C1 => n14654, C2 => n14311, ZN => n9288);
   U5106 : OAI222_X1 port map( A1 => n14907, A2 => n14317, B1 => n7654, B2 => 
                           n14312, C1 => n14648, C2 => n14311, ZN => n9287);
   U5107 : OAI222_X1 port map( A1 => n14901, A2 => n14317, B1 => n7648, B2 => 
                           n14312, C1 => n14642, C2 => n14311, ZN => n9286);
   U5108 : OAI222_X1 port map( A1 => n14895, A2 => n14317, B1 => n7642, B2 => 
                           n14312, C1 => n14636, C2 => n14311, ZN => n9285);
   U5109 : OAI222_X1 port map( A1 => n14936, A2 => n14400, B1 => n7682, B2 => 
                           n14396, C1 => n14678, C2 => n14394, ZN => n9580);
   U5110 : OAI222_X1 port map( A1 => n14930, A2 => n14400, B1 => n7676, B2 => 
                           n14395, C1 => n14672, C2 => n14394, ZN => n9579);
   U5111 : OAI222_X1 port map( A1 => n14924, A2 => n14400, B1 => n7670, B2 => 
                           n14395, C1 => n14666, C2 => n14394, ZN => n9578);
   U5112 : OAI222_X1 port map( A1 => n14918, A2 => n14400, B1 => n7664, B2 => 
                           n14395, C1 => n14660, C2 => n14394, ZN => n9577);
   U5113 : OAI222_X1 port map( A1 => n14912, A2 => n14400, B1 => n7658, B2 => 
                           n14395, C1 => n14654, C2 => n14394, ZN => n9576);
   U5114 : OAI222_X1 port map( A1 => n14906, A2 => n14400, B1 => n7652, B2 => 
                           n14395, C1 => n14648, C2 => n14394, ZN => n9575);
   U5115 : OAI222_X1 port map( A1 => n14900, A2 => n14400, B1 => n7646, B2 => 
                           n14395, C1 => n14642, C2 => n14394, ZN => n9574);
   U5116 : OAI222_X1 port map( A1 => n14894, A2 => n14400, B1 => n7640, B2 => 
                           n14395, C1 => n14636, C2 => n14394, ZN => n9573);
   U5117 : OAI222_X1 port map( A1 => n14940, A2 => n13297, B1 => n6740, B2 => 
                           n13294, C1 => n14682, C2 => n13291, ZN => n10284);
   U5118 : OAI222_X1 port map( A1 => n14934, A2 => n13297, B1 => n6764, B2 => 
                           n13294, C1 => n14676, C2 => n13291, ZN => n10283);
   U5119 : OAI222_X1 port map( A1 => n14928, A2 => n13297, B1 => n6788, B2 => 
                           n13294, C1 => n14670, C2 => n13291, ZN => n10282);
   U5120 : OAI222_X1 port map( A1 => n14922, A2 => n13297, B1 => n6812, B2 => 
                           n13294, C1 => n14664, C2 => n13291, ZN => n10281);
   U5121 : OAI222_X1 port map( A1 => n14916, A2 => n13297, B1 => n6836, B2 => 
                           n13294, C1 => n14658, C2 => n13291, ZN => n10280);
   U5122 : OAI222_X1 port map( A1 => n14910, A2 => n13297, B1 => n6860, B2 => 
                           n13294, C1 => n14652, C2 => n13291, ZN => n10279);
   U5123 : OAI222_X1 port map( A1 => n14904, A2 => n13297, B1 => n6884, B2 => 
                           n13294, C1 => n14646, C2 => n13291, ZN => n10278);
   U5124 : OAI222_X1 port map( A1 => n14898, A2 => n13297, B1 => n6908, B2 => 
                           n13294, C1 => n14640, C2 => n13291, ZN => n10277);
   U5125 : OAI222_X1 port map( A1 => n14934, A2 => n13315, B1 => n6762, B2 => 
                           n13312, C1 => n14676, C2 => n13309, ZN => n10347);
   U5126 : OAI222_X1 port map( A1 => n14928, A2 => n13315, B1 => n6786, B2 => 
                           n13312, C1 => n14670, C2 => n13309, ZN => n10346);
   U5127 : OAI222_X1 port map( A1 => n14922, A2 => n13315, B1 => n6810, B2 => 
                           n13312, C1 => n14664, C2 => n13309, ZN => n10345);
   U5128 : OAI222_X1 port map( A1 => n14916, A2 => n13315, B1 => n6834, B2 => 
                           n13312, C1 => n14658, C2 => n13309, ZN => n10344);
   U5129 : OAI222_X1 port map( A1 => n14910, A2 => n13315, B1 => n6858, B2 => 
                           n13312, C1 => n14652, C2 => n13309, ZN => n10343);
   U5130 : OAI222_X1 port map( A1 => n14904, A2 => n13315, B1 => n6882, B2 => 
                           n13312, C1 => n14646, C2 => n13309, ZN => n10342);
   U5131 : OAI222_X1 port map( A1 => n14898, A2 => n13315, B1 => n6906, B2 => 
                           n13312, C1 => n14640, C2 => n13309, ZN => n10341);
   U5132 : OAI222_X1 port map( A1 => n14940, A2 => n13342, B1 => n7812, B2 => 
                           n13339, C1 => n14681, C2 => n13336, ZN => n10444);
   U5133 : OAI222_X1 port map( A1 => n14934, A2 => n13342, B1 => n7808, B2 => 
                           n13339, C1 => n14675, C2 => n13336, ZN => n10443);
   U5134 : OAI222_X1 port map( A1 => n14928, A2 => n13342, B1 => n7804, B2 => 
                           n13339, C1 => n14669, C2 => n13336, ZN => n10442);
   U5135 : OAI222_X1 port map( A1 => n14922, A2 => n13342, B1 => n7800, B2 => 
                           n13339, C1 => n14663, C2 => n13336, ZN => n10441);
   U5136 : OAI222_X1 port map( A1 => n14916, A2 => n13342, B1 => n7796, B2 => 
                           n13339, C1 => n14657, C2 => n13336, ZN => n10440);
   U5137 : OAI222_X1 port map( A1 => n14910, A2 => n13342, B1 => n7792, B2 => 
                           n13339, C1 => n14651, C2 => n13336, ZN => n10439);
   U5138 : OAI222_X1 port map( A1 => n14904, A2 => n13342, B1 => n7788, B2 => 
                           n13339, C1 => n14645, C2 => n13336, ZN => n10438);
   U5139 : OAI222_X1 port map( A1 => n14898, A2 => n13342, B1 => n7784, B2 => 
                           n13339, C1 => n14639, C2 => n13336, ZN => n10437);
   U5140 : OAI222_X1 port map( A1 => n14933, A2 => n13351, B1 => n7809, B2 => 
                           n13348, C1 => n14675, C2 => n13345, ZN => n10475);
   U5141 : OAI222_X1 port map( A1 => n14927, A2 => n13351, B1 => n7805, B2 => 
                           n13348, C1 => n14669, C2 => n13345, ZN => n10474);
   U5142 : OAI222_X1 port map( A1 => n14921, A2 => n13351, B1 => n7801, B2 => 
                           n13348, C1 => n14663, C2 => n13345, ZN => n10473);
   U5143 : OAI222_X1 port map( A1 => n14915, A2 => n13351, B1 => n7797, B2 => 
                           n13348, C1 => n14657, C2 => n13345, ZN => n10472);
   U5144 : OAI222_X1 port map( A1 => n14909, A2 => n13351, B1 => n7793, B2 => 
                           n13348, C1 => n14651, C2 => n13345, ZN => n10471);
   U5145 : OAI222_X1 port map( A1 => n14903, A2 => n13351, B1 => n7789, B2 => 
                           n13348, C1 => n14645, C2 => n13345, ZN => n10470);
   U5146 : OAI222_X1 port map( A1 => n14897, A2 => n13351, B1 => n7785, B2 => 
                           n13348, C1 => n14639, C2 => n13345, ZN => n10469);
   U5147 : OAI222_X1 port map( A1 => n14939, A2 => n13378, B1 => n6737, B2 => 
                           n13375, C1 => n14681, C2 => n13372, ZN => n10572);
   U5148 : OAI222_X1 port map( A1 => n14933, A2 => n13378, B1 => n6761, B2 => 
                           n13375, C1 => n14675, C2 => n13372, ZN => n10571);
   U5149 : OAI222_X1 port map( A1 => n14927, A2 => n13378, B1 => n6785, B2 => 
                           n13375, C1 => n14669, C2 => n13372, ZN => n10570);
   U5150 : OAI222_X1 port map( A1 => n14921, A2 => n13378, B1 => n6809, B2 => 
                           n13375, C1 => n14663, C2 => n13372, ZN => n10569);
   U5151 : OAI222_X1 port map( A1 => n14915, A2 => n13378, B1 => n6833, B2 => 
                           n13375, C1 => n14657, C2 => n13372, ZN => n10568);
   U5152 : OAI222_X1 port map( A1 => n14909, A2 => n13378, B1 => n6857, B2 => 
                           n13375, C1 => n14651, C2 => n13372, ZN => n10567);
   U5153 : OAI222_X1 port map( A1 => n14903, A2 => n13378, B1 => n6881, B2 => 
                           n13375, C1 => n14645, C2 => n13372, ZN => n10566);
   U5154 : OAI222_X1 port map( A1 => n14897, A2 => n13378, B1 => n6905, B2 => 
                           n13375, C1 => n14639, C2 => n13372, ZN => n10565);
   U5155 : OAI222_X1 port map( A1 => n14938, A2 => n13459, B1 => n6734, B2 => 
                           n13456, C1 => n14680, C2 => n13453, ZN => n10860);
   U5156 : OAI222_X1 port map( A1 => n14932, A2 => n13459, B1 => n6758, B2 => 
                           n13456, C1 => n14674, C2 => n13453, ZN => n10859);
   U5157 : OAI222_X1 port map( A1 => n14926, A2 => n13459, B1 => n6782, B2 => 
                           n13456, C1 => n14668, C2 => n13453, ZN => n10858);
   U5158 : OAI222_X1 port map( A1 => n14920, A2 => n13459, B1 => n6806, B2 => 
                           n13456, C1 => n14662, C2 => n13453, ZN => n10857);
   U5159 : OAI222_X1 port map( A1 => n14914, A2 => n13459, B1 => n6830, B2 => 
                           n13456, C1 => n14656, C2 => n13453, ZN => n10856);
   U5160 : OAI222_X1 port map( A1 => n14908, A2 => n13459, B1 => n6854, B2 => 
                           n13456, C1 => n14650, C2 => n13453, ZN => n10855);
   U5161 : OAI222_X1 port map( A1 => n14902, A2 => n13459, B1 => n6878, B2 => 
                           n13456, C1 => n14644, C2 => n13453, ZN => n10854);
   U5162 : OAI222_X1 port map( A1 => n14896, A2 => n13459, B1 => n6902, B2 => 
                           n13456, C1 => n14638, C2 => n13453, ZN => n10853);
   U5163 : OAI222_X1 port map( A1 => n14932, A2 => n13477, B1 => n6756, B2 => 
                           n13474, C1 => n14674, C2 => n13471, ZN => n10923);
   U5164 : OAI222_X1 port map( A1 => n14920, A2 => n13477, B1 => n6804, B2 => 
                           n13474, C1 => n14662, C2 => n13471, ZN => n10921);
   U5165 : OAI222_X1 port map( A1 => n14914, A2 => n13477, B1 => n6828, B2 => 
                           n13474, C1 => n14656, C2 => n13471, ZN => n10920);
   U5166 : OAI222_X1 port map( A1 => n14908, A2 => n13477, B1 => n6852, B2 => 
                           n13474, C1 => n14650, C2 => n13471, ZN => n10919);
   U5167 : OAI222_X1 port map( A1 => n14902, A2 => n13477, B1 => n6876, B2 => 
                           n13474, C1 => n14644, C2 => n13471, ZN => n10918);
   U5168 : OAI222_X1 port map( A1 => n14896, A2 => n13477, B1 => n6900, B2 => 
                           n13474, C1 => n14638, C2 => n13471, ZN => n10917);
   U5169 : OAI222_X1 port map( A1 => n14938, A2 => n13540, B1 => n6731, B2 => 
                           n13537, C1 => n14679, C2 => n13534, ZN => n11148);
   U5170 : OAI222_X1 port map( A1 => n14932, A2 => n13540, B1 => n6755, B2 => 
                           n13537, C1 => n14673, C2 => n13534, ZN => n11147);
   U5171 : OAI222_X1 port map( A1 => n14926, A2 => n13540, B1 => n6779, B2 => 
                           n13537, C1 => n14667, C2 => n13534, ZN => n11146);
   U5172 : OAI222_X1 port map( A1 => n14920, A2 => n13540, B1 => n6803, B2 => 
                           n13537, C1 => n14661, C2 => n13534, ZN => n11145);
   U5173 : OAI222_X1 port map( A1 => n14914, A2 => n13540, B1 => n6827, B2 => 
                           n13537, C1 => n14655, C2 => n13534, ZN => n11144);
   U5174 : OAI222_X1 port map( A1 => n14908, A2 => n13540, B1 => n6851, B2 => 
                           n13537, C1 => n14649, C2 => n13534, ZN => n11143);
   U5175 : OAI222_X1 port map( A1 => n14902, A2 => n13540, B1 => n6875, B2 => 
                           n13537, C1 => n14643, C2 => n13534, ZN => n11142);
   U5176 : OAI222_X1 port map( A1 => n14896, A2 => n13540, B1 => n6899, B2 => 
                           n13537, C1 => n14637, C2 => n13534, ZN => n11141);
   U5177 : OAI222_X1 port map( A1 => n14937, A2 => n13621, B1 => n6728, B2 => 
                           n13618, C1 => n14679, C2 => n13615, ZN => n11436);
   U5178 : OAI222_X1 port map( A1 => n14931, A2 => n13621, B1 => n6752, B2 => 
                           n13618, C1 => n14673, C2 => n13615, ZN => n11435);
   U5179 : OAI222_X1 port map( A1 => n14925, A2 => n13621, B1 => n6776, B2 => 
                           n13618, C1 => n14667, C2 => n13615, ZN => n11434);
   U5180 : OAI222_X1 port map( A1 => n14919, A2 => n13621, B1 => n6800, B2 => 
                           n13618, C1 => n14661, C2 => n13615, ZN => n11433);
   U5181 : OAI222_X1 port map( A1 => n14913, A2 => n13621, B1 => n6824, B2 => 
                           n13618, C1 => n14655, C2 => n13615, ZN => n11432);
   U5182 : OAI222_X1 port map( A1 => n14907, A2 => n13621, B1 => n6848, B2 => 
                           n13618, C1 => n14649, C2 => n13615, ZN => n11431);
   U5183 : OAI222_X1 port map( A1 => n14901, A2 => n13621, B1 => n6872, B2 => 
                           n13618, C1 => n14643, C2 => n13615, ZN => n11430);
   U5184 : OAI222_X1 port map( A1 => n14895, A2 => n13621, B1 => n6896, B2 => 
                           n13618, C1 => n14637, C2 => n13615, ZN => n11429);
   U5185 : OAI222_X1 port map( A1 => n14937, A2 => n13630, B1 => n6727, B2 => 
                           n13627, C1 => n14679, C2 => n13624, ZN => n11468);
   U5186 : OAI222_X1 port map( A1 => n14887, A2 => n14498, B1 => n14494, B2 => 
                           n1649, C1 => n14629, C2 => n14493, ZN => n9924);
   U5187 : OAI222_X1 port map( A1 => n14887, A2 => n14507, B1 => n14503, B2 => 
                           n1628, C1 => n14629, C2 => n14502, ZN => n9956);
   U5188 : OAI222_X1 port map( A1 => n14891, A2 => n13359, B1 => n1510, B2 => 
                           n13356, C1 => n14633, C2 => n13354, ZN => n10500);
   U5189 : OAI222_X1 port map( A1 => n14891, A2 => n13368, B1 => n1486, B2 => 
                           n13365, C1 => n14633, C2 => n13363, ZN => n10532);
   U5190 : OAI222_X1 port map( A1 => n14891, A2 => n13404, B1 => n1447, B2 => 
                           n13401, C1 => n14633, C2 => n13399, ZN => n10660);
   U5191 : OAI222_X1 port map( A1 => n14891, A2 => n13440, B1 => n1351, B2 => 
                           n13437, C1 => n14632, C2 => n13435, ZN => n10788);
   U5192 : OAI222_X1 port map( A1 => n14891, A2 => n13449, B1 => n1327, B2 => 
                           n13446, C1 => n14632, C2 => n13444, ZN => n10820);
   U5193 : OAI222_X1 port map( A1 => n14890, A2 => n13521, B1 => n1192, B2 => 
                           n13518, C1 => n14632, C2 => n13516, ZN => n11076);
   U5194 : OAI222_X1 port map( A1 => n14890, A2 => n13530, B1 => n1168, B2 => 
                           n13527, C1 => n14632, C2 => n13525, ZN => n11108);
   U5195 : OAI222_X1 port map( A1 => n14888, A2 => n14343, B1 => n14339, B2 => 
                           n1036, C1 => n14630, C2 => n14338, ZN => n9380);
   U5196 : OAI222_X1 port map( A1 => n14888, A2 => n14334, B1 => n14330, B2 => 
                           n555, C1 => n14630, C2 => n14329, ZN => n9348);
   U5197 : OAI222_X1 port map( A1 => n14888, A2 => n14417, B1 => n14413, B2 => 
                           n459, C1 => n14629, C2 => n14412, ZN => n9636);
   U5198 : OAI222_X1 port map( A1 => n14888, A2 => n14426, B1 => n14422, B2 => 
                           n435, C1 => n14629, C2 => n14421, ZN => n9668);
   U5199 : OAI222_X1 port map( A1 => n14935, A2 => n14499, B1 => n14495, B2 => 
                           n388, C1 => n14677, C2 => n14493, ZN => n9932);
   U5200 : OAI222_X1 port map( A1 => n14929, A2 => n14499, B1 => n14494, B2 => 
                           n387, C1 => n14671, C2 => n14493, ZN => n9931);
   U5201 : OAI222_X1 port map( A1 => n14923, A2 => n14499, B1 => n14494, B2 => 
                           n386, C1 => n14665, C2 => n14493, ZN => n9930);
   U5202 : OAI222_X1 port map( A1 => n14917, A2 => n14499, B1 => n14494, B2 => 
                           n385, C1 => n14659, C2 => n14493, ZN => n9929);
   U5203 : OAI222_X1 port map( A1 => n14911, A2 => n14499, B1 => n14494, B2 => 
                           n384, C1 => n14653, C2 => n14493, ZN => n9928);
   U5204 : OAI222_X1 port map( A1 => n14905, A2 => n14499, B1 => n14494, B2 => 
                           n383, C1 => n14647, C2 => n14493, ZN => n9927);
   U5205 : OAI222_X1 port map( A1 => n14899, A2 => n14499, B1 => n14494, B2 => 
                           n382, C1 => n14641, C2 => n14493, ZN => n9926);
   U5206 : OAI222_X1 port map( A1 => n14893, A2 => n14499, B1 => n14494, B2 => 
                           n381, C1 => n14635, C2 => n14493, ZN => n9925);
   U5207 : OAI222_X1 port map( A1 => n14935, A2 => n14508, B1 => n14504, B2 => 
                           n380, C1 => n14677, C2 => n14502, ZN => n9964);
   U5208 : OAI222_X1 port map( A1 => n14929, A2 => n14508, B1 => n14503, B2 => 
                           n379, C1 => n14671, C2 => n14502, ZN => n9963);
   U5209 : OAI222_X1 port map( A1 => n14923, A2 => n14508, B1 => n14503, B2 => 
                           n378, C1 => n14665, C2 => n14502, ZN => n9962);
   U5210 : OAI222_X1 port map( A1 => n14917, A2 => n14508, B1 => n14503, B2 => 
                           n377, C1 => n14659, C2 => n14502, ZN => n9961);
   U5211 : OAI222_X1 port map( A1 => n14911, A2 => n14508, B1 => n14503, B2 => 
                           n376, C1 => n14653, C2 => n14502, ZN => n9960);
   U5212 : OAI222_X1 port map( A1 => n14905, A2 => n14508, B1 => n14503, B2 => 
                           n375, C1 => n14647, C2 => n14502, ZN => n9959);
   U5213 : OAI222_X1 port map( A1 => n14899, A2 => n14508, B1 => n14503, B2 => 
                           n374, C1 => n14641, C2 => n14502, ZN => n9958);
   U5214 : OAI222_X1 port map( A1 => n14893, A2 => n14508, B1 => n14503, B2 => 
                           n373, C1 => n14635, C2 => n14502, ZN => n9957);
   U5215 : OAI222_X1 port map( A1 => n14936, A2 => n14335, B1 => n14331, B2 => 
                           n348, C1 => n14678, C2 => n14329, ZN => n9356);
   U5216 : OAI222_X1 port map( A1 => n14930, A2 => n14335, B1 => n14330, B2 => 
                           n347, C1 => n14672, C2 => n14329, ZN => n9355);
   U5217 : OAI222_X1 port map( A1 => n14924, A2 => n14335, B1 => n14330, B2 => 
                           n346, C1 => n14666, C2 => n14329, ZN => n9354);
   U5218 : OAI222_X1 port map( A1 => n14918, A2 => n14335, B1 => n14330, B2 => 
                           n345, C1 => n14660, C2 => n14329, ZN => n9353);
   U5219 : OAI222_X1 port map( A1 => n14912, A2 => n14335, B1 => n14330, B2 => 
                           n344, C1 => n14654, C2 => n14329, ZN => n9352);
   U5220 : OAI222_X1 port map( A1 => n14906, A2 => n14335, B1 => n14330, B2 => 
                           n343, C1 => n14648, C2 => n14329, ZN => n9351);
   U5221 : OAI222_X1 port map( A1 => n14900, A2 => n14335, B1 => n14330, B2 => 
                           n342, C1 => n14642, C2 => n14329, ZN => n9350);
   U5222 : OAI222_X1 port map( A1 => n14894, A2 => n14335, B1 => n14330, B2 => 
                           n341, C1 => n14636, C2 => n14329, ZN => n9349);
   U5223 : OAI222_X1 port map( A1 => n14936, A2 => n14344, B1 => n14340, B2 => 
                           n340, C1 => n14678, C2 => n14338, ZN => n9388);
   U5224 : OAI222_X1 port map( A1 => n14930, A2 => n14344, B1 => n14339, B2 => 
                           n339, C1 => n14672, C2 => n14338, ZN => n9387);
   U5225 : OAI222_X1 port map( A1 => n14924, A2 => n14344, B1 => n14339, B2 => 
                           n338, C1 => n14666, C2 => n14338, ZN => n9386);
   U5226 : OAI222_X1 port map( A1 => n14918, A2 => n14344, B1 => n14339, B2 => 
                           n337, C1 => n14660, C2 => n14338, ZN => n9385);
   U5227 : OAI222_X1 port map( A1 => n14912, A2 => n14344, B1 => n14339, B2 => 
                           n336, C1 => n14654, C2 => n14338, ZN => n9384);
   U5228 : OAI222_X1 port map( A1 => n14906, A2 => n14344, B1 => n14339, B2 => 
                           n335, C1 => n14648, C2 => n14338, ZN => n9383);
   U5229 : OAI222_X1 port map( A1 => n14900, A2 => n14344, B1 => n14339, B2 => 
                           n334, C1 => n14642, C2 => n14338, ZN => n9382);
   U5230 : OAI222_X1 port map( A1 => n14894, A2 => n14344, B1 => n14339, B2 => 
                           n333, C1 => n14636, C2 => n14338, ZN => n9381);
   U5231 : OAI222_X1 port map( A1 => n14936, A2 => n14418, B1 => n14414, B2 => 
                           n284, C1 => n14677, C2 => n14412, ZN => n9644);
   U5232 : OAI222_X1 port map( A1 => n14930, A2 => n14418, B1 => n14413, B2 => 
                           n283, C1 => n14671, C2 => n14412, ZN => n9643);
   U5233 : OAI222_X1 port map( A1 => n14924, A2 => n14418, B1 => n14413, B2 => 
                           n282, C1 => n14665, C2 => n14412, ZN => n9642);
   U5234 : OAI222_X1 port map( A1 => n14918, A2 => n14418, B1 => n14413, B2 => 
                           n281, C1 => n14659, C2 => n14412, ZN => n9641);
   U5235 : OAI222_X1 port map( A1 => n14912, A2 => n14418, B1 => n14413, B2 => 
                           n280, C1 => n14653, C2 => n14412, ZN => n9640);
   U5236 : OAI222_X1 port map( A1 => n14906, A2 => n14418, B1 => n14413, B2 => 
                           n279, C1 => n14647, C2 => n14412, ZN => n9639);
   U5237 : OAI222_X1 port map( A1 => n14900, A2 => n14418, B1 => n14413, B2 => 
                           n278, C1 => n14641, C2 => n14412, ZN => n9638);
   U5238 : OAI222_X1 port map( A1 => n14894, A2 => n14418, B1 => n14413, B2 => 
                           n277, C1 => n14635, C2 => n14412, ZN => n9637);
   U5239 : OAI222_X1 port map( A1 => n14936, A2 => n14427, B1 => n14423, B2 => 
                           n276, C1 => n14677, C2 => n14421, ZN => n9676);
   U5240 : OAI222_X1 port map( A1 => n14930, A2 => n14427, B1 => n14422, B2 => 
                           n275, C1 => n14671, C2 => n14421, ZN => n9675);
   U5241 : OAI222_X1 port map( A1 => n14924, A2 => n14427, B1 => n14422, B2 => 
                           n274, C1 => n14665, C2 => n14421, ZN => n9674);
   U5242 : OAI222_X1 port map( A1 => n14918, A2 => n14427, B1 => n14422, B2 => 
                           n273, C1 => n14659, C2 => n14421, ZN => n9673);
   U5243 : OAI222_X1 port map( A1 => n14912, A2 => n14427, B1 => n14422, B2 => 
                           n272, C1 => n14653, C2 => n14421, ZN => n9672);
   U5244 : OAI222_X1 port map( A1 => n14906, A2 => n14427, B1 => n14422, B2 => 
                           n271, C1 => n14647, C2 => n14421, ZN => n9671);
   U5245 : OAI222_X1 port map( A1 => n14900, A2 => n14427, B1 => n14422, B2 => 
                           n270, C1 => n14641, C2 => n14421, ZN => n9670);
   U5246 : OAI222_X1 port map( A1 => n14894, A2 => n14427, B1 => n14422, B2 => 
                           n269, C1 => n14635, C2 => n14421, ZN => n9669);
   U5247 : OAI222_X1 port map( A1 => n14939, A2 => n13360, B1 => n211, B2 => 
                           n13357, C1 => n14681, C2 => n13354, ZN => n10508);
   U5248 : OAI222_X1 port map( A1 => n14933, A2 => n13360, B1 => n210, B2 => 
                           n13357, C1 => n14675, C2 => n13354, ZN => n10507);
   U5249 : OAI222_X1 port map( A1 => n14927, A2 => n13360, B1 => n209, B2 => 
                           n13357, C1 => n14669, C2 => n13354, ZN => n10506);
   U5250 : OAI222_X1 port map( A1 => n14921, A2 => n13360, B1 => n208, B2 => 
                           n13357, C1 => n14663, C2 => n13354, ZN => n10505);
   U5251 : OAI222_X1 port map( A1 => n14915, A2 => n13360, B1 => n207, B2 => 
                           n13357, C1 => n14657, C2 => n13354, ZN => n10504);
   U5252 : OAI222_X1 port map( A1 => n14909, A2 => n13360, B1 => n206, B2 => 
                           n13357, C1 => n14651, C2 => n13354, ZN => n10503);
   U5253 : OAI222_X1 port map( A1 => n14903, A2 => n13360, B1 => n205, B2 => 
                           n13357, C1 => n14645, C2 => n13354, ZN => n10502);
   U5254 : OAI222_X1 port map( A1 => n14897, A2 => n13360, B1 => n204, B2 => 
                           n13357, C1 => n14639, C2 => n13354, ZN => n10501);
   U5255 : OAI222_X1 port map( A1 => n14939, A2 => n13369, B1 => n203, B2 => 
                           n13366, C1 => n14681, C2 => n13363, ZN => n10540);
   U5256 : OAI222_X1 port map( A1 => n14933, A2 => n13369, B1 => n202, B2 => 
                           n13366, C1 => n14675, C2 => n13363, ZN => n10539);
   U5257 : OAI222_X1 port map( A1 => n14927, A2 => n13369, B1 => n201, B2 => 
                           n13366, C1 => n14669, C2 => n13363, ZN => n10538);
   U5258 : OAI222_X1 port map( A1 => n14921, A2 => n13369, B1 => n200, B2 => 
                           n13366, C1 => n14663, C2 => n13363, ZN => n10537);
   U5259 : OAI222_X1 port map( A1 => n14915, A2 => n13369, B1 => n199, B2 => 
                           n13366, C1 => n14657, C2 => n13363, ZN => n10536);
   U5260 : OAI222_X1 port map( A1 => n14909, A2 => n13369, B1 => n198, B2 => 
                           n13366, C1 => n14651, C2 => n13363, ZN => n10535);
   U5261 : OAI222_X1 port map( A1 => n14903, A2 => n13369, B1 => n197, B2 => 
                           n13366, C1 => n14645, C2 => n13363, ZN => n10534);
   U5262 : OAI222_X1 port map( A1 => n14897, A2 => n13369, B1 => n196, B2 => 
                           n13366, C1 => n14639, C2 => n13363, ZN => n10533);
   U5263 : OAI222_X1 port map( A1 => n14939, A2 => n13405, B1 => n187, B2 => 
                           n13402, C1 => n14681, C2 => n13399, ZN => n10668);
   U5264 : OAI222_X1 port map( A1 => n14933, A2 => n13405, B1 => n186, B2 => 
                           n13402, C1 => n14675, C2 => n13399, ZN => n10667);
   U5265 : OAI222_X1 port map( A1 => n14927, A2 => n13405, B1 => n185, B2 => 
                           n13402, C1 => n14669, C2 => n13399, ZN => n10666);
   U5266 : OAI222_X1 port map( A1 => n14921, A2 => n13405, B1 => n184, B2 => 
                           n13402, C1 => n14663, C2 => n13399, ZN => n10665);
   U5267 : OAI222_X1 port map( A1 => n14915, A2 => n13405, B1 => n183, B2 => 
                           n13402, C1 => n14657, C2 => n13399, ZN => n10664);
   U5268 : OAI222_X1 port map( A1 => n14909, A2 => n13405, B1 => n182, B2 => 
                           n13402, C1 => n14651, C2 => n13399, ZN => n10663);
   U5269 : OAI222_X1 port map( A1 => n14903, A2 => n13405, B1 => n181, B2 => 
                           n13402, C1 => n14645, C2 => n13399, ZN => n10662);
   U5270 : OAI222_X1 port map( A1 => n14897, A2 => n13405, B1 => n180, B2 => 
                           n13402, C1 => n14639, C2 => n13399, ZN => n10661);
   U5271 : OAI222_X1 port map( A1 => n14939, A2 => n13441, B1 => n155, B2 => 
                           n13438, C1 => n14680, C2 => n13435, ZN => n10796);
   U5272 : OAI222_X1 port map( A1 => n14933, A2 => n13441, B1 => n154, B2 => 
                           n13438, C1 => n14674, C2 => n13435, ZN => n10795);
   U5273 : OAI222_X1 port map( A1 => n14927, A2 => n13441, B1 => n153, B2 => 
                           n13438, C1 => n14668, C2 => n13435, ZN => n10794);
   U5274 : OAI222_X1 port map( A1 => n14921, A2 => n13441, B1 => n152, B2 => 
                           n13438, C1 => n14662, C2 => n13435, ZN => n10793);
   U5275 : OAI222_X1 port map( A1 => n14915, A2 => n13441, B1 => n151, B2 => 
                           n13438, C1 => n14656, C2 => n13435, ZN => n10792);
   U5276 : OAI222_X1 port map( A1 => n14909, A2 => n13441, B1 => n150, B2 => 
                           n13438, C1 => n14650, C2 => n13435, ZN => n10791);
   U5277 : OAI222_X1 port map( A1 => n14903, A2 => n13441, B1 => n149, B2 => 
                           n13438, C1 => n14644, C2 => n13435, ZN => n10790);
   U5278 : OAI222_X1 port map( A1 => n14897, A2 => n13441, B1 => n148, B2 => 
                           n13438, C1 => n14638, C2 => n13435, ZN => n10789);
   U5279 : OAI222_X1 port map( A1 => n14939, A2 => n13450, B1 => n147, B2 => 
                           n13447, C1 => n14680, C2 => n13444, ZN => n10828);
   U5280 : OAI222_X1 port map( A1 => n14933, A2 => n13450, B1 => n146, B2 => 
                           n13447, C1 => n14674, C2 => n13444, ZN => n10827);
   U5281 : OAI222_X1 port map( A1 => n14927, A2 => n13450, B1 => n145, B2 => 
                           n13447, C1 => n14668, C2 => n13444, ZN => n10826);
   U5282 : OAI222_X1 port map( A1 => n14921, A2 => n13450, B1 => n144, B2 => 
                           n13447, C1 => n14662, C2 => n13444, ZN => n10825);
   U5283 : OAI222_X1 port map( A1 => n14915, A2 => n13450, B1 => n143, B2 => 
                           n13447, C1 => n14656, C2 => n13444, ZN => n10824);
   U5284 : OAI222_X1 port map( A1 => n14909, A2 => n13450, B1 => n142, B2 => 
                           n13447, C1 => n14650, C2 => n13444, ZN => n10823);
   U5285 : OAI222_X1 port map( A1 => n14903, A2 => n13450, B1 => n141, B2 => 
                           n13447, C1 => n14644, C2 => n13444, ZN => n10822);
   U5286 : OAI222_X1 port map( A1 => n14897, A2 => n13450, B1 => n140, B2 => 
                           n13447, C1 => n14638, C2 => n13444, ZN => n10821);
   U5287 : OAI222_X1 port map( A1 => n14938, A2 => n13522, B1 => n98, B2 => 
                           n13519, C1 => n14680, C2 => n13516, ZN => n11084);
   U5288 : OAI222_X1 port map( A1 => n14932, A2 => n13522, B1 => n97, B2 => 
                           n13519, C1 => n14674, C2 => n13516, ZN => n11083);
   U5289 : OAI222_X1 port map( A1 => n14926, A2 => n13522, B1 => n92, B2 => 
                           n13519, C1 => n14668, C2 => n13516, ZN => n11082);
   U5290 : OAI222_X1 port map( A1 => n14920, A2 => n13522, B1 => n91, B2 => 
                           n13519, C1 => n14662, C2 => n13516, ZN => n11081);
   U5291 : OAI222_X1 port map( A1 => n14914, A2 => n13522, B1 => n86, B2 => 
                           n13519, C1 => n14656, C2 => n13516, ZN => n11080);
   U5292 : OAI222_X1 port map( A1 => n14908, A2 => n13522, B1 => n85, B2 => 
                           n13519, C1 => n14650, C2 => n13516, ZN => n11079);
   U5293 : OAI222_X1 port map( A1 => n14902, A2 => n13522, B1 => n80, B2 => 
                           n13519, C1 => n14644, C2 => n13516, ZN => n11078);
   U5294 : OAI222_X1 port map( A1 => n14896, A2 => n13522, B1 => n79, B2 => 
                           n13519, C1 => n14638, C2 => n13516, ZN => n11077);
   U5295 : OAI222_X1 port map( A1 => n14938, A2 => n13531, B1 => n74, B2 => 
                           n13528, C1 => n14680, C2 => n13525, ZN => n11116);
   U5296 : OAI222_X1 port map( A1 => n14932, A2 => n13531, B1 => n73, B2 => 
                           n13528, C1 => n14674, C2 => n13525, ZN => n11115);
   U5297 : OAI222_X1 port map( A1 => n14926, A2 => n13531, B1 => n70, B2 => 
                           n13528, C1 => n14668, C2 => n13525, ZN => n11114);
   U5298 : OAI222_X1 port map( A1 => n14920, A2 => n13531, B1 => n69, B2 => 
                           n13528, C1 => n14662, C2 => n13525, ZN => n11113);
   U5299 : OAI222_X1 port map( A1 => n14914, A2 => n13531, B1 => n68, B2 => 
                           n13528, C1 => n14656, C2 => n13525, ZN => n11112);
   U5300 : OAI222_X1 port map( A1 => n14908, A2 => n13531, B1 => n67, B2 => 
                           n13528, C1 => n14650, C2 => n13525, ZN => n11111);
   U5301 : OAI222_X1 port map( A1 => n14902, A2 => n13531, B1 => n66, B2 => 
                           n13528, C1 => n14644, C2 => n13525, ZN => n11110);
   U5302 : OAI222_X1 port map( A1 => n14896, A2 => n13531, B1 => n65, B2 => 
                           n13528, C1 => n14638, C2 => n13525, ZN => n11109);
   U5303 : OAI222_X1 port map( A1 => n14940, A2 => n13261, B1 => n8898, B2 => 
                           n13258, C1 => n14682, C2 => n13255, ZN => n10156);
   U5304 : OAI222_X1 port map( A1 => n14934, A2 => n13261, B1 => n7904, B2 => 
                           n13258, C1 => n14676, C2 => n13255, ZN => n10155);
   U5305 : OAI222_X1 port map( A1 => n14928, A2 => n13261, B1 => n7901, B2 => 
                           n13258, C1 => n14670, C2 => n13255, ZN => n10154);
   U5306 : OAI222_X1 port map( A1 => n14922, A2 => n13261, B1 => n7898, B2 => 
                           n13258, C1 => n14664, C2 => n13255, ZN => n10153);
   U5307 : OAI222_X1 port map( A1 => n14916, A2 => n13261, B1 => n7895, B2 => 
                           n13258, C1 => n14658, C2 => n13255, ZN => n10152);
   U5308 : OAI222_X1 port map( A1 => n14910, A2 => n13261, B1 => n7892, B2 => 
                           n13258, C1 => n14652, C2 => n13255, ZN => n10151);
   U5309 : OAI222_X1 port map( A1 => n14904, A2 => n13261, B1 => n7889, B2 => 
                           n13258, C1 => n14646, C2 => n13255, ZN => n10150);
   U5310 : OAI222_X1 port map( A1 => n14898, A2 => n13261, B1 => n7886, B2 => 
                           n13258, C1 => n14640, C2 => n13255, ZN => n10149);
   U5311 : OAI222_X1 port map( A1 => n14934, A2 => n13270, B1 => n7905, B2 => 
                           n13267, C1 => n14676, C2 => n13264, ZN => n10187);
   U5312 : OAI222_X1 port map( A1 => n14928, A2 => n13270, B1 => n7902, B2 => 
                           n13267, C1 => n14670, C2 => n13264, ZN => n10186);
   U5313 : OAI222_X1 port map( A1 => n14922, A2 => n13270, B1 => n7899, B2 => 
                           n13267, C1 => n14664, C2 => n13264, ZN => n10185);
   U5314 : OAI222_X1 port map( A1 => n14916, A2 => n13270, B1 => n7896, B2 => 
                           n13267, C1 => n14658, C2 => n13264, ZN => n10184);
   U5315 : OAI222_X1 port map( A1 => n14910, A2 => n13270, B1 => n7893, B2 => 
                           n13267, C1 => n14652, C2 => n13264, ZN => n10183);
   U5316 : OAI222_X1 port map( A1 => n14904, A2 => n13270, B1 => n7890, B2 => 
                           n13267, C1 => n14646, C2 => n13264, ZN => n10182);
   U5317 : OAI222_X1 port map( A1 => n14898, A2 => n13270, B1 => n7887, B2 => 
                           n13267, C1 => n14640, C2 => n13264, ZN => n10181);
   U5318 : OAI222_X1 port map( A1 => n14940, A2 => n13279, B1 => n251, B2 => 
                           n13276, C1 => n14682, C2 => n13273, ZN => n10220);
   U5319 : OAI222_X1 port map( A1 => n14934, A2 => n13279, B1 => n250, B2 => 
                           n13276, C1 => n14676, C2 => n13273, ZN => n10219);
   U5320 : OAI222_X1 port map( A1 => n14928, A2 => n13279, B1 => n249, B2 => 
                           n13276, C1 => n14670, C2 => n13273, ZN => n10218);
   U5321 : OAI222_X1 port map( A1 => n14922, A2 => n13279, B1 => n248, B2 => 
                           n13276, C1 => n14664, C2 => n13273, ZN => n10217);
   U5322 : OAI222_X1 port map( A1 => n14916, A2 => n13279, B1 => n247, B2 => 
                           n13276, C1 => n14658, C2 => n13273, ZN => n10216);
   U5323 : OAI222_X1 port map( A1 => n14910, A2 => n13279, B1 => n246, B2 => 
                           n13276, C1 => n14652, C2 => n13273, ZN => n10215);
   U5324 : OAI222_X1 port map( A1 => n14904, A2 => n13279, B1 => n245, B2 => 
                           n13276, C1 => n14646, C2 => n13273, ZN => n10214);
   U5325 : OAI222_X1 port map( A1 => n14898, A2 => n13279, B1 => n244, B2 => 
                           n13276, C1 => n14640, C2 => n13273, ZN => n10213);
   U5326 : OAI222_X1 port map( A1 => n14940, A2 => n13288, B1 => n243, B2 => 
                           n13285, C1 => n14682, C2 => n13282, ZN => n10252);
   U5327 : OAI222_X1 port map( A1 => n14934, A2 => n13288, B1 => n242, B2 => 
                           n13285, C1 => n14676, C2 => n13282, ZN => n10251);
   U5328 : OAI222_X1 port map( A1 => n14928, A2 => n13288, B1 => n241, B2 => 
                           n13285, C1 => n14670, C2 => n13282, ZN => n10250);
   U5329 : OAI222_X1 port map( A1 => n14922, A2 => n13288, B1 => n240, B2 => 
                           n13285, C1 => n14664, C2 => n13282, ZN => n10249);
   U5330 : OAI222_X1 port map( A1 => n14916, A2 => n13288, B1 => n239, B2 => 
                           n13285, C1 => n14658, C2 => n13282, ZN => n10248);
   U5331 : OAI222_X1 port map( A1 => n14910, A2 => n13288, B1 => n238, B2 => 
                           n13285, C1 => n14652, C2 => n13282, ZN => n10247);
   U5332 : OAI222_X1 port map( A1 => n14904, A2 => n13288, B1 => n237, B2 => 
                           n13285, C1 => n14646, C2 => n13282, ZN => n10246);
   U5333 : OAI222_X1 port map( A1 => n14898, A2 => n13288, B1 => n236, B2 => 
                           n13285, C1 => n14640, C2 => n13282, ZN => n10245);
   U5334 : OAI222_X1 port map( A1 => n14772, A2 => n13234, B1 => n7413, B2 => 
                           n13231, C1 => n14514, C2 => n13228, ZN => n10032);
   U5335 : OAI222_X1 port map( A1 => n14797, A2 => n13234, B1 => n7293, B2 => 
                           n13231, C1 => n14544, C2 => n13228, ZN => n10037);
   U5336 : OAI222_X1 port map( A1 => n14791, A2 => n13234, B1 => n7317, B2 => 
                           n13231, C1 => n14538, C2 => n13228, ZN => n10036);
   U5337 : OAI222_X1 port map( A1 => n14785, A2 => n13234, B1 => n7341, B2 => 
                           n13231, C1 => n14532, C2 => n13228, ZN => n10035);
   U5338 : OAI222_X1 port map( A1 => n14779, A2 => n13234, B1 => n7365, B2 => 
                           n13231, C1 => n14526, C2 => n13228, ZN => n10034);
   U5339 : OAI222_X1 port map( A1 => n14773, A2 => n13234, B1 => n7389, B2 => 
                           n13231, C1 => n14520, C2 => n13228, ZN => n10033);
   U5340 : OAI222_X1 port map( A1 => n2615, A2 => n14087, B1 => n4251, B2 => 
                           n14084, C1 => n14076, C2 => n2156, ZN => n9160);
   U5341 : NOR4_X1 port map( A1 => n4252, A2 => n4253, A3 => n4254, A4 => n4255
                           , ZN => n4251);
   U5342 : NAND4_X1 port map( A1 => n4280, A2 => n4281, A3 => n4282, A4 => 
                           n4283, ZN => n4252);
   U5343 : NAND4_X1 port map( A1 => n4272, A2 => n4273, A3 => n4274, A4 => 
                           n4275, ZN => n4253);
   U5344 : OAI222_X1 port map( A1 => n2620, A2 => n13867, B1 => n5387, B2 => 
                           n13864, C1 => n13856, C2 => n2183, ZN => n9132);
   U5345 : NOR4_X1 port map( A1 => n5388, A2 => n5389, A3 => n5390, A4 => n5391
                           , ZN => n5387);
   U5346 : NAND4_X1 port map( A1 => n5416, A2 => n5417, A3 => n5418, A4 => 
                           n5419, ZN => n5388);
   U5347 : NAND4_X1 port map( A1 => n5408, A2 => n5409, A3 => n5410, A4 => 
                           n5411, ZN => n5389);
   U5348 : OAI222_X1 port map( A1 => n2618, A2 => n13867, B1 => n5461, B2 => 
                           n13864, C1 => n13856, C2 => n2185, ZN => n9130);
   U5349 : NOR4_X1 port map( A1 => n5462, A2 => n5463, A3 => n5464, A4 => n5465
                           , ZN => n5461);
   U5350 : NAND4_X1 port map( A1 => n5490, A2 => n5491, A3 => n5492, A4 => 
                           n5493, ZN => n5462);
   U5351 : NAND4_X1 port map( A1 => n5482, A2 => n5483, A3 => n5484, A4 => 
                           n5485, ZN => n5463);
   U5352 : OAI222_X1 port map( A1 => n2617, A2 => n13867, B1 => n5498, B2 => 
                           n13864, C1 => n13856, C2 => n2186, ZN => n9129);
   U5353 : NOR4_X1 port map( A1 => n5499, A2 => n5500, A3 => n5501, A4 => n5502
                           , ZN => n5498);
   U5354 : NAND4_X1 port map( A1 => n5527, A2 => n5528, A3 => n5529, A4 => 
                           n5530, ZN => n5499);
   U5355 : NAND4_X1 port map( A1 => n5519, A2 => n5520, A3 => n5521, A4 => 
                           n5522, ZN => n5500);
   U5356 : OAI222_X1 port map( A1 => n2616, A2 => n13867, B1 => n5535, B2 => 
                           n13864, C1 => n13856, C2 => n2187, ZN => n9128);
   U5357 : NOR4_X1 port map( A1 => n5536, A2 => n5537, A3 => n5538, A4 => n5539
                           , ZN => n5535);
   U5358 : NAND4_X1 port map( A1 => n5564, A2 => n5565, A3 => n5566, A4 => 
                           n5567, ZN => n5536);
   U5359 : NAND4_X1 port map( A1 => n5556, A2 => n5557, A3 => n5558, A4 => 
                           n5559, ZN => n5537);
   U5360 : OAI222_X1 port map( A1 => n2615, A2 => n13867, B1 => n5572, B2 => 
                           n13864, C1 => n13856, C2 => n2188, ZN => n9127);
   U5361 : NOR4_X1 port map( A1 => n5573, A2 => n5574, A3 => n5575, A4 => n5576
                           , ZN => n5572);
   U5362 : NAND4_X1 port map( A1 => n5601, A2 => n5602, A3 => n5603, A4 => 
                           n5604, ZN => n5573);
   U5363 : NAND4_X1 port map( A1 => n5593, A2 => n5594, A3 => n5595, A4 => 
                           n5596, ZN => n5574);
   U5364 : OAI222_X1 port map( A1 => n2601, A2 => n14085, B1 => n4769, B2 => 
                           n14082, C1 => n14077, C2 => n2170, ZN => n9146);
   U5365 : NOR4_X1 port map( A1 => n4770, A2 => n4771, A3 => n4772, A4 => n4773
                           , ZN => n4769);
   U5366 : NAND4_X1 port map( A1 => n4798, A2 => n4799, A3 => n4800, A4 => 
                           n4801, ZN => n4770);
   U5367 : NAND4_X1 port map( A1 => n4790, A2 => n4791, A3 => n4792, A4 => 
                           n4793, ZN => n4771);
   U5368 : OAI222_X1 port map( A1 => n2601, A2 => n13865, B1 => n6090, B2 => 
                           n13862, C1 => n13857, C2 => n2202, ZN => n9113);
   U5369 : NOR4_X1 port map( A1 => n6091, A2 => n6092, A3 => n6093, A4 => n6094
                           , ZN => n6090);
   U5370 : NAND4_X1 port map( A1 => n6119, A2 => n6120, A3 => n6121, A4 => 
                           n6122, ZN => n6091);
   U5371 : NAND4_X1 port map( A1 => n6111, A2 => n6112, A3 => n6113, A4 => 
                           n6114, ZN => n6092);
   U5372 : OAI222_X1 port map( A1 => n2600, A2 => n13865, B1 => n6127, B2 => 
                           n13862, C1 => n13857, C2 => n2203, ZN => n9112);
   U5373 : NOR4_X1 port map( A1 => n6128, A2 => n6129, A3 => n6130, A4 => n6131
                           , ZN => n6127);
   U5374 : NAND4_X1 port map( A1 => n6156, A2 => n6157, A3 => n6158, A4 => 
                           n6159, ZN => n6128);
   U5375 : NAND4_X1 port map( A1 => n6148, A2 => n6149, A3 => n6150, A4 => 
                           n6151, ZN => n6129);
   U5376 : OAI222_X1 port map( A1 => n2599, A2 => n13865, B1 => n6164, B2 => 
                           n13862, C1 => n13857, C2 => n2204, ZN => n9111);
   U5377 : NOR4_X1 port map( A1 => n6165, A2 => n6166, A3 => n6167, A4 => n6168
                           , ZN => n6164);
   U5378 : NAND4_X1 port map( A1 => n6193, A2 => n6194, A3 => n6195, A4 => 
                           n6196, ZN => n6165);
   U5379 : NAND4_X1 port map( A1 => n6185, A2 => n6186, A3 => n6187, A4 => 
                           n6188, ZN => n6166);
   U5380 : OAI222_X1 port map( A1 => n2598, A2 => n13865, B1 => n6201, B2 => 
                           n13862, C1 => n13857, C2 => n2205, ZN => n9110);
   U5381 : NOR4_X1 port map( A1 => n6202, A2 => n6203, A3 => n6204, A4 => n6205
                           , ZN => n6201);
   U5382 : NAND4_X1 port map( A1 => n6230, A2 => n6231, A3 => n6232, A4 => 
                           n6233, ZN => n6202);
   U5383 : NAND4_X1 port map( A1 => n6222, A2 => n6223, A3 => n6224, A4 => 
                           n6225, ZN => n6203);
   U5384 : OAI222_X1 port map( A1 => n2597, A2 => n13865, B1 => n6238, B2 => 
                           n13862, C1 => n13858, C2 => n2206, ZN => n9109);
   U5385 : NOR4_X1 port map( A1 => n6239, A2 => n6240, A3 => n6241, A4 => n6242
                           , ZN => n6238);
   U5386 : NAND4_X1 port map( A1 => n6267, A2 => n6268, A3 => n6269, A4 => 
                           n6270, ZN => n6239);
   U5387 : NAND4_X1 port map( A1 => n6259, A2 => n6260, A3 => n6261, A4 => 
                           n6262, ZN => n6240);
   U5388 : OAI222_X1 port map( A1 => n2596, A2 => n13865, B1 => n6275, B2 => 
                           n13862, C1 => n13858, C2 => n2207, ZN => n9108);
   U5389 : NOR4_X1 port map( A1 => n6276, A2 => n6277, A3 => n6278, A4 => n6279
                           , ZN => n6275);
   U5390 : NAND4_X1 port map( A1 => n6304, A2 => n6305, A3 => n6306, A4 => 
                           n6307, ZN => n6276);
   U5391 : NAND4_X1 port map( A1 => n6296, A2 => n6297, A3 => n6298, A4 => 
                           n6299, ZN => n6277);
   U5392 : OAI222_X1 port map( A1 => n2595, A2 => n13865, B1 => n6312, B2 => 
                           n13862, C1 => n13858, C2 => n2208, ZN => n9107);
   U5393 : NOR4_X1 port map( A1 => n6313, A2 => n6314, A3 => n6315, A4 => n6316
                           , ZN => n6312);
   U5394 : NAND4_X1 port map( A1 => n6341, A2 => n6342, A3 => n6343, A4 => 
                           n6344, ZN => n6313);
   U5395 : NAND4_X1 port map( A1 => n6333, A2 => n6334, A3 => n6335, A4 => 
                           n6336, ZN => n6314);
   U5396 : OAI222_X1 port map( A1 => n2594, A2 => n13865, B1 => n6349, B2 => 
                           n13862, C1 => n13858, C2 => n2209, ZN => n9106);
   U5397 : NOR4_X1 port map( A1 => n6350, A2 => n6351, A3 => n6352, A4 => n6353
                           , ZN => n6349);
   U5398 : NAND4_X1 port map( A1 => n6378, A2 => n6379, A3 => n6380, A4 => 
                           n6381, ZN => n6350);
   U5399 : NAND4_X1 port map( A1 => n6370, A2 => n6371, A3 => n6372, A4 => 
                           n6373, ZN => n6351);
   U5400 : OAI222_X1 port map( A1 => n2593, A2 => n13865, B1 => n6386, B2 => 
                           n13862, C1 => n13858, C2 => n2210, ZN => n9105);
   U5401 : NOR4_X1 port map( A1 => n6387, A2 => n6388, A3 => n6389, A4 => n6390
                           , ZN => n6386);
   U5402 : NAND4_X1 port map( A1 => n6415, A2 => n6416, A3 => n6417, A4 => 
                           n6418, ZN => n6387);
   U5403 : NAND4_X1 port map( A1 => n6407, A2 => n6408, A3 => n6409, A4 => 
                           n6410, ZN => n6388);
   U5404 : OAI222_X1 port map( A1 => n2592, A2 => n13865, B1 => n6423, B2 => 
                           n13862, C1 => n13858, C2 => n2211, ZN => n9104);
   U5405 : NOR4_X1 port map( A1 => n6424, A2 => n6425, A3 => n6426, A4 => n6427
                           , ZN => n6423);
   U5406 : NAND4_X1 port map( A1 => n6452, A2 => n6453, A3 => n6454, A4 => 
                           n6455, ZN => n6424);
   U5407 : NAND4_X1 port map( A1 => n6444, A2 => n6445, A3 => n6446, A4 => 
                           n6447, ZN => n6425);
   U5408 : OAI222_X1 port map( A1 => n2591, A2 => n13865, B1 => n6460, B2 => 
                           n13862, C1 => n13858, C2 => n2212, ZN => n9103);
   U5409 : NOR4_X1 port map( A1 => n6461, A2 => n6462, A3 => n6463, A4 => n6464
                           , ZN => n6460);
   U5410 : NAND4_X1 port map( A1 => n6489, A2 => n6490, A3 => n6491, A4 => 
                           n6492, ZN => n6461);
   U5411 : NAND4_X1 port map( A1 => n6481, A2 => n6482, A3 => n6483, A4 => 
                           n6484, ZN => n6462);
   U5412 : OAI222_X1 port map( A1 => n2603, A2 => n14086, B1 => n4695, B2 => 
                           n14083, C1 => n14077, C2 => n2168, ZN => n9148);
   U5413 : NOR4_X1 port map( A1 => n4696, A2 => n4697, A3 => n4698, A4 => n4699
                           , ZN => n4695);
   U5414 : NAND4_X1 port map( A1 => n4724, A2 => n4725, A3 => n4726, A4 => 
                           n4727, ZN => n4696);
   U5415 : NAND4_X1 port map( A1 => n4716, A2 => n4717, A3 => n4718, A4 => 
                           n4719, ZN => n4697);
   U5416 : OAI222_X1 port map( A1 => n2602, A2 => n14086, B1 => n4732, B2 => 
                           n14083, C1 => n14077, C2 => n2169, ZN => n9147);
   U5417 : NOR4_X1 port map( A1 => n4733, A2 => n4734, A3 => n4735, A4 => n4736
                           , ZN => n4732);
   U5418 : NAND4_X1 port map( A1 => n4761, A2 => n4762, A3 => n4763, A4 => 
                           n4764, ZN => n4733);
   U5419 : NAND4_X1 port map( A1 => n4753, A2 => n4754, A3 => n4755, A4 => 
                           n4756, ZN => n4734);
   U5420 : OAI222_X1 port map( A1 => n2603, A2 => n13866, B1 => n6016, B2 => 
                           n13863, C1 => n13857, C2 => n2200, ZN => n9115);
   U5421 : NOR4_X1 port map( A1 => n6017, A2 => n6018, A3 => n6019, A4 => n6020
                           , ZN => n6016);
   U5422 : NAND4_X1 port map( A1 => n6045, A2 => n6046, A3 => n6047, A4 => 
                           n6048, ZN => n6017);
   U5423 : NAND4_X1 port map( A1 => n6037, A2 => n6038, A3 => n6039, A4 => 
                           n6040, ZN => n6018);
   U5424 : OAI222_X1 port map( A1 => n2602, A2 => n13866, B1 => n6053, B2 => 
                           n13863, C1 => n13857, C2 => n2201, ZN => n9114);
   U5425 : NOR4_X1 port map( A1 => n6054, A2 => n6055, A3 => n6056, A4 => n6057
                           , ZN => n6053);
   U5426 : NAND4_X1 port map( A1 => n6082, A2 => n6083, A3 => n6084, A4 => 
                           n6085, ZN => n6054);
   U5427 : NAND4_X1 port map( A1 => n6074, A2 => n6075, A3 => n6076, A4 => 
                           n6077, ZN => n6055);
   U5428 : OAI222_X1 port map( A1 => n2590, A2 => n13865, B1 => n6497, B2 => 
                           n13862, C1 => n13858, C2 => n2213, ZN => n9102);
   U5429 : NOR4_X1 port map( A1 => n6498, A2 => n6499, A3 => n6500, A4 => n6501
                           , ZN => n6497);
   U5430 : NAND4_X1 port map( A1 => n6541, A2 => n6542, A3 => n6543, A4 => 
                           n6544, ZN => n6498);
   U5431 : NAND4_X1 port map( A1 => n6531, A2 => n6532, A3 => n6533, A4 => 
                           n6534, ZN => n6499);
   U5432 : OAI222_X1 port map( A1 => n2621, A2 => n14087, B1 => n3955, B2 => 
                           n14084, C1 => n14076, C2 => n2150, ZN => n9166);
   U5433 : NOR4_X1 port map( A1 => n3958, A2 => n3959, A3 => n3960, A4 => n3961
                           , ZN => n3955);
   U5434 : NAND4_X1 port map( A1 => n4038, A2 => n4039, A3 => n4040, A4 => 
                           n4041, ZN => n3958);
   U5435 : NAND4_X1 port map( A1 => n4014, A2 => n4015, A3 => n4016, A4 => 
                           n4017, ZN => n3959);
   U5436 : OAI222_X1 port map( A1 => n2621, A2 => n13867, B1 => n5276, B2 => 
                           n13864, C1 => n13856, C2 => n2182, ZN => n9133);
   U5437 : NOR4_X1 port map( A1 => n5279, A2 => n5280, A3 => n5281, A4 => n5282
                           , ZN => n5276);
   U5438 : NAND4_X1 port map( A1 => n5361, A2 => n5362, A3 => n5363, A4 => 
                           n5364, ZN => n5279);
   U5439 : NAND4_X1 port map( A1 => n5335, A2 => n5336, A3 => n5337, A4 => 
                           n5338, ZN => n5280);
   U5440 : OAI222_X1 port map( A1 => n7398, A2 => n13637, B1 => n14767, B2 => 
                           n13634, C1 => n14510, C2 => n13631, ZN => n11472);
   U5441 : OAI222_X1 port map( A1 => n14767, A2 => n14706, B1 => n7414, B2 => 
                           n14718, C1 => n14707, C2 => n14514, ZN => n10000);
   U5442 : OAI222_X1 port map( A1 => n14887, A2 => n13232, B1 => n6933, B2 => 
                           n13229, C1 => n14634, C2 => n13226, ZN => n10052);
   U5443 : OAI222_X1 port map( A1 => n14881, A2 => n13232, B1 => n6957, B2 => 
                           n13229, C1 => n14628, C2 => n13226, ZN => n10051);
   U5444 : OAI222_X1 port map( A1 => n14875, A2 => n13233, B1 => n6981, B2 => 
                           n13230, C1 => n14622, C2 => n13226, ZN => n10050);
   U5445 : OAI222_X1 port map( A1 => n14869, A2 => n13233, B1 => n7005, B2 => 
                           n13230, C1 => n14616, C2 => n13227, ZN => n10049);
   U5446 : OAI222_X1 port map( A1 => n14863, A2 => n13233, B1 => n7029, B2 => 
                           n13230, C1 => n14610, C2 => n13227, ZN => n10048);
   U5447 : OAI222_X1 port map( A1 => n14833, A2 => n13233, B1 => n7149, B2 => 
                           n13230, C1 => n14580, C2 => n13227, ZN => n10043);
   U5448 : OAI222_X1 port map( A1 => n14827, A2 => n13233, B1 => n7173, B2 => 
                           n13230, C1 => n14574, C2 => n13227, ZN => n10042);
   U5449 : OAI222_X1 port map( A1 => n6942, A2 => n13638, B1 => n14881, B2 => 
                           n13635, C1 => n14624, C2 => n13632, ZN => n11491);
   U5450 : OAI222_X1 port map( A1 => n6966, A2 => n13638, B1 => n14875, B2 => 
                           n13635, C1 => n14618, C2 => n13632, ZN => n11490);
   U5451 : OAI222_X1 port map( A1 => n6990, A2 => n13638, B1 => n14869, B2 => 
                           n13635, C1 => n14612, C2 => n13632, ZN => n11489);
   U5452 : OAI222_X1 port map( A1 => n7014, A2 => n13638, B1 => n14863, B2 => 
                           n13635, C1 => n14606, C2 => n13632, ZN => n11488);
   U5453 : OAI222_X1 port map( A1 => n7038, A2 => n13638, B1 => n14857, B2 => 
                           n13635, C1 => n14600, C2 => n13632, ZN => n11487);
   U5454 : OAI222_X1 port map( A1 => n7062, A2 => n13638, B1 => n14851, B2 => 
                           n13635, C1 => n14594, C2 => n13632, ZN => n11486);
   U5455 : OAI222_X1 port map( A1 => n7086, A2 => n13638, B1 => n14845, B2 => 
                           n13635, C1 => n14588, C2 => n13632, ZN => n11485);
   U5456 : OAI222_X1 port map( A1 => n7110, A2 => n13638, B1 => n14839, B2 => 
                           n13635, C1 => n14582, C2 => n13632, ZN => n11484);
   U5457 : OAI222_X1 port map( A1 => n7134, A2 => n13638, B1 => n14833, B2 => 
                           n13635, C1 => n14576, C2 => n13632, ZN => n11483);
   U5458 : OAI222_X1 port map( A1 => n7158, A2 => n13638, B1 => n14827, B2 => 
                           n13635, C1 => n14570, C2 => n13632, ZN => n11482);
   U5459 : OAI222_X1 port map( A1 => n7182, A2 => n13638, B1 => n14821, B2 => 
                           n13635, C1 => n14564, C2 => n13632, ZN => n11481);
   U5460 : OAI222_X1 port map( A1 => n7254, A2 => n13637, B1 => n14803, B2 => 
                           n13634, C1 => n14546, C2 => n13631, ZN => n11478);
   U5461 : OAI222_X1 port map( A1 => n7278, A2 => n13637, B1 => n14797, B2 => 
                           n13634, C1 => n14540, C2 => n13631, ZN => n11477);
   U5462 : OAI222_X1 port map( A1 => n7302, A2 => n13637, B1 => n14791, B2 => 
                           n13634, C1 => n14534, C2 => n13631, ZN => n11476);
   U5463 : OAI222_X1 port map( A1 => n7326, A2 => n13637, B1 => n14785, B2 => 
                           n13634, C1 => n14528, C2 => n13631, ZN => n11475);
   U5464 : OAI222_X1 port map( A1 => n7350, A2 => n13637, B1 => n14779, B2 => 
                           n13634, C1 => n14522, C2 => n13631, ZN => n11474);
   U5465 : OAI222_X1 port map( A1 => n7374, A2 => n13637, B1 => n14773, B2 => 
                           n13634, C1 => n14516, C2 => n13631, ZN => n11473);
   U5466 : OAI222_X1 port map( A1 => n7470, A2 => n13637, B1 => n14749, B2 => 
                           n13634, C1 => n14695, C2 => n13631, ZN => n11469);
   U5467 : OAI222_X1 port map( A1 => n14809, A2 => n13234, B1 => n7245, B2 => 
                           n13231, C1 => n14556, C2 => n13227, ZN => n10039);
   U5468 : OAI222_X1 port map( A1 => n14803, A2 => n13234, B1 => n7269, B2 => 
                           n13231, C1 => n14550, C2 => n13227, ZN => n10038);
   U5469 : OAI222_X1 port map( A1 => n7422, A2 => n13637, B1 => n14761, B2 => 
                           n13634, C1 => n14712, C2 => n13631, ZN => n11471);
   U5470 : OAI222_X1 port map( A1 => n7446, A2 => n13637, B1 => n14755, B2 => 
                           n13634, C1 => n14700, C2 => n13631, ZN => n11470);
   U5471 : OAI222_X1 port map( A1 => n14749, A2 => n13232, B1 => n7485, B2 => 
                           n13229, C1 => n14692, C2 => n13226, ZN => n10029);
   U5472 : OAI222_X1 port map( A1 => n14935, A2 => n13233, B1 => n6741, B2 => 
                           n13230, C1 => n14682, C2 => n13226, ZN => n10060);
   U5473 : OAI222_X1 port map( A1 => n14929, A2 => n13232, B1 => n6765, B2 => 
                           n13229, C1 => n14676, C2 => n13226, ZN => n10059);
   U5474 : OAI222_X1 port map( A1 => n14923, A2 => n13232, B1 => n6789, B2 => 
                           n13229, C1 => n14670, C2 => n13226, ZN => n10058);
   U5475 : OAI222_X1 port map( A1 => n14917, A2 => n13232, B1 => n6813, B2 => 
                           n13229, C1 => n14664, C2 => n13226, ZN => n10057);
   U5476 : OAI222_X1 port map( A1 => n14911, A2 => n13232, B1 => n6837, B2 => 
                           n13229, C1 => n14658, C2 => n13226, ZN => n10056);
   U5477 : OAI222_X1 port map( A1 => n14905, A2 => n13232, B1 => n6861, B2 => 
                           n13229, C1 => n14652, C2 => n13226, ZN => n10055);
   U5478 : OAI222_X1 port map( A1 => n14899, A2 => n13232, B1 => n6885, B2 => 
                           n13229, C1 => n14646, C2 => n13226, ZN => n10054);
   U5479 : OAI222_X1 port map( A1 => n14893, A2 => n13232, B1 => n6909, B2 => 
                           n13229, C1 => n14640, C2 => n13227, ZN => n10053);
   U5480 : OAI222_X1 port map( A1 => n14767, A2 => n14443, B1 => n7417, B2 => 
                           n14442, C1 => n14509, C2 => n14437, ZN => n9712);
   U5481 : OAI222_X1 port map( A1 => n14767, A2 => n14479, B1 => n7702, B2 => 
                           n14478, C1 => n14509, C2 => n14473, ZN => n9840);
   U5482 : OAI222_X1 port map( A1 => n14767, A2 => n14488, B1 => n7703, B2 => 
                           n14487, C1 => n14509, C2 => n14482, ZN => n9872);
   U5483 : OAI222_X1 port map( A1 => n14767, A2 => n14434, B1 => n7418, B2 => 
                           n14433, C1 => n14509, C2 => n14428, ZN => n9680);
   U5484 : OAI222_X1 port map( A1 => n14827, A2 => n14444, B1 => n7177, B2 => 
                           n14441, C1 => n14569, C2 => n14438, ZN => n9722);
   U5485 : OAI222_X1 port map( A1 => n14809, A2 => n14443, B1 => n7249, B2 => 
                           n14441, C1 => n14551, C2 => n14437, ZN => n9719);
   U5486 : OAI222_X1 port map( A1 => n14803, A2 => n14443, B1 => n7273, B2 => 
                           n14441, C1 => n14545, C2 => n14437, ZN => n9718);
   U5487 : OAI222_X1 port map( A1 => n14797, A2 => n14443, B1 => n7297, B2 => 
                           n14441, C1 => n14539, C2 => n14437, ZN => n9717);
   U5488 : OAI222_X1 port map( A1 => n14791, A2 => n14443, B1 => n7321, B2 => 
                           n14442, C1 => n14533, C2 => n14437, ZN => n9716);
   U5489 : OAI222_X1 port map( A1 => n14785, A2 => n14443, B1 => n7345, B2 => 
                           n14442, C1 => n14527, C2 => n14437, ZN => n9715);
   U5490 : OAI222_X1 port map( A1 => n14779, A2 => n14443, B1 => n7369, B2 => 
                           n14442, C1 => n14521, C2 => n14437, ZN => n9714);
   U5491 : OAI222_X1 port map( A1 => n14773, A2 => n14443, B1 => n7393, B2 => 
                           n14442, C1 => n14515, C2 => n14437, ZN => n9713);
   U5492 : OAI222_X1 port map( A1 => n14749, A2 => n14443, B1 => n7489, B2 => 
                           n14442, C1 => n14697, C2 => n14437, ZN => n9709);
   U5493 : OAI222_X1 port map( A1 => n14881, A2 => n14453, B1 => n6960, B2 => 
                           n14450, C1 => n14623, C2 => n14447, ZN => n9763);
   U5494 : OAI222_X1 port map( A1 => n14875, A2 => n14453, B1 => n6984, B2 => 
                           n14450, C1 => n14617, C2 => n14447, ZN => n9762);
   U5495 : OAI222_X1 port map( A1 => n14869, A2 => n14453, B1 => n7008, B2 => 
                           n14450, C1 => n14611, C2 => n14447, ZN => n9761);
   U5496 : OAI222_X1 port map( A1 => n14833, A2 => n14453, B1 => n7152, B2 => 
                           n14450, C1 => n14575, C2 => n14447, ZN => n9755);
   U5497 : OAI222_X1 port map( A1 => n14827, A2 => n14453, B1 => n7176, B2 => 
                           n14450, C1 => n14569, C2 => n14447, ZN => n9754);
   U5498 : OAI222_X1 port map( A1 => n14809, A2 => n14452, B1 => n7248, B2 => 
                           n14450, C1 => n14551, C2 => n14446, ZN => n9751);
   U5499 : OAI222_X1 port map( A1 => n14803, A2 => n14452, B1 => n7272, B2 => 
                           n14450, C1 => n14545, C2 => n14446, ZN => n9750);
   U5500 : OAI222_X1 port map( A1 => n14797, A2 => n14452, B1 => n7296, B2 => 
                           n14450, C1 => n14539, C2 => n14446, ZN => n9749);
   U5501 : OAI222_X1 port map( A1 => n14791, A2 => n14452, B1 => n7320, B2 => 
                           n14451, C1 => n14533, C2 => n14446, ZN => n9748);
   U5502 : OAI222_X1 port map( A1 => n14785, A2 => n14452, B1 => n7344, B2 => 
                           n14451, C1 => n14527, C2 => n14446, ZN => n9747);
   U5503 : OAI222_X1 port map( A1 => n14779, A2 => n14452, B1 => n7368, B2 => 
                           n14451, C1 => n14521, C2 => n14446, ZN => n9746);
   U5504 : OAI222_X1 port map( A1 => n14773, A2 => n14452, B1 => n7392, B2 => 
                           n14451, C1 => n14515, C2 => n14446, ZN => n9745);
   U5505 : OAI222_X1 port map( A1 => n14749, A2 => n14452, B1 => n7488, B2 => 
                           n14449, C1 => n14697, C2 => n14446, ZN => n9741);
   U5506 : OAI222_X1 port map( A1 => n14881, A2 => n14480, B1 => n7778, B2 => 
                           n14476, C1 => n14623, C2 => n14474, ZN => n9859);
   U5507 : OAI222_X1 port map( A1 => n14875, A2 => n14480, B1 => n7774, B2 => 
                           n14476, C1 => n14617, C2 => n14474, ZN => n9858);
   U5508 : OAI222_X1 port map( A1 => n14869, A2 => n14480, B1 => n7770, B2 => 
                           n14476, C1 => n14611, C2 => n14474, ZN => n9857);
   U5509 : OAI222_X1 port map( A1 => n14863, A2 => n14480, B1 => n7766, B2 => 
                           n14477, C1 => n14605, C2 => n14474, ZN => n9856);
   U5510 : OAI222_X1 port map( A1 => n14857, A2 => n14480, B1 => n7762, B2 => 
                           n14477, C1 => n14599, C2 => n14474, ZN => n9855);
   U5511 : OAI222_X1 port map( A1 => n14851, A2 => n14480, B1 => n7758, B2 => 
                           n14477, C1 => n14593, C2 => n14474, ZN => n9854);
   U5512 : OAI222_X1 port map( A1 => n14845, A2 => n14480, B1 => n7754, B2 => 
                           n14477, C1 => n14587, C2 => n14474, ZN => n9853);
   U5513 : OAI222_X1 port map( A1 => n14839, A2 => n14480, B1 => n7750, B2 => 
                           n14477, C1 => n14581, C2 => n14474, ZN => n9852);
   U5514 : OAI222_X1 port map( A1 => n14833, A2 => n14480, B1 => n7746, B2 => 
                           n14477, C1 => n14575, C2 => n14474, ZN => n9851);
   U5515 : OAI222_X1 port map( A1 => n14827, A2 => n14480, B1 => n7742, B2 => 
                           n14477, C1 => n14569, C2 => n14474, ZN => n9850);
   U5516 : OAI222_X1 port map( A1 => n14815, A2 => n14479, B1 => n7734, B2 => 
                           n14477, C1 => n14557, C2 => n14474, ZN => n9848);
   U5517 : OAI222_X1 port map( A1 => n14809, A2 => n14479, B1 => n7730, B2 => 
                           n14477, C1 => n14551, C2 => n14473, ZN => n9847);
   U5518 : OAI222_X1 port map( A1 => n14803, A2 => n14479, B1 => n7726, B2 => 
                           n14477, C1 => n14545, C2 => n14473, ZN => n9846);
   U5519 : OAI222_X1 port map( A1 => n14797, A2 => n14479, B1 => n7722, B2 => 
                           n14477, C1 => n14539, C2 => n14473, ZN => n9845);
   U5520 : OAI222_X1 port map( A1 => n14791, A2 => n14479, B1 => n7718, B2 => 
                           n14477, C1 => n14533, C2 => n14473, ZN => n9844);
   U5521 : OAI222_X1 port map( A1 => n14785, A2 => n14479, B1 => n7714, B2 => 
                           n14478, C1 => n14527, C2 => n14473, ZN => n9843);
   U5522 : OAI222_X1 port map( A1 => n14779, A2 => n14479, B1 => n7710, B2 => 
                           n14478, C1 => n14521, C2 => n14473, ZN => n9842);
   U5523 : OAI222_X1 port map( A1 => n14773, A2 => n14479, B1 => n7706, B2 => 
                           n14478, C1 => n14515, C2 => n14473, ZN => n9841);
   U5524 : OAI222_X1 port map( A1 => n14749, A2 => n14479, B1 => n7690, B2 => 
                           n14476, C1 => n14697, C2 => n14473, ZN => n9837);
   U5525 : OAI222_X1 port map( A1 => n14881, A2 => n14489, B1 => n7779, B2 => 
                           n14485, C1 => n14623, C2 => n14483, ZN => n9891);
   U5526 : OAI222_X1 port map( A1 => n14875, A2 => n14489, B1 => n7775, B2 => 
                           n14485, C1 => n14617, C2 => n14483, ZN => n9890);
   U5527 : OAI222_X1 port map( A1 => n14869, A2 => n14489, B1 => n7771, B2 => 
                           n14485, C1 => n14611, C2 => n14483, ZN => n9889);
   U5528 : OAI222_X1 port map( A1 => n14863, A2 => n14489, B1 => n7767, B2 => 
                           n14486, C1 => n14605, C2 => n14483, ZN => n9888);
   U5529 : OAI222_X1 port map( A1 => n14857, A2 => n14489, B1 => n7763, B2 => 
                           n14486, C1 => n14599, C2 => n14483, ZN => n9887);
   U5530 : OAI222_X1 port map( A1 => n14851, A2 => n14489, B1 => n7759, B2 => 
                           n14486, C1 => n14593, C2 => n14483, ZN => n9886);
   U5531 : OAI222_X1 port map( A1 => n14845, A2 => n14489, B1 => n7755, B2 => 
                           n14486, C1 => n14587, C2 => n14483, ZN => n9885);
   U5532 : OAI222_X1 port map( A1 => n14839, A2 => n14489, B1 => n7751, B2 => 
                           n14486, C1 => n14581, C2 => n14483, ZN => n9884);
   U5533 : OAI222_X1 port map( A1 => n14833, A2 => n14489, B1 => n7747, B2 => 
                           n14486, C1 => n14575, C2 => n14483, ZN => n9883);
   U5534 : OAI222_X1 port map( A1 => n14827, A2 => n14489, B1 => n7743, B2 => 
                           n14486, C1 => n14569, C2 => n14483, ZN => n9882);
   U5535 : OAI222_X1 port map( A1 => n14815, A2 => n14488, B1 => n7735, B2 => 
                           n14486, C1 => n14557, C2 => n14483, ZN => n9880);
   U5536 : OAI222_X1 port map( A1 => n14809, A2 => n14488, B1 => n7731, B2 => 
                           n14486, C1 => n14551, C2 => n14482, ZN => n9879);
   U5537 : OAI222_X1 port map( A1 => n14803, A2 => n14488, B1 => n7727, B2 => 
                           n14486, C1 => n14545, C2 => n14482, ZN => n9878);
   U5538 : OAI222_X1 port map( A1 => n14797, A2 => n14488, B1 => n7723, B2 => 
                           n14486, C1 => n14539, C2 => n14482, ZN => n9877);
   U5539 : OAI222_X1 port map( A1 => n14791, A2 => n14488, B1 => n7719, B2 => 
                           n14486, C1 => n14533, C2 => n14482, ZN => n9876);
   U5540 : OAI222_X1 port map( A1 => n14785, A2 => n14488, B1 => n7715, B2 => 
                           n14487, C1 => n14527, C2 => n14482, ZN => n9875);
   U5541 : OAI222_X1 port map( A1 => n14779, A2 => n14488, B1 => n7711, B2 => 
                           n14487, C1 => n14521, C2 => n14482, ZN => n9874);
   U5542 : OAI222_X1 port map( A1 => n14773, A2 => n14488, B1 => n7707, B2 => 
                           n14487, C1 => n14515, C2 => n14482, ZN => n9873);
   U5543 : OAI222_X1 port map( A1 => n14749, A2 => n14488, B1 => n7691, B2 => 
                           n14485, C1 => n14697, C2 => n14482, ZN => n9869);
   U5544 : OAI222_X1 port map( A1 => n14749, A2 => n14689, B1 => n7487, B2 => 
                           n14686, C1 => n14697, C2 => n14685, ZN => n9965);
   U5545 : OAI222_X1 port map( A1 => n14881, A2 => n14435, B1 => n6962, B2 => 
                           n14431, C1 => n14623, C2 => n14429, ZN => n9699);
   U5546 : OAI222_X1 port map( A1 => n14875, A2 => n14435, B1 => n6986, B2 => 
                           n14431, C1 => n14617, C2 => n14429, ZN => n9698);
   U5547 : OAI222_X1 port map( A1 => n14869, A2 => n14435, B1 => n7010, B2 => 
                           n14432, C1 => n14611, C2 => n14429, ZN => n9697);
   U5548 : OAI222_X1 port map( A1 => n14863, A2 => n14435, B1 => n7034, B2 => 
                           n14432, C1 => n14605, C2 => n14429, ZN => n9696);
   U5549 : OAI222_X1 port map( A1 => n14857, A2 => n14435, B1 => n7058, B2 => 
                           n14432, C1 => n14599, C2 => n14429, ZN => n9695);
   U5550 : OAI222_X1 port map( A1 => n14851, A2 => n14435, B1 => n7082, B2 => 
                           n14432, C1 => n14593, C2 => n14429, ZN => n9694);
   U5551 : OAI222_X1 port map( A1 => n14845, A2 => n14435, B1 => n7106, B2 => 
                           n14432, C1 => n14587, C2 => n14429, ZN => n9693);
   U5552 : OAI222_X1 port map( A1 => n14839, A2 => n14435, B1 => n7130, B2 => 
                           n14432, C1 => n14581, C2 => n14429, ZN => n9692);
   U5553 : OAI222_X1 port map( A1 => n14833, A2 => n14435, B1 => n7154, B2 => 
                           n14432, C1 => n14575, C2 => n14429, ZN => n9691);
   U5554 : OAI222_X1 port map( A1 => n14827, A2 => n14435, B1 => n7178, B2 => 
                           n14432, C1 => n14569, C2 => n14429, ZN => n9690);
   U5555 : OAI222_X1 port map( A1 => n14809, A2 => n14434, B1 => n7250, B2 => 
                           n14432, C1 => n14551, C2 => n14428, ZN => n9687);
   U5556 : OAI222_X1 port map( A1 => n14803, A2 => n14434, B1 => n7274, B2 => 
                           n14432, C1 => n14545, C2 => n14428, ZN => n9686);
   U5557 : OAI222_X1 port map( A1 => n14797, A2 => n14434, B1 => n7298, B2 => 
                           n14432, C1 => n14539, C2 => n14428, ZN => n9685);
   U5558 : OAI222_X1 port map( A1 => n14791, A2 => n14434, B1 => n7322, B2 => 
                           n14432, C1 => n14533, C2 => n14428, ZN => n9684);
   U5559 : OAI222_X1 port map( A1 => n14785, A2 => n14434, B1 => n7346, B2 => 
                           n14433, C1 => n14527, C2 => n14428, ZN => n9683);
   U5560 : OAI222_X1 port map( A1 => n14779, A2 => n14434, B1 => n7370, B2 => 
                           n14433, C1 => n14521, C2 => n14428, ZN => n9682);
   U5561 : OAI222_X1 port map( A1 => n14773, A2 => n14434, B1 => n7394, B2 => 
                           n14433, C1 => n14515, C2 => n14428, ZN => n9681);
   U5562 : OAI222_X1 port map( A1 => n14761, A2 => n14443, B1 => n7441, B2 => 
                           n14442, C1 => n14710, C2 => n14437, ZN => n9711);
   U5563 : OAI222_X1 port map( A1 => n14755, A2 => n14443, B1 => n7465, B2 => 
                           n14442, C1 => n14698, C2 => n14437, ZN => n9710);
   U5564 : OAI222_X1 port map( A1 => n14762, A2 => n14452, B1 => n7440, B2 => 
                           n14451, C1 => n14710, C2 => n14446, ZN => n9743);
   U5565 : OAI222_X1 port map( A1 => n14756, A2 => n14452, B1 => n7464, B2 => 
                           n14451, C1 => n14698, C2 => n14446, ZN => n9742);
   U5566 : OAI222_X1 port map( A1 => n14761, A2 => n14479, B1 => n7698, B2 => 
                           n14478, C1 => n14710, C2 => n14473, ZN => n9839);
   U5567 : OAI222_X1 port map( A1 => n14755, A2 => n14479, B1 => n7694, B2 => 
                           n14478, C1 => n14698, C2 => n14473, ZN => n9838);
   U5568 : OAI222_X1 port map( A1 => n14761, A2 => n14488, B1 => n7699, B2 => 
                           n14487, C1 => n14710, C2 => n14482, ZN => n9871);
   U5569 : OAI222_X1 port map( A1 => n14755, A2 => n14488, B1 => n7695, B2 => 
                           n14487, C1 => n14698, C2 => n14482, ZN => n9870);
   U5570 : OAI222_X1 port map( A1 => n14761, A2 => n14689, B1 => n7439, B2 => 
                           n14688, C1 => n14710, C2 => n14685, ZN => n9967);
   U5571 : OAI222_X1 port map( A1 => n14755, A2 => n14689, B1 => n7463, B2 => 
                           n14688, C1 => n14698, C2 => n14685, ZN => n9966);
   U5572 : OAI222_X1 port map( A1 => n14762, A2 => n14434, B1 => n7442, B2 => 
                           n14433, C1 => n14710, C2 => n14428, ZN => n9679);
   U5573 : OAI222_X1 port map( A1 => n14756, A2 => n14434, B1 => n7466, B2 => 
                           n14433, C1 => n14698, C2 => n14428, ZN => n9678);
   U5574 : OAI222_X1 port map( A1 => n14886, A2 => n13296, B1 => n6956, B2 => 
                           n13293, C1 => n14628, C2 => n13290, ZN => n10275);
   U5575 : OAI222_X1 port map( A1 => n14880, A2 => n13296, B1 => n6980, B2 => 
                           n13293, C1 => n14622, C2 => n13290, ZN => n10274);
   U5576 : OAI222_X1 port map( A1 => n14874, A2 => n13296, B1 => n7004, B2 => 
                           n13293, C1 => n14616, C2 => n13290, ZN => n10273);
   U5577 : OAI222_X1 port map( A1 => n14868, A2 => n13296, B1 => n7028, B2 => 
                           n13293, C1 => n14610, C2 => n13290, ZN => n10272);
   U5578 : OAI222_X1 port map( A1 => n14862, A2 => n13296, B1 => n7052, B2 => 
                           n13293, C1 => n14604, C2 => n13290, ZN => n10271);
   U5579 : OAI222_X1 port map( A1 => n14856, A2 => n13296, B1 => n7076, B2 => 
                           n13293, C1 => n14598, C2 => n13290, ZN => n10270);
   U5580 : OAI222_X1 port map( A1 => n14850, A2 => n13296, B1 => n7100, B2 => 
                           n13293, C1 => n14592, C2 => n13290, ZN => n10269);
   U5581 : OAI222_X1 port map( A1 => n14844, A2 => n13296, B1 => n7124, B2 => 
                           n13293, C1 => n14586, C2 => n13290, ZN => n10268);
   U5582 : OAI222_X1 port map( A1 => n14838, A2 => n13296, B1 => n7148, B2 => 
                           n13293, C1 => n14580, C2 => n13290, ZN => n10267);
   U5583 : OAI222_X1 port map( A1 => n14832, A2 => n13296, B1 => n7172, B2 => 
                           n13293, C1 => n14574, C2 => n13290, ZN => n10266);
   U5584 : OAI222_X1 port map( A1 => n14826, A2 => n13296, B1 => n7196, B2 => 
                           n13293, C1 => n14568, C2 => n13290, ZN => n10265);
   U5585 : OAI222_X1 port map( A1 => n14814, A2 => n13295, B1 => n7244, B2 => 
                           n13292, C1 => n14556, C2 => n13289, ZN => n10263);
   U5586 : OAI222_X1 port map( A1 => n14808, A2 => n13295, B1 => n7268, B2 => 
                           n13292, C1 => n14550, C2 => n13289, ZN => n10262);
   U5587 : OAI222_X1 port map( A1 => n14802, A2 => n13295, B1 => n7292, B2 => 
                           n13292, C1 => n14544, C2 => n13289, ZN => n10261);
   U5588 : OAI222_X1 port map( A1 => n14796, A2 => n13295, B1 => n7316, B2 => 
                           n13292, C1 => n14538, C2 => n13289, ZN => n10260);
   U5589 : OAI222_X1 port map( A1 => n14790, A2 => n13295, B1 => n7340, B2 => 
                           n13292, C1 => n14532, C2 => n13289, ZN => n10259);
   U5590 : OAI222_X1 port map( A1 => n14784, A2 => n13295, B1 => n7364, B2 => 
                           n13292, C1 => n14526, C2 => n13289, ZN => n10258);
   U5591 : OAI222_X1 port map( A1 => n14778, A2 => n13295, B1 => n7388, B2 => 
                           n13292, C1 => n14520, C2 => n13289, ZN => n10257);
   U5592 : OAI222_X1 port map( A1 => n14772, A2 => n13295, B1 => n7412, B2 => 
                           n13292, C1 => n14514, C2 => n13289, ZN => n10256);
   U5593 : OAI222_X1 port map( A1 => n14766, A2 => n13295, B1 => n7436, B2 => 
                           n13292, C1 => n14715, C2 => n13289, ZN => n10255);
   U5594 : OAI222_X1 port map( A1 => n14760, A2 => n13295, B1 => n7460, B2 => 
                           n13292, C1 => n14703, C2 => n13289, ZN => n10254);
   U5595 : OAI222_X1 port map( A1 => n14754, A2 => n13295, B1 => n7484, B2 => 
                           n13292, C1 => n14692, C2 => n13289, ZN => n10253);
   U5596 : OAI222_X1 port map( A1 => n14886, A2 => n13314, B1 => n6954, B2 => 
                           n13311, C1 => n14628, C2 => n13308, ZN => n10339);
   U5597 : OAI222_X1 port map( A1 => n14880, A2 => n13314, B1 => n6978, B2 => 
                           n13311, C1 => n14622, C2 => n13308, ZN => n10338);
   U5598 : OAI222_X1 port map( A1 => n14874, A2 => n13314, B1 => n7002, B2 => 
                           n13311, C1 => n14616, C2 => n13308, ZN => n10337);
   U5599 : OAI222_X1 port map( A1 => n14838, A2 => n13314, B1 => n7146, B2 => 
                           n13311, C1 => n14580, C2 => n13308, ZN => n10331);
   U5600 : OAI222_X1 port map( A1 => n14886, A2 => n13341, B1 => n7776, B2 => 
                           n13338, C1 => n14627, C2 => n13335, ZN => n10435);
   U5601 : OAI222_X1 port map( A1 => n14880, A2 => n13341, B1 => n7772, B2 => 
                           n13338, C1 => n14621, C2 => n13335, ZN => n10434);
   U5602 : OAI222_X1 port map( A1 => n14874, A2 => n13341, B1 => n7768, B2 => 
                           n13338, C1 => n14615, C2 => n13335, ZN => n10433);
   U5603 : OAI222_X1 port map( A1 => n14868, A2 => n13341, B1 => n7764, B2 => 
                           n13338, C1 => n14609, C2 => n13335, ZN => n10432);
   U5604 : OAI222_X1 port map( A1 => n14862, A2 => n13341, B1 => n7760, B2 => 
                           n13338, C1 => n14603, C2 => n13335, ZN => n10431);
   U5605 : OAI222_X1 port map( A1 => n14856, A2 => n13341, B1 => n7756, B2 => 
                           n13338, C1 => n14597, C2 => n13335, ZN => n10430);
   U5606 : OAI222_X1 port map( A1 => n14850, A2 => n13341, B1 => n7752, B2 => 
                           n13338, C1 => n14591, C2 => n13335, ZN => n10429);
   U5607 : OAI222_X1 port map( A1 => n14844, A2 => n13341, B1 => n7748, B2 => 
                           n13338, C1 => n14585, C2 => n13335, ZN => n10428);
   U5608 : OAI222_X1 port map( A1 => n14838, A2 => n13341, B1 => n7744, B2 => 
                           n13338, C1 => n14579, C2 => n13335, ZN => n10427);
   U5609 : OAI222_X1 port map( A1 => n14832, A2 => n13341, B1 => n7740, B2 => 
                           n13338, C1 => n14573, C2 => n13335, ZN => n10426);
   U5610 : OAI222_X1 port map( A1 => n14826, A2 => n13341, B1 => n7736, B2 => 
                           n13338, C1 => n14567, C2 => n13335, ZN => n10425);
   U5611 : OAI222_X1 port map( A1 => n14820, A2 => n13340, B1 => n7732, B2 => 
                           n13337, C1 => n14561, C2 => n13335, ZN => n10424);
   U5612 : OAI222_X1 port map( A1 => n14814, A2 => n13340, B1 => n7728, B2 => 
                           n13337, C1 => n14555, C2 => n13334, ZN => n10423);
   U5613 : OAI222_X1 port map( A1 => n14808, A2 => n13340, B1 => n7724, B2 => 
                           n13337, C1 => n14549, C2 => n13334, ZN => n10422);
   U5614 : OAI222_X1 port map( A1 => n14802, A2 => n13340, B1 => n7720, B2 => 
                           n13337, C1 => n14543, C2 => n13334, ZN => n10421);
   U5615 : OAI222_X1 port map( A1 => n14796, A2 => n13340, B1 => n7716, B2 => 
                           n13337, C1 => n14537, C2 => n13334, ZN => n10420);
   U5616 : OAI222_X1 port map( A1 => n14790, A2 => n13340, B1 => n7712, B2 => 
                           n13337, C1 => n14531, C2 => n13334, ZN => n10419);
   U5617 : OAI222_X1 port map( A1 => n14784, A2 => n13340, B1 => n7708, B2 => 
                           n13337, C1 => n14525, C2 => n13334, ZN => n10418);
   U5618 : OAI222_X1 port map( A1 => n14778, A2 => n13340, B1 => n7704, B2 => 
                           n13337, C1 => n14519, C2 => n13334, ZN => n10417);
   U5619 : OAI222_X1 port map( A1 => n14771, A2 => n13340, B1 => n7700, B2 => 
                           n13337, C1 => n14513, C2 => n13334, ZN => n10416);
   U5620 : OAI222_X1 port map( A1 => n14766, A2 => n13340, B1 => n7696, B2 => 
                           n13337, C1 => n14714, C2 => n13334, ZN => n10415);
   U5621 : OAI222_X1 port map( A1 => n14760, A2 => n13340, B1 => n7692, B2 => 
                           n13337, C1 => n14702, C2 => n13334, ZN => n10414);
   U5622 : OAI222_X1 port map( A1 => n14754, A2 => n13340, B1 => n7688, B2 => 
                           n13337, C1 => n14693, C2 => n13334, ZN => n10413);
   U5623 : OAI222_X1 port map( A1 => n14885, A2 => n13350, B1 => n7777, B2 => 
                           n13347, C1 => n14627, C2 => n13344, ZN => n10467);
   U5624 : OAI222_X1 port map( A1 => n14879, A2 => n13350, B1 => n7773, B2 => 
                           n13347, C1 => n14621, C2 => n13344, ZN => n10466);
   U5625 : OAI222_X1 port map( A1 => n14873, A2 => n13350, B1 => n7769, B2 => 
                           n13347, C1 => n14615, C2 => n13344, ZN => n10465);
   U5626 : OAI222_X1 port map( A1 => n14867, A2 => n13350, B1 => n7765, B2 => 
                           n13347, C1 => n14609, C2 => n13344, ZN => n10464);
   U5627 : OAI222_X1 port map( A1 => n14861, A2 => n13350, B1 => n7761, B2 => 
                           n13347, C1 => n14603, C2 => n13344, ZN => n10463);
   U5628 : OAI222_X1 port map( A1 => n14855, A2 => n13350, B1 => n7757, B2 => 
                           n13347, C1 => n14597, C2 => n13344, ZN => n10462);
   U5629 : OAI222_X1 port map( A1 => n14849, A2 => n13350, B1 => n7753, B2 => 
                           n13347, C1 => n14591, C2 => n13344, ZN => n10461);
   U5630 : OAI222_X1 port map( A1 => n14843, A2 => n13350, B1 => n7749, B2 => 
                           n13347, C1 => n14585, C2 => n13344, ZN => n10460);
   U5631 : OAI222_X1 port map( A1 => n14837, A2 => n13350, B1 => n7745, B2 => 
                           n13347, C1 => n14579, C2 => n13344, ZN => n10459);
   U5632 : OAI222_X1 port map( A1 => n14831, A2 => n13350, B1 => n7741, B2 => 
                           n13347, C1 => n14573, C2 => n13344, ZN => n10458);
   U5633 : OAI222_X1 port map( A1 => n14825, A2 => n13350, B1 => n7737, B2 => 
                           n13347, C1 => n14567, C2 => n13344, ZN => n10457);
   U5634 : OAI222_X1 port map( A1 => n14819, A2 => n13349, B1 => n2314, B2 => 
                           n13346, C1 => n14561, C2 => n13344, ZN => n10456);
   U5635 : OAI222_X1 port map( A1 => n14813, A2 => n13349, B1 => n7729, B2 => 
                           n13346, C1 => n14555, C2 => n13343, ZN => n10455);
   U5636 : OAI222_X1 port map( A1 => n14807, A2 => n13349, B1 => n7725, B2 => 
                           n13346, C1 => n14549, C2 => n13343, ZN => n10454);
   U5637 : OAI222_X1 port map( A1 => n14801, A2 => n13349, B1 => n7721, B2 => 
                           n13346, C1 => n14543, C2 => n13343, ZN => n10453);
   U5638 : OAI222_X1 port map( A1 => n14795, A2 => n13349, B1 => n7717, B2 => 
                           n13346, C1 => n14537, C2 => n13343, ZN => n10452);
   U5639 : OAI222_X1 port map( A1 => n14789, A2 => n13349, B1 => n7713, B2 => 
                           n13346, C1 => n14531, C2 => n13343, ZN => n10451);
   U5640 : OAI222_X1 port map( A1 => n14783, A2 => n13349, B1 => n7709, B2 => 
                           n13346, C1 => n14525, C2 => n13343, ZN => n10450);
   U5641 : OAI222_X1 port map( A1 => n14777, A2 => n13349, B1 => n7705, B2 => 
                           n13346, C1 => n14519, C2 => n13343, ZN => n10449);
   U5642 : OAI222_X1 port map( A1 => n14771, A2 => n13349, B1 => n7701, B2 => 
                           n13346, C1 => n14513, C2 => n13343, ZN => n10448);
   U5643 : OAI222_X1 port map( A1 => n14766, A2 => n13349, B1 => n7697, B2 => 
                           n13346, C1 => n14714, C2 => n13343, ZN => n10447);
   U5644 : OAI222_X1 port map( A1 => n14760, A2 => n13349, B1 => n7693, B2 => 
                           n13346, C1 => n14702, C2 => n13343, ZN => n10446);
   U5645 : OAI222_X1 port map( A1 => n14885, A2 => n13377, B1 => n6953, B2 => 
                           n13374, C1 => n14627, C2 => n13371, ZN => n10563);
   U5646 : OAI222_X1 port map( A1 => n14879, A2 => n13377, B1 => n6977, B2 => 
                           n13374, C1 => n14621, C2 => n13371, ZN => n10562);
   U5647 : OAI222_X1 port map( A1 => n14873, A2 => n13377, B1 => n7001, B2 => 
                           n13374, C1 => n14615, C2 => n13371, ZN => n10561);
   U5648 : OAI222_X1 port map( A1 => n14867, A2 => n13377, B1 => n7025, B2 => 
                           n13374, C1 => n14609, C2 => n13371, ZN => n10560);
   U5649 : OAI222_X1 port map( A1 => n14861, A2 => n13377, B1 => n7049, B2 => 
                           n13374, C1 => n14603, C2 => n13371, ZN => n10559);
   U5650 : OAI222_X1 port map( A1 => n14855, A2 => n13377, B1 => n7073, B2 => 
                           n13374, C1 => n14597, C2 => n13371, ZN => n10558);
   U5651 : OAI222_X1 port map( A1 => n14849, A2 => n13377, B1 => n7097, B2 => 
                           n13374, C1 => n14591, C2 => n13371, ZN => n10557);
   U5652 : OAI222_X1 port map( A1 => n14843, A2 => n13377, B1 => n7121, B2 => 
                           n13374, C1 => n14585, C2 => n13371, ZN => n10556);
   U5653 : OAI222_X1 port map( A1 => n14837, A2 => n13377, B1 => n7145, B2 => 
                           n13374, C1 => n14579, C2 => n13371, ZN => n10555);
   U5654 : OAI222_X1 port map( A1 => n14831, A2 => n13377, B1 => n7169, B2 => 
                           n13374, C1 => n14573, C2 => n13371, ZN => n10554);
   U5655 : OAI222_X1 port map( A1 => n14825, A2 => n13377, B1 => n7193, B2 => 
                           n13374, C1 => n14567, C2 => n13371, ZN => n10553);
   U5656 : OAI222_X1 port map( A1 => n14813, A2 => n13376, B1 => n7241, B2 => 
                           n13373, C1 => n14555, C2 => n13370, ZN => n10551);
   U5657 : OAI222_X1 port map( A1 => n14807, A2 => n13376, B1 => n7265, B2 => 
                           n13373, C1 => n14549, C2 => n13370, ZN => n10550);
   U5658 : OAI222_X1 port map( A1 => n14801, A2 => n13376, B1 => n7289, B2 => 
                           n13373, C1 => n14543, C2 => n13370, ZN => n10549);
   U5659 : OAI222_X1 port map( A1 => n14795, A2 => n13376, B1 => n7313, B2 => 
                           n13373, C1 => n14537, C2 => n13370, ZN => n10548);
   U5660 : OAI222_X1 port map( A1 => n14789, A2 => n13376, B1 => n7337, B2 => 
                           n13373, C1 => n14531, C2 => n13370, ZN => n10547);
   U5661 : OAI222_X1 port map( A1 => n14783, A2 => n13376, B1 => n7361, B2 => 
                           n13373, C1 => n14525, C2 => n13370, ZN => n10546);
   U5662 : OAI222_X1 port map( A1 => n14777, A2 => n13376, B1 => n7385, B2 => 
                           n13373, C1 => n14519, C2 => n13370, ZN => n10545);
   U5663 : OAI222_X1 port map( A1 => n14771, A2 => n13376, B1 => n7409, B2 => 
                           n13373, C1 => n14513, C2 => n13370, ZN => n10544);
   U5664 : OAI222_X1 port map( A1 => n14765, A2 => n13376, B1 => n7433, B2 => 
                           n13373, C1 => n14714, C2 => n13370, ZN => n10543);
   U5665 : OAI222_X1 port map( A1 => n14759, A2 => n13376, B1 => n7457, B2 => 
                           n13373, C1 => n14702, C2 => n13370, ZN => n10542);
   U5666 : OAI222_X1 port map( A1 => n14753, A2 => n13376, B1 => n7481, B2 => 
                           n13373, C1 => n14693, C2 => n13370, ZN => n10541);
   U5667 : OAI222_X1 port map( A1 => n14884, A2 => n13458, B1 => n6950, B2 => 
                           n13455, C1 => n14626, C2 => n13452, ZN => n10851);
   U5668 : OAI222_X1 port map( A1 => n14878, A2 => n13458, B1 => n6974, B2 => 
                           n13455, C1 => n14620, C2 => n13452, ZN => n10850);
   U5669 : OAI222_X1 port map( A1 => n14872, A2 => n13458, B1 => n6998, B2 => 
                           n13455, C1 => n14614, C2 => n13452, ZN => n10849);
   U5670 : OAI222_X1 port map( A1 => n14866, A2 => n13458, B1 => n7022, B2 => 
                           n13455, C1 => n14608, C2 => n13452, ZN => n10848);
   U5671 : OAI222_X1 port map( A1 => n14860, A2 => n13458, B1 => n7046, B2 => 
                           n13455, C1 => n14602, C2 => n13452, ZN => n10847);
   U5672 : OAI222_X1 port map( A1 => n14854, A2 => n13458, B1 => n7070, B2 => 
                           n13455, C1 => n14596, C2 => n13452, ZN => n10846);
   U5673 : OAI222_X1 port map( A1 => n14848, A2 => n13458, B1 => n7094, B2 => 
                           n13455, C1 => n14590, C2 => n13452, ZN => n10845);
   U5674 : OAI222_X1 port map( A1 => n14842, A2 => n13458, B1 => n7118, B2 => 
                           n13455, C1 => n14584, C2 => n13452, ZN => n10844);
   U5675 : OAI222_X1 port map( A1 => n14836, A2 => n13458, B1 => n7142, B2 => 
                           n13455, C1 => n14578, C2 => n13452, ZN => n10843);
   U5676 : OAI222_X1 port map( A1 => n14830, A2 => n13458, B1 => n7166, B2 => 
                           n13455, C1 => n14572, C2 => n13452, ZN => n10842);
   U5677 : OAI222_X1 port map( A1 => n14824, A2 => n13458, B1 => n7190, B2 => 
                           n13455, C1 => n14566, C2 => n13452, ZN => n10841);
   U5678 : OAI222_X1 port map( A1 => n14812, A2 => n13457, B1 => n7238, B2 => 
                           n13454, C1 => n14554, C2 => n13451, ZN => n10839);
   U5679 : OAI222_X1 port map( A1 => n14806, A2 => n13457, B1 => n7262, B2 => 
                           n13454, C1 => n14548, C2 => n13451, ZN => n10838);
   U5680 : OAI222_X1 port map( A1 => n14800, A2 => n13457, B1 => n7286, B2 => 
                           n13454, C1 => n14542, C2 => n13451, ZN => n10837);
   U5681 : OAI222_X1 port map( A1 => n14794, A2 => n13457, B1 => n7310, B2 => 
                           n13454, C1 => n14536, C2 => n13451, ZN => n10836);
   U5682 : OAI222_X1 port map( A1 => n14788, A2 => n13457, B1 => n7334, B2 => 
                           n13454, C1 => n14530, C2 => n13451, ZN => n10835);
   U5683 : OAI222_X1 port map( A1 => n14782, A2 => n13457, B1 => n7358, B2 => 
                           n13454, C1 => n14524, C2 => n13451, ZN => n10834);
   U5684 : OAI222_X1 port map( A1 => n14776, A2 => n13457, B1 => n7382, B2 => 
                           n13454, C1 => n14518, C2 => n13451, ZN => n10833);
   U5685 : OAI222_X1 port map( A1 => n14770, A2 => n13457, B1 => n7406, B2 => 
                           n13454, C1 => n14512, C2 => n13451, ZN => n10832);
   U5686 : OAI222_X1 port map( A1 => n14765, A2 => n13457, B1 => n7430, B2 => 
                           n13454, C1 => n14713, C2 => n13451, ZN => n10831);
   U5687 : OAI222_X1 port map( A1 => n14759, A2 => n13457, B1 => n7454, B2 => 
                           n13454, C1 => n14701, C2 => n13451, ZN => n10830);
   U5688 : OAI222_X1 port map( A1 => n14752, A2 => n13457, B1 => n7478, B2 => 
                           n13454, C1 => n14694, C2 => n13451, ZN => n10829);
   U5689 : OAI222_X1 port map( A1 => n14884, A2 => n13476, B1 => n6948, B2 => 
                           n13473, C1 => n14626, C2 => n13470, ZN => n10915);
   U5690 : OAI222_X1 port map( A1 => n14878, A2 => n13476, B1 => n6972, B2 => 
                           n13473, C1 => n14620, C2 => n13470, ZN => n10914);
   U5691 : OAI222_X1 port map( A1 => n14872, A2 => n13476, B1 => n6996, B2 => 
                           n13473, C1 => n14614, C2 => n13470, ZN => n10913);
   U5692 : OAI222_X1 port map( A1 => n14866, A2 => n13476, B1 => n7020, B2 => 
                           n13473, C1 => n14608, C2 => n13470, ZN => n10912);
   U5693 : OAI222_X1 port map( A1 => n14884, A2 => n13539, B1 => n6947, B2 => 
                           n13536, C1 => n14625, C2 => n13533, ZN => n11139);
   U5694 : OAI222_X1 port map( A1 => n14878, A2 => n13539, B1 => n6971, B2 => 
                           n13536, C1 => n14619, C2 => n13533, ZN => n11138);
   U5695 : OAI222_X1 port map( A1 => n14872, A2 => n13539, B1 => n6995, B2 => 
                           n13536, C1 => n14613, C2 => n13533, ZN => n11137);
   U5696 : OAI222_X1 port map( A1 => n14866, A2 => n13539, B1 => n7019, B2 => 
                           n13536, C1 => n14607, C2 => n13533, ZN => n11136);
   U5697 : OAI222_X1 port map( A1 => n14860, A2 => n13539, B1 => n7043, B2 => 
                           n13536, C1 => n14601, C2 => n13533, ZN => n11135);
   U5698 : OAI222_X1 port map( A1 => n14854, A2 => n13539, B1 => n7067, B2 => 
                           n13536, C1 => n14595, C2 => n13533, ZN => n11134);
   U5699 : OAI222_X1 port map( A1 => n14848, A2 => n13539, B1 => n7091, B2 => 
                           n13536, C1 => n14589, C2 => n13533, ZN => n11133);
   U5700 : OAI222_X1 port map( A1 => n14842, A2 => n13539, B1 => n7115, B2 => 
                           n13536, C1 => n14583, C2 => n13533, ZN => n11132);
   U5701 : OAI222_X1 port map( A1 => n14836, A2 => n13539, B1 => n7139, B2 => 
                           n13536, C1 => n14577, C2 => n13533, ZN => n11131);
   U5702 : OAI222_X1 port map( A1 => n14830, A2 => n13539, B1 => n7163, B2 => 
                           n13536, C1 => n14571, C2 => n13533, ZN => n11130);
   U5703 : OAI222_X1 port map( A1 => n14824, A2 => n13539, B1 => n7187, B2 => 
                           n13536, C1 => n14565, C2 => n13533, ZN => n11129);
   U5704 : OAI222_X1 port map( A1 => n14806, A2 => n13538, B1 => n7259, B2 => 
                           n13535, C1 => n14547, C2 => n13532, ZN => n11126);
   U5705 : OAI222_X1 port map( A1 => n14800, A2 => n13538, B1 => n7283, B2 => 
                           n13535, C1 => n14541, C2 => n13532, ZN => n11125);
   U5706 : OAI222_X1 port map( A1 => n14794, A2 => n13538, B1 => n7307, B2 => 
                           n13535, C1 => n14535, C2 => n13532, ZN => n11124);
   U5707 : OAI222_X1 port map( A1 => n14788, A2 => n13538, B1 => n7331, B2 => 
                           n13535, C1 => n14529, C2 => n13532, ZN => n11123);
   U5708 : OAI222_X1 port map( A1 => n14782, A2 => n13538, B1 => n7355, B2 => 
                           n13535, C1 => n14523, C2 => n13532, ZN => n11122);
   U5709 : OAI222_X1 port map( A1 => n14776, A2 => n13538, B1 => n7379, B2 => 
                           n13535, C1 => n14517, C2 => n13532, ZN => n11121);
   U5710 : OAI222_X1 port map( A1 => n14770, A2 => n13538, B1 => n7403, B2 => 
                           n13535, C1 => n14511, C2 => n13532, ZN => n11120);
   U5711 : OAI222_X1 port map( A1 => n14764, A2 => n13538, B1 => n7427, B2 => 
                           n13535, C1 => n14713, C2 => n13532, ZN => n11119);
   U5712 : OAI222_X1 port map( A1 => n14758, A2 => n13538, B1 => n7451, B2 => 
                           n13535, C1 => n14701, C2 => n13532, ZN => n11118);
   U5713 : OAI222_X1 port map( A1 => n14752, A2 => n13538, B1 => n7475, B2 => 
                           n13535, C1 => n14694, C2 => n13532, ZN => n11117);
   U5714 : OAI222_X1 port map( A1 => n14767, A2 => n14452, B1 => n7416, B2 => 
                           n14451, C1 => n14509, C2 => n14446, ZN => n9744);
   U5715 : OAI222_X1 port map( A1 => n14890, A2 => n14690, B1 => n6935, B2 => 
                           n14686, C1 => n14683, C2 => n14634, ZN => n9988);
   U5716 : OAI222_X1 port map( A1 => n14884, A2 => n14690, B1 => n6959, B2 => 
                           n14686, C1 => n14683, C2 => n14628, ZN => n9987);
   U5717 : OAI222_X1 port map( A1 => n14878, A2 => n14690, B1 => n6983, B2 => 
                           n14686, C1 => n14683, C2 => n14622, ZN => n9986);
   U5718 : OAI222_X1 port map( A1 => n14872, A2 => n14690, B1 => n7007, B2 => 
                           n14687, C1 => n14683, C2 => n14616, ZN => n9985);
   U5719 : OAI222_X1 port map( A1 => n14866, A2 => n14690, B1 => n7031, B2 => 
                           n14687, C1 => n14683, C2 => n14610, ZN => n9984);
   U5720 : OAI222_X1 port map( A1 => n14860, A2 => n14690, B1 => n7055, B2 => 
                           n14687, C1 => n14684, C2 => n14604, ZN => n9983);
   U5721 : OAI222_X1 port map( A1 => n14854, A2 => n14690, B1 => n7079, B2 => 
                           n14687, C1 => n14684, C2 => n14598, ZN => n9982);
   U5722 : OAI222_X1 port map( A1 => n14848, A2 => n14690, B1 => n7103, B2 => 
                           n14687, C1 => n14684, C2 => n14592, ZN => n9981);
   U5723 : OAI222_X1 port map( A1 => n14842, A2 => n14690, B1 => n7127, B2 => 
                           n14687, C1 => n14684, C2 => n14586, ZN => n9980);
   U5724 : OAI222_X1 port map( A1 => n14836, A2 => n14690, B1 => n7151, B2 => 
                           n14687, C1 => n14684, C2 => n14580, ZN => n9979);
   U5725 : OAI222_X1 port map( A1 => n14830, A2 => n14690, B1 => n7175, B2 => 
                           n14687, C1 => n14684, C2 => n14574, ZN => n9978);
   U5726 : OAI222_X1 port map( A1 => n14812, A2 => n14689, B1 => n7247, B2 => 
                           n14687, C1 => n14684, C2 => n14556, ZN => n9975);
   U5727 : OAI222_X1 port map( A1 => n14806, A2 => n14689, B1 => n7271, B2 => 
                           n14687, C1 => n14684, C2 => n14550, ZN => n9974);
   U5728 : OAI222_X1 port map( A1 => n14800, A2 => n14689, B1 => n7295, B2 => 
                           n14687, C1 => n14684, C2 => n14544, ZN => n9973);
   U5729 : OAI222_X1 port map( A1 => n14794, A2 => n14689, B1 => n7319, B2 => 
                           n14687, C1 => n14685, C2 => n14538, ZN => n9972);
   U5730 : OAI222_X1 port map( A1 => n14788, A2 => n14689, B1 => n7343, B2 => 
                           n14688, C1 => n14685, C2 => n14532, ZN => n9971);
   U5731 : OAI222_X1 port map( A1 => n14782, A2 => n14689, B1 => n7367, B2 => 
                           n14688, C1 => n14685, C2 => n14526, ZN => n9970);
   U5732 : OAI222_X1 port map( A1 => n14776, A2 => n14689, B1 => n7391, B2 => 
                           n14688, C1 => n14685, C2 => n14520, ZN => n9969);
   U5733 : OAI222_X1 port map( A1 => n14770, A2 => n14689, B1 => n7415, B2 => 
                           n14688, C1 => n14685, C2 => n14514, ZN => n9968);
   U5734 : OAI222_X1 port map( A1 => n14892, A2 => n13260, B1 => n7883, B2 => 
                           n13257, C1 => n14634, C2 => n13254, ZN => n10148);
   U5735 : OAI222_X1 port map( A1 => n14886, A2 => n13260, B1 => n7880, B2 => 
                           n13257, C1 => n14628, C2 => n13254, ZN => n10147);
   U5736 : OAI222_X1 port map( A1 => n14880, A2 => n13260, B1 => n7877, B2 => 
                           n13257, C1 => n14622, C2 => n13254, ZN => n10146);
   U5737 : OAI222_X1 port map( A1 => n14874, A2 => n13260, B1 => n7874, B2 => 
                           n13257, C1 => n14616, C2 => n13254, ZN => n10145);
   U5738 : OAI222_X1 port map( A1 => n14868, A2 => n13260, B1 => n7871, B2 => 
                           n13257, C1 => n14610, C2 => n13254, ZN => n10144);
   U5739 : OAI222_X1 port map( A1 => n14862, A2 => n13260, B1 => n7868, B2 => 
                           n13257, C1 => n14604, C2 => n13254, ZN => n10143);
   U5740 : OAI222_X1 port map( A1 => n14856, A2 => n13260, B1 => n7865, B2 => 
                           n13257, C1 => n14598, C2 => n13254, ZN => n10142);
   U5741 : OAI222_X1 port map( A1 => n14850, A2 => n13260, B1 => n7862, B2 => 
                           n13257, C1 => n14592, C2 => n13254, ZN => n10141);
   U5742 : OAI222_X1 port map( A1 => n14844, A2 => n13260, B1 => n7859, B2 => 
                           n13257, C1 => n14586, C2 => n13254, ZN => n10140);
   U5743 : OAI222_X1 port map( A1 => n14838, A2 => n13260, B1 => n7856, B2 => 
                           n13257, C1 => n14580, C2 => n13254, ZN => n10139);
   U5744 : OAI222_X1 port map( A1 => n14832, A2 => n13260, B1 => n7853, B2 => 
                           n13257, C1 => n14574, C2 => n13254, ZN => n10138);
   U5745 : OAI222_X1 port map( A1 => n14826, A2 => n13260, B1 => n7850, B2 => 
                           n13257, C1 => n14568, C2 => n13254, ZN => n10137);
   U5746 : OAI222_X1 port map( A1 => n14820, A2 => n13259, B1 => n7847, B2 => 
                           n13256, C1 => n14562, C2 => n13254, ZN => n10136);
   U5747 : OAI222_X1 port map( A1 => n14814, A2 => n13259, B1 => n7844, B2 => 
                           n13256, C1 => n14556, C2 => n13253, ZN => n10135);
   U5748 : OAI222_X1 port map( A1 => n14808, A2 => n13259, B1 => n7841, B2 => 
                           n13256, C1 => n14550, C2 => n13253, ZN => n10134);
   U5749 : OAI222_X1 port map( A1 => n14802, A2 => n13259, B1 => n7838, B2 => 
                           n13256, C1 => n14544, C2 => n13253, ZN => n10133);
   U5750 : OAI222_X1 port map( A1 => n14796, A2 => n13259, B1 => n7835, B2 => 
                           n13256, C1 => n14538, C2 => n13253, ZN => n10132);
   U5751 : OAI222_X1 port map( A1 => n14790, A2 => n13259, B1 => n7832, B2 => 
                           n13256, C1 => n14532, C2 => n13253, ZN => n10131);
   U5752 : OAI222_X1 port map( A1 => n14784, A2 => n13259, B1 => n7829, B2 => 
                           n13256, C1 => n14526, C2 => n13253, ZN => n10130);
   U5753 : OAI222_X1 port map( A1 => n14778, A2 => n13259, B1 => n7826, B2 => 
                           n13256, C1 => n14520, C2 => n13253, ZN => n10129);
   U5754 : OAI222_X1 port map( A1 => n14772, A2 => n13259, B1 => n7823, B2 => 
                           n13256, C1 => n14514, C2 => n13253, ZN => n10128);
   U5755 : OAI222_X1 port map( A1 => n14766, A2 => n13259, B1 => n7820, B2 => 
                           n13256, C1 => n14715, C2 => n13253, ZN => n10127);
   U5756 : OAI222_X1 port map( A1 => n14760, A2 => n13259, B1 => n7817, B2 => 
                           n13256, C1 => n14703, C2 => n13253, ZN => n10126);
   U5757 : OAI222_X1 port map( A1 => n14754, A2 => n13259, B1 => n7686, B2 => 
                           n13256, C1 => n14692, C2 => n13253, ZN => n10125);
   U5758 : OAI222_X1 port map( A1 => n14892, A2 => n13269, B1 => n7884, B2 => 
                           n13266, C1 => n14634, C2 => n13263, ZN => n10180);
   U5759 : OAI222_X1 port map( A1 => n14886, A2 => n13269, B1 => n7881, B2 => 
                           n13266, C1 => n14628, C2 => n13263, ZN => n10179);
   U5760 : OAI222_X1 port map( A1 => n14880, A2 => n13269, B1 => n7878, B2 => 
                           n13266, C1 => n14622, C2 => n13263, ZN => n10178);
   U5761 : OAI222_X1 port map( A1 => n14874, A2 => n13269, B1 => n7875, B2 => 
                           n13266, C1 => n14616, C2 => n13263, ZN => n10177);
   U5762 : OAI222_X1 port map( A1 => n14868, A2 => n13269, B1 => n7872, B2 => 
                           n13266, C1 => n14610, C2 => n13263, ZN => n10176);
   U5763 : OAI222_X1 port map( A1 => n14862, A2 => n13269, B1 => n7869, B2 => 
                           n13266, C1 => n14604, C2 => n13263, ZN => n10175);
   U5764 : OAI222_X1 port map( A1 => n14856, A2 => n13269, B1 => n7866, B2 => 
                           n13266, C1 => n14598, C2 => n13263, ZN => n10174);
   U5765 : OAI222_X1 port map( A1 => n14850, A2 => n13269, B1 => n7863, B2 => 
                           n13266, C1 => n14592, C2 => n13263, ZN => n10173);
   U5766 : OAI222_X1 port map( A1 => n14844, A2 => n13269, B1 => n7860, B2 => 
                           n13266, C1 => n14586, C2 => n13263, ZN => n10172);
   U5767 : OAI222_X1 port map( A1 => n14838, A2 => n13269, B1 => n7857, B2 => 
                           n13266, C1 => n14580, C2 => n13263, ZN => n10171);
   U5768 : OAI222_X1 port map( A1 => n14832, A2 => n13269, B1 => n7854, B2 => 
                           n13266, C1 => n14574, C2 => n13263, ZN => n10170);
   U5769 : OAI222_X1 port map( A1 => n14826, A2 => n13269, B1 => n7851, B2 => 
                           n13266, C1 => n14568, C2 => n13263, ZN => n10169);
   U5770 : OAI222_X1 port map( A1 => n14820, A2 => n13268, B1 => n7848, B2 => 
                           n13265, C1 => n14562, C2 => n13263, ZN => n10168);
   U5771 : OAI222_X1 port map( A1 => n14814, A2 => n13268, B1 => n7845, B2 => 
                           n13265, C1 => n14556, C2 => n13262, ZN => n10167);
   U5772 : OAI222_X1 port map( A1 => n14808, A2 => n13268, B1 => n7842, B2 => 
                           n13265, C1 => n14550, C2 => n13262, ZN => n10166);
   U5773 : OAI222_X1 port map( A1 => n14802, A2 => n13268, B1 => n7839, B2 => 
                           n13265, C1 => n14544, C2 => n13262, ZN => n10165);
   U5774 : OAI222_X1 port map( A1 => n14796, A2 => n13268, B1 => n7836, B2 => 
                           n13265, C1 => n14538, C2 => n13262, ZN => n10164);
   U5775 : OAI222_X1 port map( A1 => n14790, A2 => n13268, B1 => n7833, B2 => 
                           n13265, C1 => n14532, C2 => n13262, ZN => n10163);
   U5776 : OAI222_X1 port map( A1 => n14784, A2 => n13268, B1 => n7830, B2 => 
                           n13265, C1 => n14526, C2 => n13262, ZN => n10162);
   U5777 : OAI222_X1 port map( A1 => n14778, A2 => n13268, B1 => n7827, B2 => 
                           n13265, C1 => n14520, C2 => n13262, ZN => n10161);
   U5778 : OAI222_X1 port map( A1 => n14772, A2 => n13268, B1 => n7824, B2 => 
                           n13265, C1 => n14514, C2 => n13262, ZN => n10160);
   U5779 : OAI222_X1 port map( A1 => n14766, A2 => n13268, B1 => n7821, B2 => 
                           n13265, C1 => n14715, C2 => n13262, ZN => n10159);
   U5780 : OAI222_X1 port map( A1 => n14760, A2 => n13268, B1 => n7818, B2 => 
                           n13265, C1 => n14703, C2 => n13262, ZN => n10158);
   U5781 : OAI222_X1 port map( A1 => n14883, A2 => n13620, B1 => n6944, B2 => 
                           n13617, C1 => n14625, C2 => n13614, ZN => n11427);
   U5782 : OAI222_X1 port map( A1 => n14877, A2 => n13620, B1 => n6968, B2 => 
                           n13617, C1 => n14619, C2 => n13614, ZN => n11426);
   U5783 : OAI222_X1 port map( A1 => n14871, A2 => n13620, B1 => n6992, B2 => 
                           n13617, C1 => n14613, C2 => n13614, ZN => n11425);
   U5784 : OAI222_X1 port map( A1 => n14865, A2 => n13620, B1 => n7016, B2 => 
                           n13617, C1 => n14607, C2 => n13614, ZN => n11424);
   U5785 : OAI222_X1 port map( A1 => n14859, A2 => n13620, B1 => n7040, B2 => 
                           n13617, C1 => n14601, C2 => n13614, ZN => n11423);
   U5786 : OAI222_X1 port map( A1 => n14853, A2 => n13620, B1 => n7064, B2 => 
                           n13617, C1 => n14595, C2 => n13614, ZN => n11422);
   U5787 : OAI222_X1 port map( A1 => n14847, A2 => n13620, B1 => n7088, B2 => 
                           n13617, C1 => n14589, C2 => n13614, ZN => n11421);
   U5788 : OAI222_X1 port map( A1 => n14841, A2 => n13620, B1 => n7112, B2 => 
                           n13617, C1 => n14583, C2 => n13614, ZN => n11420);
   U5789 : OAI222_X1 port map( A1 => n14835, A2 => n13620, B1 => n7136, B2 => 
                           n13617, C1 => n14577, C2 => n13614, ZN => n11419);
   U5790 : OAI222_X1 port map( A1 => n14829, A2 => n13620, B1 => n7160, B2 => 
                           n13617, C1 => n14571, C2 => n13614, ZN => n11418);
   U5791 : OAI222_X1 port map( A1 => n14823, A2 => n13620, B1 => n7184, B2 => 
                           n13617, C1 => n14565, C2 => n13614, ZN => n11417);
   U5792 : OAI222_X1 port map( A1 => n14805, A2 => n13619, B1 => n7256, B2 => 
                           n13616, C1 => n14547, C2 => n13613, ZN => n11414);
   U5793 : OAI222_X1 port map( A1 => n14799, A2 => n13619, B1 => n7280, B2 => 
                           n13616, C1 => n14541, C2 => n13613, ZN => n11413);
   U5794 : OAI222_X1 port map( A1 => n14793, A2 => n13619, B1 => n7304, B2 => 
                           n13616, C1 => n14535, C2 => n13613, ZN => n11412);
   U5795 : OAI222_X1 port map( A1 => n14787, A2 => n13619, B1 => n7328, B2 => 
                           n13616, C1 => n14529, C2 => n13613, ZN => n11411);
   U5796 : OAI222_X1 port map( A1 => n14781, A2 => n13619, B1 => n7352, B2 => 
                           n13616, C1 => n14523, C2 => n13613, ZN => n11410);
   U5797 : OAI222_X1 port map( A1 => n14775, A2 => n13619, B1 => n7376, B2 => 
                           n13616, C1 => n14517, C2 => n13613, ZN => n11409);
   U5798 : OAI222_X1 port map( A1 => n14769, A2 => n13619, B1 => n7400, B2 => 
                           n13616, C1 => n14511, C2 => n13613, ZN => n11408);
   U5799 : OAI222_X1 port map( A1 => n14763, A2 => n13619, B1 => n7424, B2 => 
                           n13616, C1 => n14712, C2 => n13613, ZN => n11407);
   U5800 : OAI222_X1 port map( A1 => n14757, A2 => n13619, B1 => n7448, B2 => 
                           n13616, C1 => n14700, C2 => n13613, ZN => n11406);
   U5801 : OAI222_X1 port map( A1 => n14751, A2 => n13619, B1 => n7472, B2 => 
                           n13616, C1 => n14695, C2 => n13613, ZN => n11405);
   U5802 : OAI222_X1 port map( A1 => n14829, A2 => n13629, B1 => n7159, B2 => 
                           n13626, C1 => n14571, C2 => n13623, ZN => n11450);
   U5803 : OAI222_X1 port map( A1 => n14823, A2 => n13629, B1 => n7183, B2 => 
                           n13626, C1 => n14565, C2 => n13623, ZN => n11449);
   U5804 : OAI222_X1 port map( A1 => n14805, A2 => n13628, B1 => n7255, B2 => 
                           n13625, C1 => n14547, C2 => n13622, ZN => n11446);
   U5805 : OAI222_X1 port map( A1 => n14799, A2 => n13628, B1 => n7279, B2 => 
                           n13625, C1 => n14541, C2 => n13622, ZN => n11445);
   U5806 : OAI222_X1 port map( A1 => n14793, A2 => n13628, B1 => n7303, B2 => 
                           n13625, C1 => n14535, C2 => n13622, ZN => n11444);
   U5807 : OAI222_X1 port map( A1 => n14787, A2 => n13628, B1 => n7327, B2 => 
                           n13625, C1 => n14529, C2 => n13622, ZN => n11443);
   U5808 : OAI222_X1 port map( A1 => n14781, A2 => n13628, B1 => n7351, B2 => 
                           n13625, C1 => n14523, C2 => n13622, ZN => n11442);
   U5809 : OAI222_X1 port map( A1 => n14775, A2 => n13628, B1 => n7375, B2 => 
                           n13625, C1 => n14517, C2 => n13622, ZN => n11441);
   U5810 : OAI222_X1 port map( A1 => n14769, A2 => n13628, B1 => n7399, B2 => 
                           n13625, C1 => n14511, C2 => n13622, ZN => n11440);
   U5811 : OAI222_X1 port map( A1 => n14763, A2 => n13628, B1 => n7423, B2 => 
                           n13625, C1 => n14712, C2 => n13622, ZN => n11439);
   U5812 : OAI222_X1 port map( A1 => n14757, A2 => n13628, B1 => n7447, B2 => 
                           n13625, C1 => n14700, C2 => n13622, ZN => n11438);
   U5813 : OAI222_X1 port map( A1 => n14751, A2 => n13628, B1 => n7471, B2 => 
                           n13625, C1 => n14695, C2 => n13622, ZN => n11437);
   U5814 : OAI222_X1 port map( A1 => n14883, A2 => n14316, B1 => n7630, B2 => 
                           n14312, C1 => n14624, C2 => n14310, ZN => n9283);
   U5815 : OAI222_X1 port map( A1 => n14877, A2 => n14316, B1 => n7624, B2 => 
                           n14312, C1 => n14618, C2 => n14310, ZN => n9282);
   U5816 : OAI222_X1 port map( A1 => n14871, A2 => n14316, B1 => n7618, B2 => 
                           n14312, C1 => n14612, C2 => n14310, ZN => n9281);
   U5817 : OAI222_X1 port map( A1 => n14865, A2 => n14316, B1 => n7612, B2 => 
                           n14313, C1 => n14606, C2 => n14310, ZN => n9280);
   U5818 : OAI222_X1 port map( A1 => n14859, A2 => n14316, B1 => n7606, B2 => 
                           n14313, C1 => n14600, C2 => n14310, ZN => n9279);
   U5819 : OAI222_X1 port map( A1 => n14853, A2 => n14316, B1 => n7600, B2 => 
                           n14313, C1 => n14594, C2 => n14310, ZN => n9278);
   U5820 : OAI222_X1 port map( A1 => n14847, A2 => n14316, B1 => n7594, B2 => 
                           n14313, C1 => n14588, C2 => n14310, ZN => n9277);
   U5821 : OAI222_X1 port map( A1 => n14841, A2 => n14316, B1 => n7588, B2 => 
                           n14313, C1 => n14582, C2 => n14310, ZN => n9276);
   U5822 : OAI222_X1 port map( A1 => n14835, A2 => n14316, B1 => n7582, B2 => 
                           n14313, C1 => n14576, C2 => n14310, ZN => n9275);
   U5823 : OAI222_X1 port map( A1 => n14829, A2 => n14316, B1 => n7576, B2 => 
                           n14313, C1 => n14570, C2 => n14310, ZN => n9274);
   U5824 : OAI222_X1 port map( A1 => n14817, A2 => n14315, B1 => n7564, B2 => 
                           n14313, C1 => n14558, C2 => n14310, ZN => n9272);
   U5825 : OAI222_X1 port map( A1 => n14811, A2 => n14315, B1 => n7558, B2 => 
                           n14313, C1 => n14552, C2 => n14309, ZN => n9271);
   U5826 : OAI222_X1 port map( A1 => n14805, A2 => n14315, B1 => n7552, B2 => 
                           n14313, C1 => n14546, C2 => n14309, ZN => n9270);
   U5827 : OAI222_X1 port map( A1 => n14799, A2 => n14315, B1 => n7546, B2 => 
                           n14313, C1 => n14540, C2 => n14309, ZN => n9269);
   U5828 : OAI222_X1 port map( A1 => n14793, A2 => n14315, B1 => n7540, B2 => 
                           n14313, C1 => n14534, C2 => n14309, ZN => n9268);
   U5829 : OAI222_X1 port map( A1 => n14787, A2 => n14315, B1 => n7534, B2 => 
                           n14314, C1 => n14528, C2 => n14309, ZN => n9267);
   U5830 : OAI222_X1 port map( A1 => n14781, A2 => n14315, B1 => n7528, B2 => 
                           n14314, C1 => n14522, C2 => n14309, ZN => n9266);
   U5831 : OAI222_X1 port map( A1 => n14775, A2 => n14315, B1 => n7522, B2 => 
                           n14314, C1 => n14516, C2 => n14309, ZN => n9265);
   U5832 : OAI222_X1 port map( A1 => n14768, A2 => n14315, B1 => n7516, B2 => 
                           n14314, C1 => n14510, C2 => n14309, ZN => n9264);
   U5833 : OAI222_X1 port map( A1 => n14763, A2 => n14315, B1 => n7510, B2 => 
                           n14314, C1 => n14711, C2 => n14309, ZN => n9263);
   U5834 : OAI222_X1 port map( A1 => n14757, A2 => n14315, B1 => n7504, B2 => 
                           n14314, C1 => n14699, C2 => n14309, ZN => n9262);
   U5835 : OAI222_X1 port map( A1 => n14751, A2 => n14315, B1 => n7498, B2 => 
                           n14312, C1 => n14696, C2 => n14309, ZN => n9261);
   U5836 : OAI222_X1 port map( A1 => n14882, A2 => n14399, B1 => n7628, B2 => 
                           n14395, C1 => n14624, C2 => n14393, ZN => n9571);
   U5837 : OAI222_X1 port map( A1 => n14876, A2 => n14399, B1 => n7622, B2 => 
                           n14395, C1 => n14618, C2 => n14393, ZN => n9570);
   U5838 : OAI222_X1 port map( A1 => n14870, A2 => n14399, B1 => n7616, B2 => 
                           n14395, C1 => n14612, C2 => n14393, ZN => n9569);
   U5839 : OAI222_X1 port map( A1 => n14864, A2 => n14399, B1 => n7610, B2 => 
                           n14396, C1 => n14606, C2 => n14393, ZN => n9568);
   U5840 : OAI222_X1 port map( A1 => n14858, A2 => n14399, B1 => n7604, B2 => 
                           n14396, C1 => n14600, C2 => n14393, ZN => n9567);
   U5841 : OAI222_X1 port map( A1 => n14852, A2 => n14399, B1 => n7598, B2 => 
                           n14396, C1 => n14594, C2 => n14393, ZN => n9566);
   U5842 : OAI222_X1 port map( A1 => n14846, A2 => n14399, B1 => n7592, B2 => 
                           n14396, C1 => n14588, C2 => n14393, ZN => n9565);
   U5843 : OAI222_X1 port map( A1 => n14840, A2 => n14399, B1 => n7586, B2 => 
                           n14396, C1 => n14582, C2 => n14393, ZN => n9564);
   U5844 : OAI222_X1 port map( A1 => n14834, A2 => n14399, B1 => n7580, B2 => 
                           n14396, C1 => n14576, C2 => n14393, ZN => n9563);
   U5845 : OAI222_X1 port map( A1 => n14828, A2 => n14399, B1 => n7574, B2 => 
                           n14396, C1 => n14570, C2 => n14393, ZN => n9562);
   U5846 : OAI222_X1 port map( A1 => n14816, A2 => n14398, B1 => n7562, B2 => 
                           n14396, C1 => n14558, C2 => n14393, ZN => n9560);
   U5847 : OAI222_X1 port map( A1 => n14810, A2 => n14398, B1 => n7556, B2 => 
                           n14396, C1 => n14552, C2 => n14392, ZN => n9559);
   U5848 : OAI222_X1 port map( A1 => n14804, A2 => n14398, B1 => n7550, B2 => 
                           n14396, C1 => n14546, C2 => n14392, ZN => n9558);
   U5849 : OAI222_X1 port map( A1 => n14798, A2 => n14398, B1 => n7544, B2 => 
                           n14396, C1 => n14540, C2 => n14392, ZN => n9557);
   U5850 : OAI222_X1 port map( A1 => n14792, A2 => n14398, B1 => n7538, B2 => 
                           n14396, C1 => n14534, C2 => n14392, ZN => n9556);
   U5851 : OAI222_X1 port map( A1 => n14786, A2 => n14398, B1 => n7532, B2 => 
                           n14397, C1 => n14528, C2 => n14392, ZN => n9555);
   U5852 : OAI222_X1 port map( A1 => n14780, A2 => n14398, B1 => n7526, B2 => 
                           n14397, C1 => n14522, C2 => n14392, ZN => n9554);
   U5853 : OAI222_X1 port map( A1 => n14774, A2 => n14398, B1 => n7520, B2 => 
                           n14397, C1 => n14516, C2 => n14392, ZN => n9553);
   U5854 : OAI222_X1 port map( A1 => n14768, A2 => n14398, B1 => n7514, B2 => 
                           n14397, C1 => n14510, C2 => n14392, ZN => n9552);
   U5855 : OAI222_X1 port map( A1 => n14762, A2 => n14398, B1 => n7508, B2 => 
                           n14397, C1 => n14711, C2 => n14392, ZN => n9551);
   U5856 : OAI222_X1 port map( A1 => n14756, A2 => n14398, B1 => n7502, B2 => 
                           n14397, C1 => n14699, C2 => n14392, ZN => n9550);
   U5857 : OAI222_X1 port map( A1 => n14750, A2 => n14398, B1 => n7496, B2 => 
                           n14395, C1 => n14696, C2 => n14392, ZN => n9549);
   U5858 : OAI222_X1 port map( A1 => n14750, A2 => n14434, B1 => n7490, B2 => 
                           n14431, C1 => n14697, C2 => n14428, ZN => n9677);
   U5859 : OAI222_X1 port map( A1 => n14938, A2 => n14691, B1 => n6743, B2 => 
                           n14687, C1 => n14683, C2 => n14682, ZN => n9996);
   U5860 : OAI222_X1 port map( A1 => n14932, A2 => n14691, B1 => n6767, B2 => 
                           n14686, C1 => n14683, C2 => n14676, ZN => n9995);
   U5861 : OAI222_X1 port map( A1 => n14926, A2 => n14691, B1 => n6791, B2 => 
                           n14686, C1 => n14683, C2 => n14670, ZN => n9994);
   U5862 : OAI222_X1 port map( A1 => n14920, A2 => n14691, B1 => n6815, B2 => 
                           n14686, C1 => n14683, C2 => n14664, ZN => n9993);
   U5863 : OAI222_X1 port map( A1 => n14914, A2 => n14691, B1 => n6839, B2 => 
                           n14686, C1 => n14683, C2 => n14658, ZN => n9992);
   U5864 : OAI222_X1 port map( A1 => n14908, A2 => n14691, B1 => n6863, B2 => 
                           n14686, C1 => n14683, C2 => n14652, ZN => n9991);
   U5865 : OAI222_X1 port map( A1 => n14902, A2 => n14691, B1 => n6887, B2 => 
                           n14686, C1 => n14683, C2 => n14646, ZN => n9990);
   U5866 : OAI222_X1 port map( A1 => n14896, A2 => n14691, B1 => n6911, B2 => 
                           n14686, C1 => n14684, C2 => n14640, ZN => n9989);
   U5867 : OAI222_X1 port map( A1 => n14767, A2 => n14497, B1 => n14496, B2 => 
                           n1709, C1 => n14509, C2 => n14491, ZN => n9904);
   U5868 : OAI222_X1 port map( A1 => n14767, A2 => n14506, B1 => n14505, B2 => 
                           n1708, C1 => n14509, C2 => n14500, ZN => n9936);
   U5869 : OAI222_X1 port map( A1 => n14821, A2 => n14471, B1 => n820, B2 => 
                           n14469, C1 => n14563, C2 => n14465, ZN => n9817);
   U5870 : OAI222_X1 port map( A1 => n14815, A2 => n14470, B1 => n756, B2 => 
                           n14469, C1 => n14557, C2 => n14465, ZN => n9816);
   U5871 : OAI222_X1 port map( A1 => n14881, A2 => n14498, B1 => n14494, B2 => 
                           n1648, C1 => n14623, C2 => n14492, ZN => n9923);
   U5872 : OAI222_X1 port map( A1 => n14875, A2 => n14498, B1 => n14494, B2 => 
                           n1647, C1 => n14617, C2 => n14492, ZN => n9922);
   U5873 : OAI222_X1 port map( A1 => n14869, A2 => n14498, B1 => n14494, B2 => 
                           n1646, C1 => n14611, C2 => n14492, ZN => n9921);
   U5874 : OAI222_X1 port map( A1 => n14863, A2 => n14498, B1 => n14495, B2 => 
                           n1645, C1 => n14605, C2 => n14492, ZN => n9920);
   U5875 : OAI222_X1 port map( A1 => n14833, A2 => n14498, B1 => n14495, B2 => 
                           n1640, C1 => n14575, C2 => n14492, ZN => n9915);
   U5876 : OAI222_X1 port map( A1 => n14827, A2 => n14498, B1 => n14495, B2 => 
                           n1639, C1 => n14569, C2 => n14492, ZN => n9914);
   U5877 : OAI222_X1 port map( A1 => n14821, A2 => n14498, B1 => n823, B2 => 
                           n14496, C1 => n14563, C2 => n14492, ZN => n9913);
   U5878 : OAI222_X1 port map( A1 => n14809, A2 => n14497, B1 => n14495, B2 => 
                           n1636, C1 => n14551, C2 => n14491, ZN => n9911);
   U5879 : OAI222_X1 port map( A1 => n14803, A2 => n14497, B1 => n14495, B2 => 
                           n1635, C1 => n14545, C2 => n14491, ZN => n9910);
   U5880 : OAI222_X1 port map( A1 => n14797, A2 => n14497, B1 => n14495, B2 => 
                           n1634, C1 => n14539, C2 => n14491, ZN => n9909);
   U5881 : OAI222_X1 port map( A1 => n14791, A2 => n14497, B1 => n14496, B2 => 
                           n1633, C1 => n14533, C2 => n14491, ZN => n9908);
   U5882 : OAI222_X1 port map( A1 => n14785, A2 => n14497, B1 => n14496, B2 => 
                           n1632, C1 => n14527, C2 => n14491, ZN => n9907);
   U5883 : OAI222_X1 port map( A1 => n14779, A2 => n14497, B1 => n14496, B2 => 
                           n1631, C1 => n14521, C2 => n14491, ZN => n9906);
   U5884 : OAI222_X1 port map( A1 => n14773, A2 => n14497, B1 => n14496, B2 => 
                           n1630, C1 => n14515, C2 => n14491, ZN => n9905);
   U5885 : OAI222_X1 port map( A1 => n14749, A2 => n14497, B1 => n14494, B2 => 
                           n1629, C1 => n14697, C2 => n14491, ZN => n9901);
   U5886 : OAI222_X1 port map( A1 => n14881, A2 => n14507, B1 => n14503, B2 => 
                           n1627, C1 => n14623, C2 => n14501, ZN => n9955);
   U5887 : OAI222_X1 port map( A1 => n14875, A2 => n14507, B1 => n14503, B2 => 
                           n1626, C1 => n14617, C2 => n14501, ZN => n9954);
   U5888 : OAI222_X1 port map( A1 => n14869, A2 => n14507, B1 => n14503, B2 => 
                           n1625, C1 => n14611, C2 => n14501, ZN => n9953);
   U5889 : OAI222_X1 port map( A1 => n14863, A2 => n14507, B1 => n14504, B2 => 
                           n1624, C1 => n14605, C2 => n14501, ZN => n9952);
   U5890 : OAI222_X1 port map( A1 => n14833, A2 => n14507, B1 => n14504, B2 => 
                           n1619, C1 => n14575, C2 => n14501, ZN => n9947);
   U5891 : OAI222_X1 port map( A1 => n14827, A2 => n14507, B1 => n14504, B2 => 
                           n1618, C1 => n14569, C2 => n14501, ZN => n9946);
   U5892 : OAI222_X1 port map( A1 => n14821, A2 => n14507, B1 => n824, B2 => 
                           n14505, C1 => n14563, C2 => n14501, ZN => n9945);
   U5893 : OAI222_X1 port map( A1 => n14809, A2 => n14506, B1 => n14504, B2 => 
                           n1615, C1 => n14551, C2 => n14500, ZN => n9943);
   U5894 : OAI222_X1 port map( A1 => n14803, A2 => n14506, B1 => n14504, B2 => 
                           n1614, C1 => n14545, C2 => n14500, ZN => n9942);
   U5895 : OAI222_X1 port map( A1 => n14797, A2 => n14506, B1 => n14504, B2 => 
                           n1613, C1 => n14539, C2 => n14500, ZN => n9941);
   U5896 : OAI222_X1 port map( A1 => n14791, A2 => n14506, B1 => n14505, B2 => 
                           n1612, C1 => n14533, C2 => n14500, ZN => n9940);
   U5897 : OAI222_X1 port map( A1 => n14785, A2 => n14506, B1 => n14505, B2 => 
                           n1611, C1 => n14527, C2 => n14500, ZN => n9939);
   U5898 : OAI222_X1 port map( A1 => n14779, A2 => n14506, B1 => n14505, B2 => 
                           n1610, C1 => n14521, C2 => n14500, ZN => n9938);
   U5899 : OAI222_X1 port map( A1 => n14773, A2 => n14506, B1 => n14505, B2 => 
                           n1609, C1 => n14515, C2 => n14500, ZN => n9937);
   U5900 : OAI222_X1 port map( A1 => n14749, A2 => n14506, B1 => n14503, B2 => 
                           n1608, C1 => n14697, C2 => n14500, ZN => n9933);
   U5901 : OAI222_X1 port map( A1 => n14761, A2 => n14497, B1 => n14496, B2 => 
                           n1602, C1 => n14710, C2 => n14491, ZN => n9903);
   U5902 : OAI222_X1 port map( A1 => n14755, A2 => n14497, B1 => n14496, B2 => 
                           n1601, C1 => n14698, C2 => n14491, ZN => n9902);
   U5903 : OAI222_X1 port map( A1 => n14761, A2 => n14506, B1 => n14505, B2 => 
                           n1600, C1 => n14710, C2 => n14500, ZN => n9935);
   U5904 : OAI222_X1 port map( A1 => n14755, A2 => n14506, B1 => n14505, B2 => 
                           n1599, C1 => n14698, C2 => n14500, ZN => n9934);
   U5905 : OAI222_X1 port map( A1 => n14892, A2 => n13287, B1 => n1598, B2 => 
                           n13284, C1 => n14634, C2 => n13281, ZN => n10244);
   U5906 : OAI222_X1 port map( A1 => n14886, A2 => n13287, B1 => n1597, B2 => 
                           n13284, C1 => n14628, C2 => n13281, ZN => n10243);
   U5907 : OAI222_X1 port map( A1 => n14880, A2 => n13287, B1 => n1596, B2 => 
                           n13284, C1 => n14622, C2 => n13281, ZN => n10242);
   U5908 : OAI222_X1 port map( A1 => n14874, A2 => n13287, B1 => n1595, B2 => 
                           n13284, C1 => n14616, C2 => n13281, ZN => n10241);
   U5909 : OAI222_X1 port map( A1 => n14868, A2 => n13287, B1 => n1594, B2 => 
                           n13284, C1 => n14610, C2 => n13281, ZN => n10240);
   U5910 : OAI222_X1 port map( A1 => n14862, A2 => n13287, B1 => n1593, B2 => 
                           n13284, C1 => n14604, C2 => n13281, ZN => n10239);
   U5911 : OAI222_X1 port map( A1 => n14856, A2 => n13287, B1 => n1592, B2 => 
                           n13284, C1 => n14598, C2 => n13281, ZN => n10238);
   U5912 : OAI222_X1 port map( A1 => n14850, A2 => n13287, B1 => n1591, B2 => 
                           n13284, C1 => n14592, C2 => n13281, ZN => n10237);
   U5913 : OAI222_X1 port map( A1 => n14844, A2 => n13287, B1 => n1590, B2 => 
                           n13284, C1 => n14586, C2 => n13281, ZN => n10236);
   U5914 : OAI222_X1 port map( A1 => n14838, A2 => n13287, B1 => n1589, B2 => 
                           n13284, C1 => n14580, C2 => n13281, ZN => n10235);
   U5915 : OAI222_X1 port map( A1 => n14832, A2 => n13287, B1 => n1588, B2 => 
                           n13284, C1 => n14574, C2 => n13281, ZN => n10234);
   U5916 : OAI222_X1 port map( A1 => n14826, A2 => n13287, B1 => n1587, B2 => 
                           n13284, C1 => n14568, C2 => n13281, ZN => n10233);
   U5917 : OAI222_X1 port map( A1 => n14820, A2 => n13286, B1 => n1586, B2 => 
                           n13283, C1 => n14562, C2 => n13281, ZN => n10232);
   U5918 : OAI222_X1 port map( A1 => n14814, A2 => n13286, B1 => n1585, B2 => 
                           n13283, C1 => n14556, C2 => n13280, ZN => n10231);
   U5919 : OAI222_X1 port map( A1 => n14808, A2 => n13286, B1 => n1584, B2 => 
                           n13283, C1 => n14550, C2 => n13280, ZN => n10230);
   U5920 : OAI222_X1 port map( A1 => n14802, A2 => n13286, B1 => n1583, B2 => 
                           n13283, C1 => n14544, C2 => n13280, ZN => n10229);
   U5921 : OAI222_X1 port map( A1 => n14796, A2 => n13286, B1 => n1582, B2 => 
                           n13283, C1 => n14538, C2 => n13280, ZN => n10228);
   U5922 : OAI222_X1 port map( A1 => n14790, A2 => n13286, B1 => n1581, B2 => 
                           n13283, C1 => n14532, C2 => n13280, ZN => n10227);
   U5923 : OAI222_X1 port map( A1 => n14784, A2 => n13286, B1 => n1580, B2 => 
                           n13283, C1 => n14526, C2 => n13280, ZN => n10226);
   U5924 : OAI222_X1 port map( A1 => n14778, A2 => n13286, B1 => n1579, B2 => 
                           n13283, C1 => n14520, C2 => n13280, ZN => n10225);
   U5925 : OAI222_X1 port map( A1 => n14772, A2 => n13286, B1 => n1578, B2 => 
                           n13283, C1 => n14514, C2 => n13280, ZN => n10224);
   U5926 : OAI222_X1 port map( A1 => n14766, A2 => n13286, B1 => n1577, B2 => 
                           n13283, C1 => n14715, C2 => n13280, ZN => n10223);
   U5927 : OAI222_X1 port map( A1 => n14760, A2 => n13286, B1 => n1576, B2 => 
                           n13283, C1 => n14703, C2 => n13280, ZN => n10222);
   U5928 : OAI222_X1 port map( A1 => n14754, A2 => n13286, B1 => n1575, B2 => 
                           n13283, C1 => n14692, C2 => n13280, ZN => n10221);
   U5929 : OAI222_X1 port map( A1 => n14885, A2 => n13359, B1 => n1509, B2 => 
                           n13356, C1 => n14627, C2 => n13353, ZN => n10499);
   U5930 : OAI222_X1 port map( A1 => n14879, A2 => n13359, B1 => n1508, B2 => 
                           n13356, C1 => n14621, C2 => n13353, ZN => n10498);
   U5931 : OAI222_X1 port map( A1 => n14873, A2 => n13359, B1 => n1507, B2 => 
                           n13356, C1 => n14615, C2 => n13353, ZN => n10497);
   U5932 : OAI222_X1 port map( A1 => n14867, A2 => n13359, B1 => n1506, B2 => 
                           n13356, C1 => n14609, C2 => n13353, ZN => n10496);
   U5933 : OAI222_X1 port map( A1 => n14861, A2 => n13359, B1 => n1505, B2 => 
                           n13356, C1 => n14603, C2 => n13353, ZN => n10495);
   U5934 : OAI222_X1 port map( A1 => n14855, A2 => n13359, B1 => n1504, B2 => 
                           n13356, C1 => n14597, C2 => n13353, ZN => n10494);
   U5935 : OAI222_X1 port map( A1 => n14849, A2 => n13359, B1 => n1503, B2 => 
                           n13356, C1 => n14591, C2 => n13353, ZN => n10493);
   U5936 : OAI222_X1 port map( A1 => n14843, A2 => n13359, B1 => n1502, B2 => 
                           n13356, C1 => n14585, C2 => n13353, ZN => n10492);
   U5937 : OAI222_X1 port map( A1 => n14837, A2 => n13359, B1 => n1501, B2 => 
                           n13356, C1 => n14579, C2 => n13353, ZN => n10491);
   U5938 : OAI222_X1 port map( A1 => n14831, A2 => n13359, B1 => n1500, B2 => 
                           n13356, C1 => n14573, C2 => n13353, ZN => n10490);
   U5939 : OAI222_X1 port map( A1 => n14825, A2 => n13359, B1 => n1499, B2 => 
                           n13356, C1 => n14567, C2 => n13353, ZN => n10489);
   U5940 : OAI222_X1 port map( A1 => n14819, A2 => n13358, B1 => n1498, B2 => 
                           n13355, C1 => n14561, C2 => n13353, ZN => n10488);
   U5941 : OAI222_X1 port map( A1 => n14813, A2 => n13358, B1 => n1497, B2 => 
                           n13355, C1 => n14555, C2 => n13352, ZN => n10487);
   U5942 : OAI222_X1 port map( A1 => n14807, A2 => n13358, B1 => n1496, B2 => 
                           n13355, C1 => n14549, C2 => n13352, ZN => n10486);
   U5943 : OAI222_X1 port map( A1 => n14801, A2 => n13358, B1 => n1495, B2 => 
                           n13355, C1 => n14543, C2 => n13352, ZN => n10485);
   U5944 : OAI222_X1 port map( A1 => n14795, A2 => n13358, B1 => n1494, B2 => 
                           n13355, C1 => n14537, C2 => n13352, ZN => n10484);
   U5945 : OAI222_X1 port map( A1 => n14789, A2 => n13358, B1 => n1493, B2 => 
                           n13355, C1 => n14531, C2 => n13352, ZN => n10483);
   U5946 : OAI222_X1 port map( A1 => n14783, A2 => n13358, B1 => n1492, B2 => 
                           n13355, C1 => n14525, C2 => n13352, ZN => n10482);
   U5947 : OAI222_X1 port map( A1 => n14777, A2 => n13358, B1 => n1491, B2 => 
                           n13355, C1 => n14519, C2 => n13352, ZN => n10481);
   U5948 : OAI222_X1 port map( A1 => n14771, A2 => n13358, B1 => n1490, B2 => 
                           n13355, C1 => n14513, C2 => n13352, ZN => n10480);
   U5949 : OAI222_X1 port map( A1 => n14765, A2 => n13358, B1 => n1489, B2 => 
                           n13355, C1 => n14714, C2 => n13352, ZN => n10479);
   U5950 : OAI222_X1 port map( A1 => n14759, A2 => n13358, B1 => n1488, B2 => 
                           n13355, C1 => n14702, C2 => n13352, ZN => n10478);
   U5951 : OAI222_X1 port map( A1 => n14753, A2 => n13358, B1 => n1487, B2 => 
                           n13355, C1 => n14693, C2 => n13352, ZN => n10477);
   U5952 : OAI222_X1 port map( A1 => n14885, A2 => n13368, B1 => n1485, B2 => 
                           n13365, C1 => n14627, C2 => n13362, ZN => n10531);
   U5953 : OAI222_X1 port map( A1 => n14879, A2 => n13368, B1 => n1484, B2 => 
                           n13365, C1 => n14621, C2 => n13362, ZN => n10530);
   U5954 : OAI222_X1 port map( A1 => n14873, A2 => n13368, B1 => n1483, B2 => 
                           n13365, C1 => n14615, C2 => n13362, ZN => n10529);
   U5955 : OAI222_X1 port map( A1 => n14867, A2 => n13368, B1 => n1482, B2 => 
                           n13365, C1 => n14609, C2 => n13362, ZN => n10528);
   U5956 : OAI222_X1 port map( A1 => n14861, A2 => n13368, B1 => n1481, B2 => 
                           n13365, C1 => n14603, C2 => n13362, ZN => n10527);
   U5957 : OAI222_X1 port map( A1 => n14855, A2 => n13368, B1 => n1480, B2 => 
                           n13365, C1 => n14597, C2 => n13362, ZN => n10526);
   U5958 : OAI222_X1 port map( A1 => n14849, A2 => n13368, B1 => n1479, B2 => 
                           n13365, C1 => n14591, C2 => n13362, ZN => n10525);
   U5959 : OAI222_X1 port map( A1 => n14843, A2 => n13368, B1 => n1478, B2 => 
                           n13365, C1 => n14585, C2 => n13362, ZN => n10524);
   U5960 : OAI222_X1 port map( A1 => n14837, A2 => n13368, B1 => n1477, B2 => 
                           n13365, C1 => n14579, C2 => n13362, ZN => n10523);
   U5961 : OAI222_X1 port map( A1 => n14831, A2 => n13368, B1 => n1476, B2 => 
                           n13365, C1 => n14573, C2 => n13362, ZN => n10522);
   U5962 : OAI222_X1 port map( A1 => n14825, A2 => n13368, B1 => n1475, B2 => 
                           n13365, C1 => n14567, C2 => n13362, ZN => n10521);
   U5963 : OAI222_X1 port map( A1 => n14819, A2 => n13367, B1 => n1474, B2 => 
                           n13364, C1 => n14561, C2 => n13362, ZN => n10520);
   U5964 : OAI222_X1 port map( A1 => n14813, A2 => n13367, B1 => n1473, B2 => 
                           n13364, C1 => n14555, C2 => n13361, ZN => n10519);
   U5965 : OAI222_X1 port map( A1 => n14807, A2 => n13367, B1 => n1472, B2 => 
                           n13364, C1 => n14549, C2 => n13361, ZN => n10518);
   U5966 : OAI222_X1 port map( A1 => n14801, A2 => n13367, B1 => n1471, B2 => 
                           n13364, C1 => n14543, C2 => n13361, ZN => n10517);
   U5967 : OAI222_X1 port map( A1 => n14795, A2 => n13367, B1 => n1470, B2 => 
                           n13364, C1 => n14537, C2 => n13361, ZN => n10516);
   U5968 : OAI222_X1 port map( A1 => n14789, A2 => n13367, B1 => n1469, B2 => 
                           n13364, C1 => n14531, C2 => n13361, ZN => n10515);
   U5969 : OAI222_X1 port map( A1 => n14783, A2 => n13367, B1 => n1468, B2 => 
                           n13364, C1 => n14525, C2 => n13361, ZN => n10514);
   U5970 : OAI222_X1 port map( A1 => n14777, A2 => n13367, B1 => n1467, B2 => 
                           n13364, C1 => n14519, C2 => n13361, ZN => n10513);
   U5971 : OAI222_X1 port map( A1 => n14771, A2 => n13367, B1 => n1466, B2 => 
                           n13364, C1 => n14513, C2 => n13361, ZN => n10512);
   U5972 : OAI222_X1 port map( A1 => n14765, A2 => n13367, B1 => n1465, B2 => 
                           n13364, C1 => n14714, C2 => n13361, ZN => n10511);
   U5973 : OAI222_X1 port map( A1 => n14759, A2 => n13367, B1 => n1464, B2 => 
                           n13364, C1 => n14702, C2 => n13361, ZN => n10510);
   U5974 : OAI222_X1 port map( A1 => n14753, A2 => n13367, B1 => n1463, B2 => 
                           n13364, C1 => n14693, C2 => n13361, ZN => n10509);
   U5975 : OAI222_X1 port map( A1 => n14885, A2 => n13404, B1 => n1446, B2 => 
                           n13401, C1 => n14627, C2 => n13398, ZN => n10659);
   U5976 : OAI222_X1 port map( A1 => n14879, A2 => n13404, B1 => n1445, B2 => 
                           n13401, C1 => n14621, C2 => n13398, ZN => n10658);
   U5977 : OAI222_X1 port map( A1 => n14873, A2 => n13404, B1 => n1444, B2 => 
                           n13401, C1 => n14615, C2 => n13398, ZN => n10657);
   U5978 : OAI222_X1 port map( A1 => n14867, A2 => n13404, B1 => n1443, B2 => 
                           n13401, C1 => n14609, C2 => n13398, ZN => n10656);
   U5979 : OAI222_X1 port map( A1 => n14861, A2 => n13404, B1 => n1442, B2 => 
                           n13401, C1 => n14603, C2 => n13398, ZN => n10655);
   U5980 : OAI222_X1 port map( A1 => n14855, A2 => n13404, B1 => n1441, B2 => 
                           n13401, C1 => n14597, C2 => n13398, ZN => n10654);
   U5981 : OAI222_X1 port map( A1 => n14849, A2 => n13404, B1 => n1440, B2 => 
                           n13401, C1 => n14591, C2 => n13398, ZN => n10653);
   U5982 : OAI222_X1 port map( A1 => n14843, A2 => n13404, B1 => n1439, B2 => 
                           n13401, C1 => n14585, C2 => n13398, ZN => n10652);
   U5983 : OAI222_X1 port map( A1 => n14837, A2 => n13404, B1 => n1438, B2 => 
                           n13401, C1 => n14579, C2 => n13398, ZN => n10651);
   U5984 : OAI222_X1 port map( A1 => n14831, A2 => n13404, B1 => n1437, B2 => 
                           n13401, C1 => n14573, C2 => n13398, ZN => n10650);
   U5985 : OAI222_X1 port map( A1 => n14825, A2 => n13404, B1 => n1436, B2 => 
                           n13401, C1 => n14567, C2 => n13398, ZN => n10649);
   U5986 : OAI222_X1 port map( A1 => n14819, A2 => n13403, B1 => n1435, B2 => 
                           n13400, C1 => n14561, C2 => n13398, ZN => n10648);
   U5987 : OAI222_X1 port map( A1 => n14813, A2 => n13403, B1 => n1434, B2 => 
                           n13400, C1 => n14555, C2 => n13397, ZN => n10647);
   U5988 : OAI222_X1 port map( A1 => n14807, A2 => n13403, B1 => n1433, B2 => 
                           n13400, C1 => n14549, C2 => n13397, ZN => n10646);
   U5989 : OAI222_X1 port map( A1 => n14801, A2 => n13403, B1 => n1432, B2 => 
                           n13400, C1 => n14543, C2 => n13397, ZN => n10645);
   U5990 : OAI222_X1 port map( A1 => n14795, A2 => n13403, B1 => n1431, B2 => 
                           n13400, C1 => n14537, C2 => n13397, ZN => n10644);
   U5991 : OAI222_X1 port map( A1 => n14789, A2 => n13403, B1 => n1430, B2 => 
                           n13400, C1 => n14531, C2 => n13397, ZN => n10643);
   U5992 : OAI222_X1 port map( A1 => n14783, A2 => n13403, B1 => n1429, B2 => 
                           n13400, C1 => n14525, C2 => n13397, ZN => n10642);
   U5993 : OAI222_X1 port map( A1 => n14777, A2 => n13403, B1 => n1428, B2 => 
                           n13400, C1 => n14519, C2 => n13397, ZN => n10641);
   U5994 : OAI222_X1 port map( A1 => n14771, A2 => n13403, B1 => n1427, B2 => 
                           n13400, C1 => n14513, C2 => n13397, ZN => n10640);
   U5995 : OAI222_X1 port map( A1 => n14765, A2 => n13403, B1 => n1426, B2 => 
                           n13400, C1 => n14714, C2 => n13397, ZN => n10639);
   U5996 : OAI222_X1 port map( A1 => n14759, A2 => n13403, B1 => n1425, B2 => 
                           n13400, C1 => n14702, C2 => n13397, ZN => n10638);
   U5997 : OAI222_X1 port map( A1 => n14753, A2 => n13403, B1 => n1424, B2 => 
                           n13400, C1 => n14693, C2 => n13397, ZN => n10637);
   U5998 : OAI222_X1 port map( A1 => n14885, A2 => n13440, B1 => n1350, B2 => 
                           n13437, C1 => n14626, C2 => n13434, ZN => n10787);
   U5999 : OAI222_X1 port map( A1 => n14879, A2 => n13440, B1 => n1349, B2 => 
                           n13437, C1 => n14620, C2 => n13434, ZN => n10786);
   U6000 : OAI222_X1 port map( A1 => n14873, A2 => n13440, B1 => n1348, B2 => 
                           n13437, C1 => n14614, C2 => n13434, ZN => n10785);
   U6001 : OAI222_X1 port map( A1 => n14867, A2 => n13440, B1 => n1347, B2 => 
                           n13437, C1 => n14608, C2 => n13434, ZN => n10784);
   U6002 : OAI222_X1 port map( A1 => n14861, A2 => n13440, B1 => n1346, B2 => 
                           n13437, C1 => n14602, C2 => n13434, ZN => n10783);
   U6003 : OAI222_X1 port map( A1 => n14855, A2 => n13440, B1 => n1345, B2 => 
                           n13437, C1 => n14596, C2 => n13434, ZN => n10782);
   U6004 : OAI222_X1 port map( A1 => n14849, A2 => n13440, B1 => n1344, B2 => 
                           n13437, C1 => n14590, C2 => n13434, ZN => n10781);
   U6005 : OAI222_X1 port map( A1 => n14843, A2 => n13440, B1 => n1343, B2 => 
                           n13437, C1 => n14584, C2 => n13434, ZN => n10780);
   U6006 : OAI222_X1 port map( A1 => n14837, A2 => n13440, B1 => n1342, B2 => 
                           n13437, C1 => n14578, C2 => n13434, ZN => n10779);
   U6007 : OAI222_X1 port map( A1 => n14831, A2 => n13440, B1 => n1341, B2 => 
                           n13437, C1 => n14572, C2 => n13434, ZN => n10778);
   U6008 : OAI222_X1 port map( A1 => n14825, A2 => n13440, B1 => n1340, B2 => 
                           n13437, C1 => n14566, C2 => n13434, ZN => n10777);
   U6009 : OAI222_X1 port map( A1 => n14819, A2 => n13439, B1 => n1339, B2 => 
                           n13436, C1 => n14560, C2 => n13434, ZN => n10776);
   U6010 : OAI222_X1 port map( A1 => n14813, A2 => n13439, B1 => n1338, B2 => 
                           n13436, C1 => n14554, C2 => n13433, ZN => n10775);
   U6011 : OAI222_X1 port map( A1 => n14807, A2 => n13439, B1 => n1337, B2 => 
                           n13436, C1 => n14548, C2 => n13433, ZN => n10774);
   U6012 : OAI222_X1 port map( A1 => n14801, A2 => n13439, B1 => n1336, B2 => 
                           n13436, C1 => n14542, C2 => n13433, ZN => n10773);
   U6013 : OAI222_X1 port map( A1 => n14795, A2 => n13439, B1 => n1335, B2 => 
                           n13436, C1 => n14536, C2 => n13433, ZN => n10772);
   U6014 : OAI222_X1 port map( A1 => n14789, A2 => n13439, B1 => n1334, B2 => 
                           n13436, C1 => n14530, C2 => n13433, ZN => n10771);
   U6015 : OAI222_X1 port map( A1 => n14783, A2 => n13439, B1 => n1333, B2 => 
                           n13436, C1 => n14524, C2 => n13433, ZN => n10770);
   U6016 : OAI222_X1 port map( A1 => n14777, A2 => n13439, B1 => n1332, B2 => 
                           n13436, C1 => n14518, C2 => n13433, ZN => n10769);
   U6017 : OAI222_X1 port map( A1 => n14771, A2 => n13439, B1 => n1331, B2 => 
                           n13436, C1 => n14512, C2 => n13433, ZN => n10768);
   U6018 : OAI222_X1 port map( A1 => n14765, A2 => n13439, B1 => n1330, B2 => 
                           n13436, C1 => n14713, C2 => n13433, ZN => n10767);
   U6019 : OAI222_X1 port map( A1 => n14759, A2 => n13439, B1 => n1329, B2 => 
                           n13436, C1 => n14701, C2 => n13433, ZN => n10766);
   U6020 : OAI222_X1 port map( A1 => n14753, A2 => n13439, B1 => n1328, B2 => 
                           n13436, C1 => n14693, C2 => n13433, ZN => n10765);
   U6021 : OAI222_X1 port map( A1 => n14885, A2 => n13449, B1 => n1326, B2 => 
                           n13446, C1 => n14626, C2 => n13443, ZN => n10819);
   U6022 : OAI222_X1 port map( A1 => n14879, A2 => n13449, B1 => n1325, B2 => 
                           n13446, C1 => n14620, C2 => n13443, ZN => n10818);
   U6023 : OAI222_X1 port map( A1 => n14873, A2 => n13449, B1 => n1324, B2 => 
                           n13446, C1 => n14614, C2 => n13443, ZN => n10817);
   U6024 : OAI222_X1 port map( A1 => n14867, A2 => n13449, B1 => n1323, B2 => 
                           n13446, C1 => n14608, C2 => n13443, ZN => n10816);
   U6025 : OAI222_X1 port map( A1 => n14861, A2 => n13449, B1 => n1322, B2 => 
                           n13446, C1 => n14602, C2 => n13443, ZN => n10815);
   U6026 : OAI222_X1 port map( A1 => n14855, A2 => n13449, B1 => n1321, B2 => 
                           n13446, C1 => n14596, C2 => n13443, ZN => n10814);
   U6027 : OAI222_X1 port map( A1 => n14849, A2 => n13449, B1 => n1320, B2 => 
                           n13446, C1 => n14590, C2 => n13443, ZN => n10813);
   U6028 : OAI222_X1 port map( A1 => n14843, A2 => n13449, B1 => n1319, B2 => 
                           n13446, C1 => n14584, C2 => n13443, ZN => n10812);
   U6029 : OAI222_X1 port map( A1 => n14837, A2 => n13449, B1 => n1318, B2 => 
                           n13446, C1 => n14578, C2 => n13443, ZN => n10811);
   U6030 : OAI222_X1 port map( A1 => n14831, A2 => n13449, B1 => n1317, B2 => 
                           n13446, C1 => n14572, C2 => n13443, ZN => n10810);
   U6031 : OAI222_X1 port map( A1 => n14825, A2 => n13449, B1 => n1316, B2 => 
                           n13446, C1 => n14566, C2 => n13443, ZN => n10809);
   U6032 : OAI222_X1 port map( A1 => n14819, A2 => n13448, B1 => n1315, B2 => 
                           n13445, C1 => n14560, C2 => n13443, ZN => n10808);
   U6033 : OAI222_X1 port map( A1 => n14813, A2 => n13448, B1 => n1314, B2 => 
                           n13445, C1 => n14554, C2 => n13442, ZN => n10807);
   U6034 : OAI222_X1 port map( A1 => n14807, A2 => n13448, B1 => n1313, B2 => 
                           n13445, C1 => n14548, C2 => n13442, ZN => n10806);
   U6035 : OAI222_X1 port map( A1 => n14801, A2 => n13448, B1 => n1312, B2 => 
                           n13445, C1 => n14542, C2 => n13442, ZN => n10805);
   U6036 : OAI222_X1 port map( A1 => n14795, A2 => n13448, B1 => n1311, B2 => 
                           n13445, C1 => n14536, C2 => n13442, ZN => n10804);
   U6037 : OAI222_X1 port map( A1 => n14789, A2 => n13448, B1 => n1310, B2 => 
                           n13445, C1 => n14530, C2 => n13442, ZN => n10803);
   U6038 : OAI222_X1 port map( A1 => n14783, A2 => n13448, B1 => n1309, B2 => 
                           n13445, C1 => n14524, C2 => n13442, ZN => n10802);
   U6039 : OAI222_X1 port map( A1 => n14777, A2 => n13448, B1 => n1308, B2 => 
                           n13445, C1 => n14518, C2 => n13442, ZN => n10801);
   U6040 : OAI222_X1 port map( A1 => n14770, A2 => n13448, B1 => n1307, B2 => 
                           n13445, C1 => n14512, C2 => n13442, ZN => n10800);
   U6041 : OAI222_X1 port map( A1 => n14765, A2 => n13448, B1 => n1306, B2 => 
                           n13445, C1 => n14713, C2 => n13442, ZN => n10799);
   U6042 : OAI222_X1 port map( A1 => n14759, A2 => n13448, B1 => n1305, B2 => 
                           n13445, C1 => n14701, C2 => n13442, ZN => n10798);
   U6043 : OAI222_X1 port map( A1 => n14753, A2 => n13448, B1 => n1304, B2 => 
                           n13445, C1 => n14694, C2 => n13442, ZN => n10797);
   U6044 : OAI222_X1 port map( A1 => n14818, A2 => n13493, B1 => n786, B2 => 
                           n13490, C1 => n14560, C2 => n13488, ZN => n10968);
   U6045 : OAI222_X1 port map( A1 => n14884, A2 => n13521, B1 => n1191, B2 => 
                           n13518, C1 => n14626, C2 => n13515, ZN => n11075);
   U6046 : OAI222_X1 port map( A1 => n14878, A2 => n13521, B1 => n1190, B2 => 
                           n13518, C1 => n14620, C2 => n13515, ZN => n11074);
   U6047 : OAI222_X1 port map( A1 => n14872, A2 => n13521, B1 => n1189, B2 => 
                           n13518, C1 => n14614, C2 => n13515, ZN => n11073);
   U6048 : OAI222_X1 port map( A1 => n14866, A2 => n13521, B1 => n1188, B2 => 
                           n13518, C1 => n14608, C2 => n13515, ZN => n11072);
   U6049 : OAI222_X1 port map( A1 => n14860, A2 => n13521, B1 => n1187, B2 => 
                           n13518, C1 => n14602, C2 => n13515, ZN => n11071);
   U6050 : OAI222_X1 port map( A1 => n14854, A2 => n13521, B1 => n1186, B2 => 
                           n13518, C1 => n14596, C2 => n13515, ZN => n11070);
   U6051 : OAI222_X1 port map( A1 => n14848, A2 => n13521, B1 => n1185, B2 => 
                           n13518, C1 => n14590, C2 => n13515, ZN => n11069);
   U6052 : OAI222_X1 port map( A1 => n14842, A2 => n13521, B1 => n1184, B2 => 
                           n13518, C1 => n14584, C2 => n13515, ZN => n11068);
   U6053 : OAI222_X1 port map( A1 => n14836, A2 => n13521, B1 => n1183, B2 => 
                           n13518, C1 => n14578, C2 => n13515, ZN => n11067);
   U6054 : OAI222_X1 port map( A1 => n14830, A2 => n13521, B1 => n1182, B2 => 
                           n13518, C1 => n14572, C2 => n13515, ZN => n11066);
   U6055 : OAI222_X1 port map( A1 => n14824, A2 => n13521, B1 => n1181, B2 => 
                           n13518, C1 => n14566, C2 => n13515, ZN => n11065);
   U6056 : OAI222_X1 port map( A1 => n14818, A2 => n13520, B1 => n1180, B2 => 
                           n13517, C1 => n14560, C2 => n13515, ZN => n11064);
   U6057 : OAI222_X1 port map( A1 => n14812, A2 => n13520, B1 => n1179, B2 => 
                           n13517, C1 => n14554, C2 => n13514, ZN => n11063);
   U6058 : OAI222_X1 port map( A1 => n14806, A2 => n13520, B1 => n1178, B2 => 
                           n13517, C1 => n14548, C2 => n13514, ZN => n11062);
   U6059 : OAI222_X1 port map( A1 => n14800, A2 => n13520, B1 => n1177, B2 => 
                           n13517, C1 => n14542, C2 => n13514, ZN => n11061);
   U6060 : OAI222_X1 port map( A1 => n14794, A2 => n13520, B1 => n1176, B2 => 
                           n13517, C1 => n14536, C2 => n13514, ZN => n11060);
   U6061 : OAI222_X1 port map( A1 => n14788, A2 => n13520, B1 => n1175, B2 => 
                           n13517, C1 => n14530, C2 => n13514, ZN => n11059);
   U6062 : OAI222_X1 port map( A1 => n14782, A2 => n13520, B1 => n1174, B2 => 
                           n13517, C1 => n14524, C2 => n13514, ZN => n11058);
   U6063 : OAI222_X1 port map( A1 => n14776, A2 => n13520, B1 => n1173, B2 => 
                           n13517, C1 => n14518, C2 => n13514, ZN => n11057);
   U6064 : OAI222_X1 port map( A1 => n14770, A2 => n13520, B1 => n1172, B2 => 
                           n13517, C1 => n14512, C2 => n13514, ZN => n11056);
   U6065 : OAI222_X1 port map( A1 => n14764, A2 => n13520, B1 => n1171, B2 => 
                           n13517, C1 => n14713, C2 => n13514, ZN => n11055);
   U6066 : OAI222_X1 port map( A1 => n14758, A2 => n13520, B1 => n1170, B2 => 
                           n13517, C1 => n14701, C2 => n13514, ZN => n11054);
   U6067 : OAI222_X1 port map( A1 => n14752, A2 => n13520, B1 => n1169, B2 => 
                           n13517, C1 => n14694, C2 => n13514, ZN => n11053);
   U6068 : OAI222_X1 port map( A1 => n14884, A2 => n13530, B1 => n1167, B2 => 
                           n13527, C1 => n14626, C2 => n13524, ZN => n11107);
   U6069 : OAI222_X1 port map( A1 => n14878, A2 => n13530, B1 => n1166, B2 => 
                           n13527, C1 => n14620, C2 => n13524, ZN => n11106);
   U6070 : OAI222_X1 port map( A1 => n14872, A2 => n13530, B1 => n1165, B2 => 
                           n13527, C1 => n14614, C2 => n13524, ZN => n11105);
   U6071 : OAI222_X1 port map( A1 => n14866, A2 => n13530, B1 => n1164, B2 => 
                           n13527, C1 => n14608, C2 => n13524, ZN => n11104);
   U6072 : OAI222_X1 port map( A1 => n14860, A2 => n13530, B1 => n1163, B2 => 
                           n13527, C1 => n14602, C2 => n13524, ZN => n11103);
   U6073 : OAI222_X1 port map( A1 => n14854, A2 => n13530, B1 => n1162, B2 => 
                           n13527, C1 => n14596, C2 => n13524, ZN => n11102);
   U6074 : OAI222_X1 port map( A1 => n14848, A2 => n13530, B1 => n1161, B2 => 
                           n13527, C1 => n14590, C2 => n13524, ZN => n11101);
   U6075 : OAI222_X1 port map( A1 => n14842, A2 => n13530, B1 => n1160, B2 => 
                           n13527, C1 => n14584, C2 => n13524, ZN => n11100);
   U6076 : OAI222_X1 port map( A1 => n14836, A2 => n13530, B1 => n1159, B2 => 
                           n13527, C1 => n14578, C2 => n13524, ZN => n11099);
   U6077 : OAI222_X1 port map( A1 => n14830, A2 => n13530, B1 => n1158, B2 => 
                           n13527, C1 => n14572, C2 => n13524, ZN => n11098);
   U6078 : OAI222_X1 port map( A1 => n14824, A2 => n13530, B1 => n1157, B2 => 
                           n13527, C1 => n14566, C2 => n13524, ZN => n11097);
   U6079 : OAI222_X1 port map( A1 => n14818, A2 => n13529, B1 => n1156, B2 => 
                           n13526, C1 => n14560, C2 => n13524, ZN => n11096);
   U6080 : OAI222_X1 port map( A1 => n14812, A2 => n13529, B1 => n1155, B2 => 
                           n13526, C1 => n14554, C2 => n13523, ZN => n11095);
   U6081 : OAI222_X1 port map( A1 => n14806, A2 => n13529, B1 => n1154, B2 => 
                           n13526, C1 => n14548, C2 => n13523, ZN => n11094);
   U6082 : OAI222_X1 port map( A1 => n14800, A2 => n13529, B1 => n1153, B2 => 
                           n13526, C1 => n14542, C2 => n13523, ZN => n11093);
   U6083 : OAI222_X1 port map( A1 => n14794, A2 => n13529, B1 => n1152, B2 => 
                           n13526, C1 => n14536, C2 => n13523, ZN => n11092);
   U6084 : OAI222_X1 port map( A1 => n14788, A2 => n13529, B1 => n1151, B2 => 
                           n13526, C1 => n14530, C2 => n13523, ZN => n11091);
   U6085 : OAI222_X1 port map( A1 => n14782, A2 => n13529, B1 => n1150, B2 => 
                           n13526, C1 => n14524, C2 => n13523, ZN => n11090);
   U6086 : OAI222_X1 port map( A1 => n14776, A2 => n13529, B1 => n1149, B2 => 
                           n13526, C1 => n14518, C2 => n13523, ZN => n11089);
   U6087 : OAI222_X1 port map( A1 => n14770, A2 => n13529, B1 => n1148, B2 => 
                           n13526, C1 => n14512, C2 => n13523, ZN => n11088);
   U6088 : OAI222_X1 port map( A1 => n14764, A2 => n13529, B1 => n1147, B2 => 
                           n13526, C1 => n14713, C2 => n13523, ZN => n11087);
   U6089 : OAI222_X1 port map( A1 => n14758, A2 => n13529, B1 => n1146, B2 => 
                           n13526, C1 => n14701, C2 => n13523, ZN => n11086);
   U6090 : OAI222_X1 port map( A1 => n14752, A2 => n13529, B1 => n1145, B2 => 
                           n13526, C1 => n14694, C2 => n13523, ZN => n11085);
   U6091 : OAI222_X1 port map( A1 => n14826, A2 => n13242, B1 => n828, B2 => 
                           n13239, C1 => n14568, C2 => n13236, ZN => n10073);
   U6092 : OAI222_X1 port map( A1 => n14826, A2 => n13251, B1 => n829, B2 => 
                           n13248, C1 => n14568, C2 => n13245, ZN => n10105);
   U6093 : OAI222_X1 port map( A1 => n14892, A2 => n13278, B1 => n1060, B2 => 
                           n13275, C1 => n14634, C2 => n13272, ZN => n10212);
   U6094 : OAI222_X1 port map( A1 => n14886, A2 => n13278, B1 => n1059, B2 => 
                           n13275, C1 => n14628, C2 => n13272, ZN => n10211);
   U6095 : OAI222_X1 port map( A1 => n14880, A2 => n13278, B1 => n1058, B2 => 
                           n13275, C1 => n14622, C2 => n13272, ZN => n10210);
   U6096 : OAI222_X1 port map( A1 => n14874, A2 => n13278, B1 => n1057, B2 => 
                           n13275, C1 => n14616, C2 => n13272, ZN => n10209);
   U6097 : OAI222_X1 port map( A1 => n14868, A2 => n13278, B1 => n1056, B2 => 
                           n13275, C1 => n14610, C2 => n13272, ZN => n10208);
   U6098 : OAI222_X1 port map( A1 => n14862, A2 => n13278, B1 => n1055, B2 => 
                           n13275, C1 => n14604, C2 => n13272, ZN => n10207);
   U6099 : OAI222_X1 port map( A1 => n14856, A2 => n13278, B1 => n1054, B2 => 
                           n13275, C1 => n14598, C2 => n13272, ZN => n10206);
   U6100 : OAI222_X1 port map( A1 => n14850, A2 => n13278, B1 => n1053, B2 => 
                           n13275, C1 => n14592, C2 => n13272, ZN => n10205);
   U6101 : OAI222_X1 port map( A1 => n14844, A2 => n13278, B1 => n1052, B2 => 
                           n13275, C1 => n14586, C2 => n13272, ZN => n10204);
   U6102 : OAI222_X1 port map( A1 => n14838, A2 => n13278, B1 => n1051, B2 => 
                           n13275, C1 => n14580, C2 => n13272, ZN => n10203);
   U6103 : OAI222_X1 port map( A1 => n14832, A2 => n13278, B1 => n1050, B2 => 
                           n13275, C1 => n14574, C2 => n13272, ZN => n10202);
   U6104 : OAI222_X1 port map( A1 => n14826, A2 => n13278, B1 => n1049, B2 => 
                           n13275, C1 => n14568, C2 => n13272, ZN => n10201);
   U6105 : OAI222_X1 port map( A1 => n14820, A2 => n13277, B1 => n1048, B2 => 
                           n13274, C1 => n14562, C2 => n13272, ZN => n10200);
   U6106 : OAI222_X1 port map( A1 => n14814, A2 => n13277, B1 => n1047, B2 => 
                           n13274, C1 => n14556, C2 => n13271, ZN => n10199);
   U6107 : OAI222_X1 port map( A1 => n14808, A2 => n13277, B1 => n1046, B2 => 
                           n13274, C1 => n14550, C2 => n13271, ZN => n10198);
   U6108 : OAI222_X1 port map( A1 => n14802, A2 => n13277, B1 => n1045, B2 => 
                           n13274, C1 => n14544, C2 => n13271, ZN => n10197);
   U6109 : OAI222_X1 port map( A1 => n14796, A2 => n13277, B1 => n1044, B2 => 
                           n13274, C1 => n14538, C2 => n13271, ZN => n10196);
   U6110 : OAI222_X1 port map( A1 => n14790, A2 => n13277, B1 => n1043, B2 => 
                           n13274, C1 => n14532, C2 => n13271, ZN => n10195);
   U6111 : OAI222_X1 port map( A1 => n14784, A2 => n13277, B1 => n1042, B2 => 
                           n13274, C1 => n14526, C2 => n13271, ZN => n10194);
   U6112 : OAI222_X1 port map( A1 => n14778, A2 => n13277, B1 => n1041, B2 => 
                           n13274, C1 => n14520, C2 => n13271, ZN => n10193);
   U6113 : OAI222_X1 port map( A1 => n14772, A2 => n13277, B1 => n1040, B2 => 
                           n13274, C1 => n14514, C2 => n13271, ZN => n10192);
   U6114 : OAI222_X1 port map( A1 => n14766, A2 => n13277, B1 => n1039, B2 => 
                           n13274, C1 => n14715, C2 => n13271, ZN => n10191);
   U6115 : OAI222_X1 port map( A1 => n14760, A2 => n13277, B1 => n1038, B2 => 
                           n13274, C1 => n14703, C2 => n13271, ZN => n10190);
   U6116 : OAI222_X1 port map( A1 => n14754, A2 => n13277, B1 => n1037, B2 => 
                           n13274, C1 => n14692, C2 => n13271, ZN => n10189);
   U6117 : OAI222_X1 port map( A1 => n14882, A2 => n14343, B1 => n14339, B2 => 
                           n1035, C1 => n14624, C2 => n14337, ZN => n9379);
   U6118 : OAI222_X1 port map( A1 => n14876, A2 => n14343, B1 => n14339, B2 => 
                           n1034, C1 => n14618, C2 => n14337, ZN => n9378);
   U6119 : OAI222_X1 port map( A1 => n14870, A2 => n14343, B1 => n14339, B2 => 
                           n1033, C1 => n14612, C2 => n14337, ZN => n9377);
   U6120 : OAI222_X1 port map( A1 => n14864, A2 => n14343, B1 => n14340, B2 => 
                           n1032, C1 => n14606, C2 => n14337, ZN => n9376);
   U6121 : OAI222_X1 port map( A1 => n14858, A2 => n14343, B1 => n14340, B2 => 
                           n1031, C1 => n14600, C2 => n14337, ZN => n9375);
   U6122 : OAI222_X1 port map( A1 => n14852, A2 => n14343, B1 => n14340, B2 => 
                           n1030, C1 => n14594, C2 => n14337, ZN => n9374);
   U6123 : OAI222_X1 port map( A1 => n14846, A2 => n14343, B1 => n14340, B2 => 
                           n1029, C1 => n14588, C2 => n14337, ZN => n9373);
   U6124 : OAI222_X1 port map( A1 => n14840, A2 => n14343, B1 => n14340, B2 => 
                           n1028, C1 => n14582, C2 => n14337, ZN => n9372);
   U6125 : OAI222_X1 port map( A1 => n14834, A2 => n14343, B1 => n14340, B2 => 
                           n1027, C1 => n14576, C2 => n14337, ZN => n9371);
   U6126 : OAI222_X1 port map( A1 => n14828, A2 => n14343, B1 => n14340, B2 => 
                           n1026, C1 => n14570, C2 => n14337, ZN => n9370);
   U6127 : OAI222_X1 port map( A1 => n14822, A2 => n14343, B1 => n806, B2 => 
                           n14341, C1 => n14564, C2 => n14337, ZN => n9369);
   U6128 : OAI222_X1 port map( A1 => n14816, A2 => n14342, B1 => n14340, B2 => 
                           n1024, C1 => n14558, C2 => n14337, ZN => n9368);
   U6129 : OAI222_X1 port map( A1 => n14810, A2 => n14342, B1 => n14340, B2 => 
                           n1023, C1 => n14552, C2 => n14336, ZN => n9367);
   U6130 : OAI222_X1 port map( A1 => n14804, A2 => n14342, B1 => n14340, B2 => 
                           n1022, C1 => n14546, C2 => n14336, ZN => n9366);
   U6131 : OAI222_X1 port map( A1 => n14798, A2 => n14342, B1 => n14340, B2 => 
                           n1021, C1 => n14540, C2 => n14336, ZN => n9365);
   U6132 : OAI222_X1 port map( A1 => n14792, A2 => n14342, B1 => n14341, B2 => 
                           n1020, C1 => n14534, C2 => n14336, ZN => n9364);
   U6133 : OAI222_X1 port map( A1 => n14786, A2 => n14342, B1 => n14341, B2 => 
                           n1019, C1 => n14528, C2 => n14336, ZN => n9363);
   U6134 : OAI222_X1 port map( A1 => n14780, A2 => n14342, B1 => n14341, B2 => 
                           n1018, C1 => n14522, C2 => n14336, ZN => n9362);
   U6135 : OAI222_X1 port map( A1 => n14774, A2 => n14342, B1 => n14341, B2 => 
                           n1017, C1 => n14516, C2 => n14336, ZN => n9361);
   U6136 : OAI222_X1 port map( A1 => n14768, A2 => n14342, B1 => n14341, B2 => 
                           n1016, C1 => n14510, C2 => n14336, ZN => n9360);
   U6137 : OAI222_X1 port map( A1 => n14762, A2 => n14342, B1 => n14341, B2 => 
                           n1015, C1 => n14711, C2 => n14336, ZN => n9359);
   U6138 : OAI222_X1 port map( A1 => n14756, A2 => n14342, B1 => n14341, B2 => 
                           n1014, C1 => n14699, C2 => n14336, ZN => n9358);
   U6139 : OAI222_X1 port map( A1 => n14750, A2 => n14342, B1 => n14339, B2 => 
                           n1013, C1 => n14696, C2 => n14336, ZN => n9357);
   U6140 : OAI222_X1 port map( A1 => n14822, A2 => n14352, B1 => n807, B2 => 
                           n14350, C1 => n14565, C2 => n14346, ZN => n9401);
   U6141 : OAI222_X1 port map( A1 => n14816, A2 => n14351, B1 => n743, B2 => 
                           n14350, C1 => n14559, C2 => n14346, ZN => n9400);
   U6142 : OAI222_X1 port map( A1 => n14822, A2 => n14381, B1 => n810, B2 => 
                           n14379, C1 => n14564, C2 => n14375, ZN => n9497);
   U6143 : OAI222_X1 port map( A1 => n14817, A2 => n13592, B1 => n795, B2 => 
                           n13589, C1 => n14559, C2 => n13587, ZN => n11320);
   U6144 : OAI222_X1 port map( A1 => n14811, A2 => n13592, B1 => n731, B2 => 
                           n13589, C1 => n14553, C2 => n13586, ZN => n11319);
   U6145 : OAI222_X1 port map( A1 => n14823, A2 => n14294, B1 => n801, B2 => 
                           n14292, C1 => n14564, C2 => n14288, ZN => n9191);
   U6146 : OAI222_X1 port map( A1 => n14823, A2 => n14305, B1 => n802, B2 => 
                           n14303, C1 => n14564, C2 => n14299, ZN => n9241);
   U6147 : OAI222_X1 port map( A1 => n14882, A2 => n14334, B1 => n14330, B2 => 
                           n554, C1 => n14624, C2 => n14328, ZN => n9347);
   U6148 : OAI222_X1 port map( A1 => n14876, A2 => n14334, B1 => n14330, B2 => 
                           n553, C1 => n14618, C2 => n14328, ZN => n9346);
   U6149 : OAI222_X1 port map( A1 => n14870, A2 => n14334, B1 => n14330, B2 => 
                           n552, C1 => n14612, C2 => n14328, ZN => n9345);
   U6150 : OAI222_X1 port map( A1 => n14864, A2 => n14334, B1 => n14331, B2 => 
                           n551, C1 => n14606, C2 => n14328, ZN => n9344);
   U6151 : OAI222_X1 port map( A1 => n14858, A2 => n14334, B1 => n14331, B2 => 
                           n550, C1 => n14600, C2 => n14328, ZN => n9343);
   U6152 : OAI222_X1 port map( A1 => n14852, A2 => n14334, B1 => n14331, B2 => 
                           n549, C1 => n14594, C2 => n14328, ZN => n9342);
   U6153 : OAI222_X1 port map( A1 => n14846, A2 => n14334, B1 => n14331, B2 => 
                           n548, C1 => n14588, C2 => n14328, ZN => n9341);
   U6154 : OAI222_X1 port map( A1 => n14840, A2 => n14334, B1 => n14331, B2 => 
                           n547, C1 => n14582, C2 => n14328, ZN => n9340);
   U6155 : OAI222_X1 port map( A1 => n14834, A2 => n14334, B1 => n14331, B2 => 
                           n546, C1 => n14576, C2 => n14328, ZN => n9339);
   U6156 : OAI222_X1 port map( A1 => n14828, A2 => n14334, B1 => n14331, B2 => 
                           n545, C1 => n14570, C2 => n14328, ZN => n9338);
   U6157 : OAI222_X1 port map( A1 => n14822, A2 => n14334, B1 => n805, B2 => 
                           n14332, C1 => n14564, C2 => n14328, ZN => n9337);
   U6158 : OAI222_X1 port map( A1 => n14816, A2 => n14333, B1 => n14331, B2 => 
                           n543, C1 => n14558, C2 => n14328, ZN => n9336);
   U6159 : OAI222_X1 port map( A1 => n14810, A2 => n14333, B1 => n14331, B2 => 
                           n542, C1 => n14552, C2 => n14327, ZN => n9335);
   U6160 : OAI222_X1 port map( A1 => n14804, A2 => n14333, B1 => n14331, B2 => 
                           n541, C1 => n14546, C2 => n14327, ZN => n9334);
   U6161 : OAI222_X1 port map( A1 => n14798, A2 => n14333, B1 => n14331, B2 => 
                           n540, C1 => n14540, C2 => n14327, ZN => n9333);
   U6162 : OAI222_X1 port map( A1 => n14792, A2 => n14333, B1 => n14332, B2 => 
                           n539, C1 => n14534, C2 => n14327, ZN => n9332);
   U6163 : OAI222_X1 port map( A1 => n14786, A2 => n14333, B1 => n14332, B2 => 
                           n538, C1 => n14528, C2 => n14327, ZN => n9331);
   U6164 : OAI222_X1 port map( A1 => n14780, A2 => n14333, B1 => n14332, B2 => 
                           n537, C1 => n14522, C2 => n14327, ZN => n9330);
   U6165 : OAI222_X1 port map( A1 => n14774, A2 => n14333, B1 => n14332, B2 => 
                           n536, C1 => n14516, C2 => n14327, ZN => n9329);
   U6166 : OAI222_X1 port map( A1 => n14768, A2 => n14333, B1 => n14332, B2 => 
                           n535, C1 => n14510, C2 => n14327, ZN => n9328);
   U6167 : OAI222_X1 port map( A1 => n14762, A2 => n14333, B1 => n14332, B2 => 
                           n534, C1 => n14711, C2 => n14327, ZN => n9327);
   U6168 : OAI222_X1 port map( A1 => n14756, A2 => n14333, B1 => n14332, B2 => 
                           n533, C1 => n14699, C2 => n14327, ZN => n9326);
   U6169 : OAI222_X1 port map( A1 => n14750, A2 => n14333, B1 => n14330, B2 => 
                           n532, C1 => n14696, C2 => n14327, ZN => n9325);
   U6170 : OAI222_X1 port map( A1 => n14822, A2 => n14390, B1 => n811, B2 => 
                           n14388, C1 => n14564, C2 => n14384, ZN => n9529);
   U6171 : OAI222_X1 port map( A1 => n14882, A2 => n14417, B1 => n14413, B2 => 
                           n458, C1 => n14623, C2 => n14411, ZN => n9635);
   U6172 : OAI222_X1 port map( A1 => n14876, A2 => n14417, B1 => n14413, B2 => 
                           n457, C1 => n14617, C2 => n14411, ZN => n9634);
   U6173 : OAI222_X1 port map( A1 => n14870, A2 => n14417, B1 => n14413, B2 => 
                           n456, C1 => n14611, C2 => n14411, ZN => n9633);
   U6174 : OAI222_X1 port map( A1 => n14864, A2 => n14417, B1 => n14414, B2 => 
                           n455, C1 => n14605, C2 => n14411, ZN => n9632);
   U6175 : OAI222_X1 port map( A1 => n14858, A2 => n14417, B1 => n14414, B2 => 
                           n454, C1 => n14599, C2 => n14411, ZN => n9631);
   U6176 : OAI222_X1 port map( A1 => n14852, A2 => n14417, B1 => n14414, B2 => 
                           n453, C1 => n14593, C2 => n14411, ZN => n9630);
   U6177 : OAI222_X1 port map( A1 => n14846, A2 => n14417, B1 => n14414, B2 => 
                           n452, C1 => n14587, C2 => n14411, ZN => n9629);
   U6178 : OAI222_X1 port map( A1 => n14840, A2 => n14417, B1 => n14414, B2 => 
                           n451, C1 => n14581, C2 => n14411, ZN => n9628);
   U6179 : OAI222_X1 port map( A1 => n14834, A2 => n14417, B1 => n14414, B2 => 
                           n450, C1 => n14575, C2 => n14411, ZN => n9627);
   U6180 : OAI222_X1 port map( A1 => n14828, A2 => n14417, B1 => n14414, B2 => 
                           n449, C1 => n14569, C2 => n14411, ZN => n9626);
   U6181 : OAI222_X1 port map( A1 => n14822, A2 => n14417, B1 => n814, B2 => 
                           n14415, C1 => n14563, C2 => n14411, ZN => n9625);
   U6182 : OAI222_X1 port map( A1 => n14816, A2 => n14416, B1 => n14414, B2 => 
                           n447, C1 => n14557, C2 => n14411, ZN => n9624);
   U6183 : OAI222_X1 port map( A1 => n14810, A2 => n14416, B1 => n14414, B2 => 
                           n446, C1 => n14551, C2 => n14410, ZN => n9623);
   U6184 : OAI222_X1 port map( A1 => n14804, A2 => n14416, B1 => n14414, B2 => 
                           n445, C1 => n14545, C2 => n14410, ZN => n9622);
   U6185 : OAI222_X1 port map( A1 => n14798, A2 => n14416, B1 => n14414, B2 => 
                           n444, C1 => n14539, C2 => n14410, ZN => n9621);
   U6186 : OAI222_X1 port map( A1 => n14792, A2 => n14416, B1 => n14415, B2 => 
                           n443, C1 => n14533, C2 => n14410, ZN => n9620);
   U6187 : OAI222_X1 port map( A1 => n14786, A2 => n14416, B1 => n14415, B2 => 
                           n442, C1 => n14527, C2 => n14410, ZN => n9619);
   U6188 : OAI222_X1 port map( A1 => n14780, A2 => n14416, B1 => n14415, B2 => 
                           n441, C1 => n14521, C2 => n14410, ZN => n9618);
   U6189 : OAI222_X1 port map( A1 => n14774, A2 => n14416, B1 => n14415, B2 => 
                           n440, C1 => n14515, C2 => n14410, ZN => n9617);
   U6190 : OAI222_X1 port map( A1 => n14768, A2 => n14416, B1 => n14415, B2 => 
                           n439, C1 => n14509, C2 => n14410, ZN => n9616);
   U6191 : OAI222_X1 port map( A1 => n14762, A2 => n14416, B1 => n14415, B2 => 
                           n438, C1 => n14710, C2 => n14410, ZN => n9615);
   U6192 : OAI222_X1 port map( A1 => n14756, A2 => n14416, B1 => n14415, B2 => 
                           n437, C1 => n14698, C2 => n14410, ZN => n9614);
   U6193 : OAI222_X1 port map( A1 => n14750, A2 => n14416, B1 => n14413, B2 => 
                           n436, C1 => n14696, C2 => n14410, ZN => n9613);
   U6194 : OAI222_X1 port map( A1 => n14882, A2 => n14426, B1 => n14422, B2 => 
                           n434, C1 => n14623, C2 => n14420, ZN => n9667);
   U6195 : OAI222_X1 port map( A1 => n14876, A2 => n14426, B1 => n14422, B2 => 
                           n433, C1 => n14617, C2 => n14420, ZN => n9666);
   U6196 : OAI222_X1 port map( A1 => n14870, A2 => n14426, B1 => n14422, B2 => 
                           n432, C1 => n14611, C2 => n14420, ZN => n9665);
   U6197 : OAI222_X1 port map( A1 => n14864, A2 => n14426, B1 => n14423, B2 => 
                           n431, C1 => n14605, C2 => n14420, ZN => n9664);
   U6198 : OAI222_X1 port map( A1 => n14858, A2 => n14426, B1 => n14423, B2 => 
                           n430, C1 => n14599, C2 => n14420, ZN => n9663);
   U6199 : OAI222_X1 port map( A1 => n14852, A2 => n14426, B1 => n14423, B2 => 
                           n429, C1 => n14593, C2 => n14420, ZN => n9662);
   U6200 : OAI222_X1 port map( A1 => n14846, A2 => n14426, B1 => n14423, B2 => 
                           n428, C1 => n14587, C2 => n14420, ZN => n9661);
   U6201 : OAI222_X1 port map( A1 => n14840, A2 => n14426, B1 => n14423, B2 => 
                           n427, C1 => n14581, C2 => n14420, ZN => n9660);
   U6202 : OAI222_X1 port map( A1 => n14834, A2 => n14426, B1 => n14423, B2 => 
                           n426, C1 => n14575, C2 => n14420, ZN => n9659);
   U6203 : OAI222_X1 port map( A1 => n14828, A2 => n14426, B1 => n14423, B2 => 
                           n425, C1 => n14569, C2 => n14420, ZN => n9658);
   U6204 : OAI222_X1 port map( A1 => n14822, A2 => n14426, B1 => n815, B2 => 
                           n14424, C1 => n14563, C2 => n14420, ZN => n9657);
   U6205 : OAI222_X1 port map( A1 => n14816, A2 => n14425, B1 => n14423, B2 => 
                           n423, C1 => n14557, C2 => n14420, ZN => n9656);
   U6206 : OAI222_X1 port map( A1 => n14810, A2 => n14425, B1 => n14423, B2 => 
                           n422, C1 => n14551, C2 => n14419, ZN => n9655);
   U6207 : OAI222_X1 port map( A1 => n14804, A2 => n14425, B1 => n14423, B2 => 
                           n421, C1 => n14545, C2 => n14419, ZN => n9654);
   U6208 : OAI222_X1 port map( A1 => n14798, A2 => n14425, B1 => n14423, B2 => 
                           n420, C1 => n14539, C2 => n14419, ZN => n9653);
   U6209 : OAI222_X1 port map( A1 => n14792, A2 => n14425, B1 => n14424, B2 => 
                           n419, C1 => n14533, C2 => n14419, ZN => n9652);
   U6210 : OAI222_X1 port map( A1 => n14786, A2 => n14425, B1 => n14424, B2 => 
                           n418, C1 => n14527, C2 => n14419, ZN => n9651);
   U6211 : OAI222_X1 port map( A1 => n14780, A2 => n14425, B1 => n14424, B2 => 
                           n417, C1 => n14521, C2 => n14419, ZN => n9650);
   U6212 : OAI222_X1 port map( A1 => n14774, A2 => n14425, B1 => n14424, B2 => 
                           n416, C1 => n14515, C2 => n14419, ZN => n9649);
   U6213 : OAI222_X1 port map( A1 => n14767, A2 => n14425, B1 => n14424, B2 => 
                           n415, C1 => n14509, C2 => n14419, ZN => n9648);
   U6214 : OAI222_X1 port map( A1 => n14762, A2 => n14425, B1 => n14424, B2 => 
                           n414, C1 => n14710, C2 => n14419, ZN => n9647);
   U6215 : OAI222_X1 port map( A1 => n14756, A2 => n14425, B1 => n14424, B2 => 
                           n413, C1 => n14698, C2 => n14419, ZN => n9646);
   U6216 : OAI222_X1 port map( A1 => n14750, A2 => n14425, B1 => n14422, B2 => 
                           n412, C1 => n14697, C2 => n14419, ZN => n9645);
   U6217 : OAI222_X1 port map( A1 => n2620, A2 => n14087, B1 => n4064, B2 => 
                           n14084, C1 => n14076, C2 => n2151, ZN => n9165);
   U6218 : NOR4_X1 port map( A1 => n4065, A2 => n4066, A3 => n4067, A4 => n4068
                           , ZN => n4064);
   U6219 : NAND4_X1 port map( A1 => n4095, A2 => n4096, A3 => n4097, A4 => 
                           n4098, ZN => n4065);
   U6220 : NAND4_X1 port map( A1 => n4085, A2 => n4086, A3 => n4087, A4 => 
                           n4088, ZN => n4066);
   U6221 : OAI222_X1 port map( A1 => n2619, A2 => n14087, B1 => n4103, B2 => 
                           n14084, C1 => n14076, C2 => n2152, ZN => n9164);
   U6222 : NOR4_X1 port map( A1 => n4104, A2 => n4105, A3 => n4106, A4 => n4107
                           , ZN => n4103);
   U6223 : NAND4_X1 port map( A1 => n4132, A2 => n4133, A3 => n4134, A4 => 
                           n4135, ZN => n4104);
   U6224 : NAND4_X1 port map( A1 => n4124, A2 => n4125, A3 => n4126, A4 => 
                           n4127, ZN => n4105);
   U6225 : OAI222_X1 port map( A1 => n2619, A2 => n13867, B1 => n5424, B2 => 
                           n13864, C1 => n13856, C2 => n2184, ZN => n9131);
   U6226 : NOR4_X1 port map( A1 => n5425, A2 => n5426, A3 => n5427, A4 => n5428
                           , ZN => n5424);
   U6227 : NAND4_X1 port map( A1 => n5453, A2 => n5454, A3 => n5455, A4 => 
                           n5456, ZN => n5425);
   U6228 : NAND4_X1 port map( A1 => n5445, A2 => n5446, A3 => n5447, A4 => 
                           n5448, ZN => n5426);
   U6229 : OAI222_X1 port map( A1 => n2618, A2 => n14087, B1 => n4140, B2 => 
                           n14084, C1 => n14076, C2 => n2153, ZN => n9163);
   U6230 : NOR4_X1 port map( A1 => n4141, A2 => n4142, A3 => n4143, A4 => n4144
                           , ZN => n4140);
   U6231 : NAND4_X1 port map( A1 => n4169, A2 => n4170, A3 => n4171, A4 => 
                           n4172, ZN => n4141);
   U6232 : NAND4_X1 port map( A1 => n4161, A2 => n4162, A3 => n4163, A4 => 
                           n4164, ZN => n4142);
   U6233 : OAI222_X1 port map( A1 => n2617, A2 => n14087, B1 => n4177, B2 => 
                           n14084, C1 => n14076, C2 => n2154, ZN => n9162);
   U6234 : NOR4_X1 port map( A1 => n4178, A2 => n4179, A3 => n4180, A4 => n4181
                           , ZN => n4177);
   U6235 : NAND4_X1 port map( A1 => n4206, A2 => n4207, A3 => n4208, A4 => 
                           n4209, ZN => n4178);
   U6236 : NAND4_X1 port map( A1 => n4198, A2 => n4199, A3 => n4200, A4 => 
                           n4201, ZN => n4179);
   U6237 : OAI222_X1 port map( A1 => n2616, A2 => n14087, B1 => n4214, B2 => 
                           n14084, C1 => n14076, C2 => n2155, ZN => n9161);
   U6238 : NOR4_X1 port map( A1 => n4215, A2 => n4216, A3 => n4217, A4 => n4218
                           , ZN => n4214);
   U6239 : NAND4_X1 port map( A1 => n4243, A2 => n4244, A3 => n4245, A4 => 
                           n4246, ZN => n4215);
   U6240 : NAND4_X1 port map( A1 => n4235, A2 => n4236, A3 => n4237, A4 => 
                           n4238, ZN => n4216);
   U6241 : OAI222_X1 port map( A1 => n2614, A2 => n13866, B1 => n5609, B2 => 
                           n13864, C1 => n13856, C2 => n2189, ZN => n9126);
   U6242 : NOR4_X1 port map( A1 => n5610, A2 => n5611, A3 => n5612, A4 => n5613
                           , ZN => n5609);
   U6243 : NAND4_X1 port map( A1 => n5638, A2 => n5639, A3 => n5640, A4 => 
                           n5641, ZN => n5610);
   U6244 : NAND4_X1 port map( A1 => n5630, A2 => n5631, A3 => n5632, A4 => 
                           n5633, ZN => n5611);
   U6245 : OAI222_X1 port map( A1 => n2613, A2 => n14086, B1 => n4325, B2 => 
                           n14083, C1 => n14076, C2 => n2158, ZN => n9158);
   U6246 : NOR4_X1 port map( A1 => n4326, A2 => n4327, A3 => n4328, A4 => n4329
                           , ZN => n4325);
   U6247 : NAND4_X1 port map( A1 => n4354, A2 => n4355, A3 => n4356, A4 => 
                           n4357, ZN => n4326);
   U6248 : NAND4_X1 port map( A1 => n4346, A2 => n4347, A3 => n4348, A4 => 
                           n4349, ZN => n4327);
   U6249 : OAI222_X1 port map( A1 => n2613, A2 => n13866, B1 => n5646, B2 => 
                           n13863, C1 => n13856, C2 => n2190, ZN => n9125);
   U6250 : NOR4_X1 port map( A1 => n5647, A2 => n5648, A3 => n5649, A4 => n5650
                           , ZN => n5646);
   U6251 : NAND4_X1 port map( A1 => n5675, A2 => n5676, A3 => n5677, A4 => 
                           n5678, ZN => n5647);
   U6252 : NAND4_X1 port map( A1 => n5667, A2 => n5668, A3 => n5669, A4 => 
                           n5670, ZN => n5648);
   U6253 : OAI222_X1 port map( A1 => n2612, A2 => n14086, B1 => n4362, B2 => 
                           n14083, C1 => n14076, C2 => n2159, ZN => n9157);
   U6254 : NOR4_X1 port map( A1 => n4363, A2 => n4364, A3 => n4365, A4 => n4366
                           , ZN => n4362);
   U6255 : NAND4_X1 port map( A1 => n4391, A2 => n4392, A3 => n4393, A4 => 
                           n4394, ZN => n4363);
   U6256 : NAND4_X1 port map( A1 => n4383, A2 => n4384, A3 => n4385, A4 => 
                           n4386, ZN => n4364);
   U6257 : OAI222_X1 port map( A1 => n2612, A2 => n13866, B1 => n5683, B2 => 
                           n13863, C1 => n13856, C2 => n2191, ZN => n9124);
   U6258 : NOR4_X1 port map( A1 => n5684, A2 => n5685, A3 => n5686, A4 => n5687
                           , ZN => n5683);
   U6259 : NAND4_X1 port map( A1 => n5712, A2 => n5713, A3 => n5714, A4 => 
                           n5715, ZN => n5684);
   U6260 : NAND4_X1 port map( A1 => n5704, A2 => n5705, A3 => n5706, A4 => 
                           n5707, ZN => n5685);
   U6261 : OAI222_X1 port map( A1 => n2611, A2 => n14086, B1 => n4399, B2 => 
                           n14083, C1 => n14076, C2 => n2160, ZN => n9156);
   U6262 : NOR4_X1 port map( A1 => n4400, A2 => n4401, A3 => n4402, A4 => n4403
                           , ZN => n4399);
   U6263 : NAND4_X1 port map( A1 => n4428, A2 => n4429, A3 => n4430, A4 => 
                           n4431, ZN => n4400);
   U6264 : NAND4_X1 port map( A1 => n4420, A2 => n4421, A3 => n4422, A4 => 
                           n4423, ZN => n4401);
   U6265 : OAI222_X1 port map( A1 => n2611, A2 => n13866, B1 => n5720, B2 => 
                           n13863, C1 => n13856, C2 => n2192, ZN => n9123);
   U6266 : NOR4_X1 port map( A1 => n5721, A2 => n5722, A3 => n5723, A4 => n5724
                           , ZN => n5720);
   U6267 : NAND4_X1 port map( A1 => n5749, A2 => n5750, A3 => n5751, A4 => 
                           n5752, ZN => n5721);
   U6268 : NAND4_X1 port map( A1 => n5741, A2 => n5742, A3 => n5743, A4 => 
                           n5744, ZN => n5722);
   U6269 : OAI222_X1 port map( A1 => n2610, A2 => n14086, B1 => n4436, B2 => 
                           n14083, C1 => n14076, C2 => n2161, ZN => n9155);
   U6270 : NOR4_X1 port map( A1 => n4437, A2 => n4438, A3 => n4439, A4 => n4440
                           , ZN => n4436);
   U6271 : NAND4_X1 port map( A1 => n4465, A2 => n4466, A3 => n4467, A4 => 
                           n4468, ZN => n4437);
   U6272 : NAND4_X1 port map( A1 => n4457, A2 => n4458, A3 => n4459, A4 => 
                           n4460, ZN => n4438);
   U6273 : OAI222_X1 port map( A1 => n2610, A2 => n13866, B1 => n5757, B2 => 
                           n13863, C1 => n13856, C2 => n2193, ZN => n9122);
   U6274 : NOR4_X1 port map( A1 => n5758, A2 => n5759, A3 => n5760, A4 => n5761
                           , ZN => n5757);
   U6275 : NAND4_X1 port map( A1 => n5786, A2 => n5787, A3 => n5788, A4 => 
                           n5789, ZN => n5758);
   U6276 : NAND4_X1 port map( A1 => n5778, A2 => n5779, A3 => n5780, A4 => 
                           n5781, ZN => n5759);
   U6277 : OAI222_X1 port map( A1 => n2609, A2 => n14086, B1 => n4473, B2 => 
                           n14083, C1 => n14077, C2 => n2162, ZN => n9154);
   U6278 : NOR4_X1 port map( A1 => n4474, A2 => n4475, A3 => n4476, A4 => n4477
                           , ZN => n4473);
   U6279 : NAND4_X1 port map( A1 => n4502, A2 => n4503, A3 => n4504, A4 => 
                           n4505, ZN => n4474);
   U6280 : NAND4_X1 port map( A1 => n4494, A2 => n4495, A3 => n4496, A4 => 
                           n4497, ZN => n4475);
   U6281 : OAI222_X1 port map( A1 => n2609, A2 => n13866, B1 => n5794, B2 => 
                           n13863, C1 => n13857, C2 => n2194, ZN => n9121);
   U6282 : NOR4_X1 port map( A1 => n5795, A2 => n5796, A3 => n5797, A4 => n5798
                           , ZN => n5794);
   U6283 : NAND4_X1 port map( A1 => n5823, A2 => n5824, A3 => n5825, A4 => 
                           n5826, ZN => n5795);
   U6284 : NAND4_X1 port map( A1 => n5815, A2 => n5816, A3 => n5817, A4 => 
                           n5818, ZN => n5796);
   U6285 : OAI222_X1 port map( A1 => n2608, A2 => n14086, B1 => n4510, B2 => 
                           n14083, C1 => n14077, C2 => n2163, ZN => n9153);
   U6286 : NOR4_X1 port map( A1 => n4511, A2 => n4512, A3 => n4513, A4 => n4514
                           , ZN => n4510);
   U6287 : NAND4_X1 port map( A1 => n4539, A2 => n4540, A3 => n4541, A4 => 
                           n4542, ZN => n4511);
   U6288 : NAND4_X1 port map( A1 => n4531, A2 => n4532, A3 => n4533, A4 => 
                           n4534, ZN => n4512);
   U6289 : OAI222_X1 port map( A1 => n2608, A2 => n13866, B1 => n5831, B2 => 
                           n13863, C1 => n13857, C2 => n2195, ZN => n9120);
   U6290 : NOR4_X1 port map( A1 => n5832, A2 => n5833, A3 => n5834, A4 => n5835
                           , ZN => n5831);
   U6291 : NAND4_X1 port map( A1 => n5860, A2 => n5861, A3 => n5862, A4 => 
                           n5863, ZN => n5832);
   U6292 : NAND4_X1 port map( A1 => n5852, A2 => n5853, A3 => n5854, A4 => 
                           n5855, ZN => n5833);
   U6293 : OAI222_X1 port map( A1 => n2607, A2 => n14086, B1 => n4547, B2 => 
                           n14083, C1 => n14077, C2 => n2164, ZN => n9152);
   U6294 : NOR4_X1 port map( A1 => n4548, A2 => n4549, A3 => n4550, A4 => n4551
                           , ZN => n4547);
   U6295 : NAND4_X1 port map( A1 => n4576, A2 => n4577, A3 => n4578, A4 => 
                           n4579, ZN => n4548);
   U6296 : NAND4_X1 port map( A1 => n4568, A2 => n4569, A3 => n4570, A4 => 
                           n4571, ZN => n4549);
   U6297 : OAI222_X1 port map( A1 => n2607, A2 => n13866, B1 => n5868, B2 => 
                           n13863, C1 => n13857, C2 => n2196, ZN => n9119);
   U6298 : NOR4_X1 port map( A1 => n5869, A2 => n5870, A3 => n5871, A4 => n5872
                           , ZN => n5868);
   U6299 : NAND4_X1 port map( A1 => n5897, A2 => n5898, A3 => n5899, A4 => 
                           n5900, ZN => n5869);
   U6300 : NAND4_X1 port map( A1 => n5889, A2 => n5890, A3 => n5891, A4 => 
                           n5892, ZN => n5870);
   U6301 : OAI222_X1 port map( A1 => n2606, A2 => n14086, B1 => n4584, B2 => 
                           n14083, C1 => n14077, C2 => n2165, ZN => n9151);
   U6302 : NOR4_X1 port map( A1 => n4585, A2 => n4586, A3 => n4587, A4 => n4588
                           , ZN => n4584);
   U6303 : NAND4_X1 port map( A1 => n4613, A2 => n4614, A3 => n4615, A4 => 
                           n4616, ZN => n4585);
   U6304 : NAND4_X1 port map( A1 => n4605, A2 => n4606, A3 => n4607, A4 => 
                           n4608, ZN => n4586);
   U6305 : OAI222_X1 port map( A1 => n2606, A2 => n13866, B1 => n5905, B2 => 
                           n13863, C1 => n13857, C2 => n2197, ZN => n9118);
   U6306 : NOR4_X1 port map( A1 => n5906, A2 => n5907, A3 => n5908, A4 => n5909
                           , ZN => n5905);
   U6307 : NAND4_X1 port map( A1 => n5934, A2 => n5935, A3 => n5936, A4 => 
                           n5937, ZN => n5906);
   U6308 : NAND4_X1 port map( A1 => n5926, A2 => n5927, A3 => n5928, A4 => 
                           n5929, ZN => n5907);
   U6309 : OAI222_X1 port map( A1 => n2605, A2 => n14086, B1 => n4621, B2 => 
                           n14083, C1 => n14077, C2 => n2166, ZN => n9150);
   U6310 : NOR4_X1 port map( A1 => n4622, A2 => n4623, A3 => n4624, A4 => n4625
                           , ZN => n4621);
   U6311 : NAND4_X1 port map( A1 => n4650, A2 => n4651, A3 => n4652, A4 => 
                           n4653, ZN => n4622);
   U6312 : NAND4_X1 port map( A1 => n4642, A2 => n4643, A3 => n4644, A4 => 
                           n4645, ZN => n4623);
   U6313 : OAI222_X1 port map( A1 => n2605, A2 => n13866, B1 => n5942, B2 => 
                           n13863, C1 => n13857, C2 => n2198, ZN => n9117);
   U6314 : NOR4_X1 port map( A1 => n5943, A2 => n5944, A3 => n5945, A4 => n5946
                           , ZN => n5942);
   U6315 : NAND4_X1 port map( A1 => n5971, A2 => n5972, A3 => n5973, A4 => 
                           n5974, ZN => n5943);
   U6316 : NAND4_X1 port map( A1 => n5963, A2 => n5964, A3 => n5965, A4 => 
                           n5966, ZN => n5944);
   U6317 : OAI222_X1 port map( A1 => n2604, A2 => n14086, B1 => n4658, B2 => 
                           n14083, C1 => n14077, C2 => n2167, ZN => n9149);
   U6318 : NOR4_X1 port map( A1 => n4659, A2 => n4660, A3 => n4661, A4 => n4662
                           , ZN => n4658);
   U6319 : NAND4_X1 port map( A1 => n4687, A2 => n4688, A3 => n4689, A4 => 
                           n4690, ZN => n4659);
   U6320 : NAND4_X1 port map( A1 => n4679, A2 => n4680, A3 => n4681, A4 => 
                           n4682, ZN => n4660);
   U6321 : OAI222_X1 port map( A1 => n2604, A2 => n13866, B1 => n5979, B2 => 
                           n13863, C1 => n13857, C2 => n2199, ZN => n9116);
   U6322 : NOR4_X1 port map( A1 => n5980, A2 => n5981, A3 => n5982, A4 => n5983
                           , ZN => n5979);
   U6323 : NAND4_X1 port map( A1 => n6008, A2 => n6009, A3 => n6010, A4 => 
                           n6011, ZN => n5980);
   U6324 : NAND4_X1 port map( A1 => n6000, A2 => n6001, A3 => n6002, A4 => 
                           n6003, ZN => n5981);
   U6325 : AOI221_X1 port map( B1 => n13896, B2 => n8761, C1 => n13893, C2 => 
                           n8729, A => n4286, ZN => n4281);
   U6326 : OAI222_X1 port map( A1 => n1726, A2 => n13890, B1 => n6875, B2 => 
                           n13889, C1 => n59, C2 => n13884, ZN => n4286);
   U6327 : AOI221_X1 port map( B1 => n13720, B2 => n8448, C1 => n13717, C2 => 
                           n8416, A => n5414, ZN => n5409);
   U6328 : OAI222_X1 port map( A1 => n1756, A2 => n13714, B1 => n6761, B2 => 
                           n13711, C1 => n195, C2 => n13708, ZN => n5414);
   U6329 : AOI221_X1 port map( B1 => n13666, B2 => n8766, C1 => n13663, C2 => 
                           n8734, A => n5422, ZN => n5417);
   U6330 : OAI222_X1 port map( A1 => n1730, A2 => n13660, B1 => n6755, B2 => 
                           n13657, C1 => n64, C2 => n13654, ZN => n5422);
   U6331 : AOI221_X1 port map( B1 => n13720, B2 => n8446, C1 => n13717, C2 => 
                           n8414, A => n5488, ZN => n5483);
   U6332 : OAI222_X1 port map( A1 => n1755, A2 => n13714, B1 => n6809, B2 => 
                           n13711, C1 => n193, C2 => n13708, ZN => n5488);
   U6333 : AOI221_X1 port map( B1 => n13666, B2 => n8764, C1 => n13663, C2 => 
                           n8732, A => n5496, ZN => n5491);
   U6334 : OAI222_X1 port map( A1 => n1729, A2 => n13660, B1 => n6803, B2 => 
                           n13657, C1 => n62, C2 => n13654, ZN => n5496);
   U6335 : AOI221_X1 port map( B1 => n13720, B2 => n8445, C1 => n13717, C2 => 
                           n8413, A => n5525, ZN => n5520);
   U6336 : OAI222_X1 port map( A1 => n1754, A2 => n13714, B1 => n6833, B2 => 
                           n13711, C1 => n192, C2 => n13708, ZN => n5525);
   U6337 : AOI221_X1 port map( B1 => n13666, B2 => n8763, C1 => n13663, C2 => 
                           n8731, A => n5533, ZN => n5528);
   U6338 : OAI222_X1 port map( A1 => n1728, A2 => n13660, B1 => n6827, B2 => 
                           n13657, C1 => n61, C2 => n13654, ZN => n5533);
   U6339 : AOI221_X1 port map( B1 => n13720, B2 => n8444, C1 => n13717, C2 => 
                           n8412, A => n5562, ZN => n5557);
   U6340 : OAI222_X1 port map( A1 => n1753, A2 => n13714, B1 => n6857, B2 => 
                           n13711, C1 => n191, C2 => n13708, ZN => n5562);
   U6341 : AOI221_X1 port map( B1 => n13666, B2 => n8762, C1 => n13663, C2 => 
                           n8730, A => n5570, ZN => n5565);
   U6342 : OAI222_X1 port map( A1 => n1727, A2 => n13660, B1 => n6851, B2 => 
                           n13657, C1 => n60, C2 => n13654, ZN => n5570);
   U6343 : AOI221_X1 port map( B1 => n13720, B2 => n8443, C1 => n13717, C2 => 
                           n8411, A => n5599, ZN => n5594);
   U6344 : OAI222_X1 port map( A1 => n1752, A2 => n13714, B1 => n6881, B2 => 
                           n13711, C1 => n190, C2 => n13708, ZN => n5599);
   U6345 : AOI221_X1 port map( B1 => n13666, B2 => n8761, C1 => n13663, C2 => 
                           n8729, A => n5607, ZN => n5602);
   U6346 : OAI222_X1 port map( A1 => n1726, A2 => n13660, B1 => n6875, B2 => 
                           n13657, C1 => n59, C2 => n13654, ZN => n5607);
   U6347 : AOI221_X1 port map( B1 => n14046, B2 => n7972, C1 => n14043, C2 => 
                           n7940, A => n5197, ZN => n5182);
   U6348 : OAI222_X1 port map( A1 => n819, A2 => n14040, B1 => n966, B2 => 
                           n14037, C1 => n508, C2 => n14034, ZN => n5197);
   U6349 : AOI221_X1 port map( B1 => n8418, B2 => n13940, C1 => n8386, C2 => 
                           n13935, A => n5218, ZN => n5211);
   U6350 : OAI222_X1 port map( A1 => n13932, A2 => n2119, B1 => n7481, B2 => 
                           n13929, C1 => n13926, C2 => n2138, ZN => n5218);
   U6351 : AOI221_X1 port map( B1 => n13939, B2 => n8429, C1 => n13936, C2 => 
                           n8397, A => n4796, ZN => n4791);
   U6352 : OAI222_X1 port map( A1 => n2130, A2 => n13933, B1 => n2291, B2 => 
                           n13929, C1 => n2149, C2 => n13927, ZN => n4796);
   U6353 : AOI221_X1 port map( B1 => n14046, B2 => n7982, C1 => n14043, C2 => 
                           n7950, A => n4817, ZN => n4812);
   U6354 : OAI222_X1 port map( A1 => n924, A2 => n14040, B1 => n996, B2 => 
                           n14037, C1 => n518, C2 => n14034, ZN => n4817);
   U6355 : AOI221_X1 port map( B1 => n13939, B2 => n8428, C1 => n13936, C2 => 
                           n8396, A => n4833, ZN => n4828);
   U6356 : OAI222_X1 port map( A1 => n2129, A2 => n13933, B1 => n7241, B2 => 
                           n13929, C1 => n2148, C2 => n13927, ZN => n4833);
   U6357 : AOI221_X1 port map( B1 => n14046, B2 => n7981, C1 => n14043, C2 => 
                           n7949, A => n4854, ZN => n4849);
   U6358 : OAI222_X1 port map( A1 => n922, A2 => n14040, B1 => n994, B2 => 
                           n14037, C1 => n517, C2 => n14034, ZN => n4854);
   U6359 : AOI221_X1 port map( B1 => n13939, B2 => n8427, C1 => n13936, C2 => 
                           n8395, A => n4870, ZN => n4865);
   U6360 : OAI222_X1 port map( A1 => n2128, A2 => n13933, B1 => n7265, B2 => 
                           n13929, C1 => n2147, C2 => n13927, ZN => n4870);
   U6361 : AOI221_X1 port map( B1 => n14046, B2 => n7980, C1 => n14043, C2 => 
                           n7948, A => n4891, ZN => n4886);
   U6362 : OAI222_X1 port map( A1 => n918, A2 => n14040, B1 => n990, B2 => 
                           n14037, C1 => n516, C2 => n14034, ZN => n4891);
   U6363 : AOI221_X1 port map( B1 => n13939, B2 => n8426, C1 => n13936, C2 => 
                           n8394, A => n4907, ZN => n4902);
   U6364 : OAI222_X1 port map( A1 => n2127, A2 => n13933, B1 => n7289, B2 => 
                           n13929, C1 => n2146, C2 => n13927, ZN => n4907);
   U6365 : AOI221_X1 port map( B1 => n14046, B2 => n7979, C1 => n14043, C2 => 
                           n7947, A => n4928, ZN => n4923);
   U6366 : OAI222_X1 port map( A1 => n916, A2 => n14040, B1 => n988, B2 => 
                           n14037, C1 => n515, C2 => n14034, ZN => n4928);
   U6367 : AOI221_X1 port map( B1 => n13898, B2 => n8737, C1 => n13893, C2 => 
                           n8705, A => n5174, ZN => n5169);
   U6368 : OAI222_X1 port map( A1 => n2011, A2 => n13890, B1 => n7451, B2 => 
                           n13887, C1 => n2030, C2 => n13884, ZN => n5174);
   U6369 : AOI221_X1 port map( B1 => n13896, B2 => n8762, C1 => n13893, C2 => 
                           n8730, A => n4249, ZN => n4244);
   U6370 : OAI222_X1 port map( A1 => n1727, A2 => n13890, B1 => n6851, B2 => 
                           n13889, C1 => n60, C2 => n13884, ZN => n4249);
   U6371 : AOI221_X1 port map( B1 => n13939, B2 => n8425, C1 => n13937, C2 => 
                           n8393, A => n4944, ZN => n4939);
   U6372 : OAI222_X1 port map( A1 => n2126, A2 => n13934, B1 => n7313, B2 => 
                           n13929, C1 => n2145, C2 => n13928, ZN => n4944);
   U6373 : AOI221_X1 port map( B1 => n13897, B2 => n8743, C1 => n13895, C2 => 
                           n8711, A => n4952, ZN => n4947);
   U6374 : OAI222_X1 port map( A1 => n2017, A2 => n13892, B1 => n7307, B2 => 
                           n13887, C1 => n2036, C2 => n13886, ZN => n4952);
   U6375 : AOI221_X1 port map( B1 => n13718, B2 => n8429, C1 => n13715, C2 => 
                           n8397, A => n6117, ZN => n6112);
   U6376 : OAI222_X1 port map( A1 => n2130, A2 => n13712, B1 => n2291, B2 => 
                           n13709, C1 => n2149, C2 => n13706, ZN => n6117);
   U6377 : AOI221_X1 port map( B1 => n13664, B2 => n8747, C1 => n13661, C2 => 
                           n8715, A => n6125, ZN => n6120);
   U6378 : OAI222_X1 port map( A1 => n2021, A2 => n13658, B1 => n2054, B2 => 
                           n13655, C1 => n2040, C2 => n13652, ZN => n6125);
   U6379 : AOI221_X1 port map( B1 => n13826, B2 => n7982, C1 => n13823, C2 => 
                           n7950, A => n6138, ZN => n6133);
   U6380 : OAI222_X1 port map( A1 => n924, A2 => n13820, B1 => n996, B2 => 
                           n13817, C1 => n518, C2 => n13814, ZN => n6138);
   U6381 : AOI221_X1 port map( B1 => n13718, B2 => n8428, C1 => n13715, C2 => 
                           n8396, A => n6154, ZN => n6149);
   U6382 : OAI222_X1 port map( A1 => n2129, A2 => n13712, B1 => n7241, B2 => 
                           n13709, C1 => n2148, C2 => n13706, ZN => n6154);
   U6383 : AOI221_X1 port map( B1 => n13664, B2 => n8746, C1 => n13661, C2 => 
                           n8714, A => n6162, ZN => n6157);
   U6384 : OAI222_X1 port map( A1 => n2020, A2 => n13658, B1 => n2053, B2 => 
                           n13655, C1 => n2039, C2 => n13652, ZN => n6162);
   U6385 : AOI221_X1 port map( B1 => n13826, B2 => n7981, C1 => n13823, C2 => 
                           n7949, A => n6175, ZN => n6170);
   U6386 : OAI222_X1 port map( A1 => n922, A2 => n13820, B1 => n994, B2 => 
                           n13817, C1 => n517, C2 => n13814, ZN => n6175);
   U6387 : AOI221_X1 port map( B1 => n13718, B2 => n8427, C1 => n13715, C2 => 
                           n8395, A => n6191, ZN => n6186);
   U6388 : OAI222_X1 port map( A1 => n2128, A2 => n13712, B1 => n7265, B2 => 
                           n13709, C1 => n2147, C2 => n13706, ZN => n6191);
   U6389 : AOI221_X1 port map( B1 => n13664, B2 => n8745, C1 => n13661, C2 => 
                           n8713, A => n6199, ZN => n6194);
   U6390 : OAI222_X1 port map( A1 => n2019, A2 => n13658, B1 => n7259, B2 => 
                           n13655, C1 => n2038, C2 => n13652, ZN => n6199);
   U6391 : AOI221_X1 port map( B1 => n13826, B2 => n7980, C1 => n13823, C2 => 
                           n7948, A => n6212, ZN => n6207);
   U6392 : OAI222_X1 port map( A1 => n918, A2 => n13820, B1 => n990, B2 => 
                           n13817, C1 => n516, C2 => n13814, ZN => n6212);
   U6393 : AOI221_X1 port map( B1 => n13718, B2 => n8426, C1 => n13715, C2 => 
                           n8394, A => n6228, ZN => n6223);
   U6394 : OAI222_X1 port map( A1 => n2127, A2 => n13712, B1 => n7289, B2 => 
                           n13709, C1 => n2146, C2 => n13706, ZN => n6228);
   U6395 : AOI221_X1 port map( B1 => n13664, B2 => n8744, C1 => n13661, C2 => 
                           n8712, A => n6236, ZN => n6231);
   U6396 : OAI222_X1 port map( A1 => n2018, A2 => n13658, B1 => n7283, B2 => 
                           n13655, C1 => n2037, C2 => n13652, ZN => n6236);
   U6397 : AOI221_X1 port map( B1 => n13826, B2 => n7979, C1 => n13823, C2 => 
                           n7947, A => n6249, ZN => n6244);
   U6398 : OAI222_X1 port map( A1 => n916, A2 => n13820, B1 => n988, B2 => 
                           n13817, C1 => n515, C2 => n13814, ZN => n6249);
   U6399 : AOI221_X1 port map( B1 => n13718, B2 => n8425, C1 => n13715, C2 => 
                           n8393, A => n6265, ZN => n6260);
   U6400 : OAI222_X1 port map( A1 => n2126, A2 => n13712, B1 => n7313, B2 => 
                           n13709, C1 => n2145, C2 => n13706, ZN => n6265);
   U6401 : AOI221_X1 port map( B1 => n13664, B2 => n8743, C1 => n13661, C2 => 
                           n8711, A => n6273, ZN => n6268);
   U6402 : OAI222_X1 port map( A1 => n2017, A2 => n13658, B1 => n7307, B2 => 
                           n13655, C1 => n2036, C2 => n13652, ZN => n6273);
   U6403 : AOI221_X1 port map( B1 => n13826, B2 => n7978, C1 => n13823, C2 => 
                           n7946, A => n6286, ZN => n6281);
   U6404 : OAI222_X1 port map( A1 => n912, A2 => n13820, B1 => n984, B2 => 
                           n13817, C1 => n514, C2 => n13814, ZN => n6286);
   U6405 : AOI221_X1 port map( B1 => n13718, B2 => n8424, C1 => n13715, C2 => 
                           n8392, A => n6302, ZN => n6297);
   U6406 : OAI222_X1 port map( A1 => n2125, A2 => n13712, B1 => n7337, B2 => 
                           n13709, C1 => n2144, C2 => n13706, ZN => n6302);
   U6407 : AOI221_X1 port map( B1 => n13664, B2 => n8742, C1 => n13661, C2 => 
                           n8710, A => n6310, ZN => n6305);
   U6408 : OAI222_X1 port map( A1 => n2016, A2 => n13658, B1 => n7331, B2 => 
                           n13655, C1 => n2035, C2 => n13652, ZN => n6310);
   U6409 : AOI221_X1 port map( B1 => n13826, B2 => n7977, C1 => n13823, C2 => 
                           n7945, A => n6323, ZN => n6318);
   U6410 : OAI222_X1 port map( A1 => n910, A2 => n13820, B1 => n982, B2 => 
                           n13817, C1 => n513, C2 => n13814, ZN => n6323);
   U6411 : AOI221_X1 port map( B1 => n13718, B2 => n8423, C1 => n13715, C2 => 
                           n8391, A => n6339, ZN => n6334);
   U6412 : OAI222_X1 port map( A1 => n2124, A2 => n13712, B1 => n7361, B2 => 
                           n13709, C1 => n2143, C2 => n13706, ZN => n6339);
   U6413 : AOI221_X1 port map( B1 => n13664, B2 => n8741, C1 => n13661, C2 => 
                           n8709, A => n6347, ZN => n6342);
   U6414 : OAI222_X1 port map( A1 => n2015, A2 => n13658, B1 => n7355, B2 => 
                           n13655, C1 => n2034, C2 => n13652, ZN => n6347);
   U6415 : AOI221_X1 port map( B1 => n13826, B2 => n7976, C1 => n13823, C2 => 
                           n7944, A => n6360, ZN => n6355);
   U6416 : OAI222_X1 port map( A1 => n906, A2 => n13820, B1 => n978, B2 => 
                           n13817, C1 => n512, C2 => n13814, ZN => n6360);
   U6417 : AOI221_X1 port map( B1 => n13718, B2 => n8422, C1 => n13715, C2 => 
                           n8390, A => n6376, ZN => n6371);
   U6418 : OAI222_X1 port map( A1 => n2123, A2 => n13712, B1 => n7385, B2 => 
                           n13709, C1 => n2142, C2 => n13706, ZN => n6376);
   U6419 : AOI221_X1 port map( B1 => n13664, B2 => n8740, C1 => n13661, C2 => 
                           n8708, A => n6384, ZN => n6379);
   U6420 : OAI222_X1 port map( A1 => n2014, A2 => n13658, B1 => n7379, B2 => 
                           n13655, C1 => n2033, C2 => n13652, ZN => n6384);
   U6421 : AOI221_X1 port map( B1 => n13826, B2 => n7975, C1 => n13823, C2 => 
                           n7943, A => n6397, ZN => n6392);
   U6422 : OAI222_X1 port map( A1 => n904, A2 => n13820, B1 => n976, B2 => 
                           n13817, C1 => n511, C2 => n13814, ZN => n6397);
   U6423 : AOI221_X1 port map( B1 => n13718, B2 => n8421, C1 => n13715, C2 => 
                           n8389, A => n6413, ZN => n6408);
   U6424 : OAI222_X1 port map( A1 => n2122, A2 => n13712, B1 => n7409, B2 => 
                           n13709, C1 => n2141, C2 => n13706, ZN => n6413);
   U6425 : AOI221_X1 port map( B1 => n13664, B2 => n8739, C1 => n13661, C2 => 
                           n8707, A => n6421, ZN => n6416);
   U6426 : OAI222_X1 port map( A1 => n2013, A2 => n13658, B1 => n7403, B2 => 
                           n13655, C1 => n2032, C2 => n13652, ZN => n6421);
   U6427 : AOI221_X1 port map( B1 => n13826, B2 => n7974, C1 => n13823, C2 => 
                           n7942, A => n6434, ZN => n6429);
   U6428 : OAI222_X1 port map( A1 => n900, A2 => n13820, B1 => n972, B2 => 
                           n13817, C1 => n510, C2 => n13814, ZN => n6434);
   U6429 : AOI221_X1 port map( B1 => n13718, B2 => n8420, C1 => n13715, C2 => 
                           n8388, A => n6450, ZN => n6445);
   U6430 : OAI222_X1 port map( A1 => n2121, A2 => n13712, B1 => n7433, B2 => 
                           n13709, C1 => n2140, C2 => n13706, ZN => n6450);
   U6431 : AOI221_X1 port map( B1 => n13664, B2 => n8738, C1 => n13661, C2 => 
                           n8706, A => n6458, ZN => n6453);
   U6432 : OAI222_X1 port map( A1 => n2012, A2 => n13658, B1 => n7427, B2 => 
                           n13655, C1 => n2031, C2 => n13652, ZN => n6458);
   U6433 : AOI221_X1 port map( B1 => n13826, B2 => n7973, C1 => n13823, C2 => 
                           n7941, A => n6471, ZN => n6466);
   U6434 : OAI222_X1 port map( A1 => n898, A2 => n13820, B1 => n970, B2 => 
                           n13817, C1 => n509, C2 => n13814, ZN => n6471);
   U6435 : AOI221_X1 port map( B1 => n13718, B2 => n8419, C1 => n13715, C2 => 
                           n8387, A => n6487, ZN => n6482);
   U6436 : OAI222_X1 port map( A1 => n2120, A2 => n13712, B1 => n7457, B2 => 
                           n13709, C1 => n2139, C2 => n13706, ZN => n6487);
   U6437 : AOI221_X1 port map( B1 => n13664, B2 => n8737, C1 => n13661, C2 => 
                           n8705, A => n6495, ZN => n6490);
   U6438 : OAI222_X1 port map( A1 => n2011, A2 => n13658, B1 => n7451, B2 => 
                           n13655, C1 => n2030, C2 => n13652, ZN => n6495);
   U6439 : AOI221_X1 port map( B1 => n14047, B2 => n7985, C1 => n14044, C2 => 
                           n7953, A => n4706, ZN => n4701);
   U6440 : OAI222_X1 port map( A1 => n934, A2 => n14041, B1 => n1002, B2 => 
                           n14038, C1 => n521, C2 => n14035, ZN => n4706);
   U6441 : AOI221_X1 port map( B1 => n13897, B2 => n8749, C1 => n13894, C2 => 
                           n8717, A => n4730, ZN => n4725);
   U6442 : OAI222_X1 port map( A1 => n2023, A2 => n13891, B1 => n7163, B2 => 
                           n13888, C1 => n2042, C2 => n13885, ZN => n4730);
   U6443 : AOI221_X1 port map( B1 => n13897, B2 => n8748, C1 => n13894, C2 => 
                           n8716, A => n4767, ZN => n4762);
   U6444 : OAI222_X1 port map( A1 => n2022, A2 => n13891, B1 => n7187, B2 => 
                           n13888, C1 => n2041, C2 => n13885, ZN => n4767);
   U6445 : AOI221_X1 port map( B1 => n13827, B2 => n7985, C1 => n13824, C2 => 
                           n7953, A => n6027, ZN => n6022);
   U6446 : OAI222_X1 port map( A1 => n934, A2 => n13821, B1 => n1002, B2 => 
                           n13818, C1 => n521, C2 => n13815, ZN => n6027);
   U6447 : AOI221_X1 port map( B1 => n13719, B2 => n8431, C1 => n13716, C2 => 
                           n8399, A => n6043, ZN => n6038);
   U6448 : OAI222_X1 port map( A1 => n2132, A2 => n13713, B1 => n7169, B2 => 
                           n13710, C1 => n2279, C2 => n13707, ZN => n6043);
   U6449 : AOI221_X1 port map( B1 => n13665, B2 => n8749, C1 => n13662, C2 => 
                           n8717, A => n6051, ZN => n6046);
   U6450 : OAI222_X1 port map( A1 => n2023, A2 => n13659, B1 => n7163, B2 => 
                           n13656, C1 => n2042, C2 => n13653, ZN => n6051);
   U6451 : AOI221_X1 port map( B1 => n13719, B2 => n8430, C1 => n13716, C2 => 
                           n8398, A => n6080, ZN => n6075);
   U6452 : OAI222_X1 port map( A1 => n2131, A2 => n13713, B1 => n7193, B2 => 
                           n13710, C1 => n2278, C2 => n13707, ZN => n6080);
   U6453 : AOI221_X1 port map( B1 => n13665, B2 => n8748, C1 => n13662, C2 => 
                           n8716, A => n6088, ZN => n6083);
   U6454 : OAI222_X1 port map( A1 => n2022, A2 => n13659, B1 => n7187, B2 => 
                           n13656, C1 => n2041, C2 => n13653, ZN => n6088);
   U6455 : AOI221_X1 port map( B1 => n13826, B2 => n7972, C1 => n13823, C2 => 
                           n7940, A => n6518, ZN => n6503);
   U6456 : OAI222_X1 port map( A1 => n819, A2 => n13820, B1 => n966, B2 => 
                           n13817, C1 => n508, C2 => n13814, ZN => n6518);
   U6457 : AOI221_X1 port map( B1 => n13718, B2 => n8418, C1 => n13715, C2 => 
                           n8386, A => n6539, ZN => n6532);
   U6458 : OAI222_X1 port map( A1 => n2119, A2 => n13712, B1 => n7481, B2 => 
                           n13709, C1 => n2138, C2 => n13706, ZN => n6539);
   U6459 : AOI221_X1 port map( B1 => n13664, B2 => n8736, C1 => n13661, C2 => 
                           n8704, A => n6548, ZN => n6542);
   U6460 : OAI222_X1 port map( A1 => n2010, A2 => n13658, B1 => n7475, B2 => 
                           n13655, C1 => n2029, C2 => n13652, ZN => n6548);
   U6461 : AOI221_X1 port map( B1 => n14046, B2 => n7978, C1 => n14043, C2 => 
                           n7946, A => n4965, ZN => n4960);
   U6462 : OAI222_X1 port map( A1 => n912, A2 => n14040, B1 => n984, B2 => 
                           n14037, C1 => n514, C2 => n14034, ZN => n4965);
   U6463 : AOI221_X1 port map( B1 => n13940, B2 => n8424, C1 => n13937, C2 => 
                           n8392, A => n4981, ZN => n4976);
   U6464 : OAI222_X1 port map( A1 => n2125, A2 => n13934, B1 => n7337, B2 => 
                           n13929, C1 => n2144, C2 => n13928, ZN => n4981);
   U6465 : AOI221_X1 port map( B1 => n13898, B2 => n8742, C1 => n13895, C2 => 
                           n8710, A => n4989, ZN => n4984);
   U6466 : OAI222_X1 port map( A1 => n2016, A2 => n13892, B1 => n7331, B2 => 
                           n13887, C1 => n2035, C2 => n13886, ZN => n4989);
   U6467 : AOI221_X1 port map( B1 => n14046, B2 => n7977, C1 => n14043, C2 => 
                           n7945, A => n5002, ZN => n4997);
   U6468 : OAI222_X1 port map( A1 => n910, A2 => n14040, B1 => n982, B2 => 
                           n14037, C1 => n513, C2 => n14034, ZN => n5002);
   U6469 : AOI221_X1 port map( B1 => n13940, B2 => n8423, C1 => n13937, C2 => 
                           n8391, A => n5018, ZN => n5013);
   U6470 : OAI222_X1 port map( A1 => n2124, A2 => n13934, B1 => n7361, B2 => 
                           n13929, C1 => n2143, C2 => n13928, ZN => n5018);
   U6471 : AOI221_X1 port map( B1 => n13898, B2 => n8741, C1 => n13895, C2 => 
                           n8709, A => n5026, ZN => n5021);
   U6472 : OAI222_X1 port map( A1 => n2015, A2 => n13892, B1 => n7355, B2 => 
                           n13887, C1 => n2034, C2 => n13886, ZN => n5026);
   U6473 : AOI221_X1 port map( B1 => n14046, B2 => n7976, C1 => n14043, C2 => 
                           n7944, A => n5039, ZN => n5034);
   U6474 : OAI222_X1 port map( A1 => n906, A2 => n14040, B1 => n978, B2 => 
                           n14037, C1 => n512, C2 => n14034, ZN => n5039);
   U6475 : AOI221_X1 port map( B1 => n13940, B2 => n8422, C1 => n13937, C2 => 
                           n8390, A => n5055, ZN => n5050);
   U6476 : OAI222_X1 port map( A1 => n2123, A2 => n13934, B1 => n7385, B2 => 
                           n13929, C1 => n2142, C2 => n13928, ZN => n5055);
   U6477 : AOI221_X1 port map( B1 => n13898, B2 => n8740, C1 => n13895, C2 => 
                           n8708, A => n5063, ZN => n5058);
   U6478 : OAI222_X1 port map( A1 => n2014, A2 => n13892, B1 => n7379, B2 => 
                           n13887, C1 => n2033, C2 => n13886, ZN => n5063);
   U6479 : AOI221_X1 port map( B1 => n14046, B2 => n7975, C1 => n14043, C2 => 
                           n7943, A => n5076, ZN => n5071);
   U6480 : OAI222_X1 port map( A1 => n904, A2 => n14040, B1 => n976, B2 => 
                           n14037, C1 => n511, C2 => n14034, ZN => n5076);
   U6481 : AOI221_X1 port map( B1 => n13940, B2 => n8421, C1 => n13937, C2 => 
                           n8389, A => n5092, ZN => n5087);
   U6482 : OAI222_X1 port map( A1 => n2122, A2 => n13934, B1 => n7409, B2 => 
                           n13929, C1 => n2141, C2 => n13928, ZN => n5092);
   U6483 : AOI221_X1 port map( B1 => n13898, B2 => n8739, C1 => n13895, C2 => 
                           n8707, A => n5100, ZN => n5095);
   U6484 : OAI222_X1 port map( A1 => n2013, A2 => n13892, B1 => n7403, B2 => 
                           n13887, C1 => n2032, C2 => n13886, ZN => n5100);
   U6485 : AOI221_X1 port map( B1 => n14046, B2 => n7974, C1 => n14043, C2 => 
                           n7942, A => n5113, ZN => n5108);
   U6486 : OAI222_X1 port map( A1 => n900, A2 => n14040, B1 => n972, B2 => 
                           n14037, C1 => n510, C2 => n14034, ZN => n5113);
   U6487 : AOI221_X1 port map( B1 => n13940, B2 => n8420, C1 => n13937, C2 => 
                           n8388, A => n5129, ZN => n5124);
   U6488 : OAI222_X1 port map( A1 => n2121, A2 => n13934, B1 => n7433, B2 => 
                           n13929, C1 => n2140, C2 => n13928, ZN => n5129);
   U6489 : AOI221_X1 port map( B1 => n13898, B2 => n8738, C1 => n13895, C2 => 
                           n8706, A => n5137, ZN => n5132);
   U6490 : OAI222_X1 port map( A1 => n2012, A2 => n13892, B1 => n7427, B2 => 
                           n13887, C1 => n2031, C2 => n13886, ZN => n5137);
   U6491 : AOI221_X1 port map( B1 => n14046, B2 => n7973, C1 => n14043, C2 => 
                           n7941, A => n5150, ZN => n5145);
   U6492 : OAI222_X1 port map( A1 => n898, A2 => n14040, B1 => n970, B2 => 
                           n14037, C1 => n509, C2 => n14034, ZN => n5150);
   U6493 : AOI221_X1 port map( B1 => n14048, B2 => n8003, C1 => n14045, C2 => 
                           n7971, A => n3979, ZN => n3963);
   U6494 : OAI222_X1 port map( A1 => n316, A2 => n14042, B1 => n332, B2 => 
                           n14039, C1 => n324, C2 => n14036, ZN => n3979);
   U6495 : AOI221_X1 port map( B1 => n8767, B2 => n13898, C1 => n8735, C2 => 
                           n13893, A => n4055, ZN => n4039);
   U6496 : OAI222_X1 port map( A1 => n13890, A2 => n1731, B1 => n6731, B2 => 
                           n13889, C1 => n13884, C2 => n1732, ZN => n4055);
   U6497 : AOI221_X1 port map( B1 => n13828, B2 => n8003, C1 => n13825, C2 => 
                           n7971, A => n5300, ZN => n5284);
   U6498 : OAI222_X1 port map( A1 => n316, A2 => n13822, B1 => n332, B2 => 
                           n13819, C1 => n324, C2 => n13816, ZN => n5300);
   U6499 : AOI221_X1 port map( B1 => n13720, B2 => n8449, C1 => n13717, C2 => 
                           n8417, A => n5352, ZN => n5336);
   U6500 : OAI222_X1 port map( A1 => n1757, A2 => n13714, B1 => n6737, B2 => 
                           n13711, C1 => n1758, C2 => n13708, ZN => n5352);
   U6501 : AOI221_X1 port map( B1 => n13666, B2 => n8767, C1 => n13663, C2 => 
                           n8735, A => n5378, ZN => n5362);
   U6502 : OAI222_X1 port map( A1 => n1731, A2 => n13660, B1 => n6731, B2 => 
                           n13657, C1 => n1732, C2 => n13654, ZN => n5378);
   U6503 : AOI221_X1 port map( B1 => n14112, B2 => n1854, C1 => n14109, C2 => 
                           n832, A => n6602, ZN => n6596);
   U6504 : OAI222_X1 port map( A1 => n308, A2 => n14106, B1 => n7682, B2 => 
                           n14103, C1 => n300, C2 => n14100, ZN => n6602);
   U6505 : AOI221_X1 port map( B1 => n13896, B2 => n8766, C1 => n13893, C2 => 
                           n8734, A => n4101, ZN => n4096);
   U6506 : OAI222_X1 port map( A1 => n1730, A2 => n13890, B1 => n6755, B2 => 
                           n13889, C1 => n64, C2 => n13884, ZN => n4101);
   U6507 : AOI221_X1 port map( B1 => n14114, B2 => n1853, C1 => n14111, C2 => 
                           n834, A => n2869, ZN => n2860);
   U6508 : OAI222_X1 port map( A1 => n307, A2 => n14108, B1 => n7676, B2 => 
                           n14105, C1 => n299, C2 => n14102, ZN => n2869);
   U6509 : AOI221_X1 port map( B1 => n13896, B2 => n8765, C1 => n13893, C2 => 
                           n8733, A => n4138, ZN => n4133);
   U6510 : OAI222_X1 port map( A1 => n57, A2 => n13890, B1 => n6779, B2 => 
                           n13889, C1 => n63, C2 => n13884, ZN => n4138);
   U6511 : AOI221_X1 port map( B1 => n13720, B2 => n8447, C1 => n13717, C2 => 
                           n8415, A => n5451, ZN => n5446);
   U6512 : OAI222_X1 port map( A1 => n188, A2 => n13714, B1 => n6785, B2 => 
                           n13711, C1 => n194, C2 => n13708, ZN => n5451);
   U6513 : AOI221_X1 port map( B1 => n13666, B2 => n8765, C1 => n13663, C2 => 
                           n8733, A => n5459, ZN => n5454);
   U6514 : OAI222_X1 port map( A1 => n57, A2 => n13660, B1 => n6779, B2 => 
                           n13657, C1 => n63, C2 => n13654, ZN => n5459);
   U6515 : AOI221_X1 port map( B1 => n14114, B2 => n1852, C1 => n14111, C2 => 
                           n836, A => n2913, ZN => n2908);
   U6516 : OAI222_X1 port map( A1 => n306, A2 => n14108, B1 => n7670, B2 => 
                           n14105, C1 => n298, C2 => n14102, ZN => n2913);
   U6517 : AOI221_X1 port map( B1 => n13896, B2 => n8764, C1 => n13893, C2 => 
                           n8732, A => n4175, ZN => n4170);
   U6518 : OAI222_X1 port map( A1 => n1729, A2 => n13890, B1 => n6803, B2 => 
                           n13889, C1 => n62, C2 => n13884, ZN => n4175);
   U6519 : AOI221_X1 port map( B1 => n14114, B2 => n1851, C1 => n14111, C2 => 
                           n838, A => n2950, ZN => n2945);
   U6520 : OAI222_X1 port map( A1 => n305, A2 => n14108, B1 => n7664, B2 => 
                           n14105, C1 => n297, C2 => n14102, ZN => n2950);
   U6521 : AOI221_X1 port map( B1 => n13896, B2 => n8763, C1 => n13893, C2 => 
                           n8731, A => n4212, ZN => n4207);
   U6522 : OAI222_X1 port map( A1 => n1728, A2 => n13890, B1 => n6827, B2 => 
                           n13889, C1 => n61, C2 => n13884, ZN => n4212);
   U6523 : AOI221_X1 port map( B1 => n14114, B2 => n1850, C1 => n14111, C2 => 
                           n840, A => n2987, ZN => n2982);
   U6524 : OAI222_X1 port map( A1 => n304, A2 => n14108, B1 => n7658, B2 => 
                           n14105, C1 => n296, C2 => n14102, ZN => n2987);
   U6525 : AOI221_X1 port map( B1 => n14114, B2 => n1849, C1 => n14111, C2 => 
                           n842, A => n3024, ZN => n3019);
   U6526 : OAI222_X1 port map( A1 => n303, A2 => n14108, B1 => n7652, B2 => 
                           n14105, C1 => n295, C2 => n14102, ZN => n3024);
   U6527 : AOI221_X1 port map( B1 => n14114, B2 => n1848, C1 => n14111, C2 => 
                           n844, A => n3061, ZN => n3056);
   U6528 : OAI222_X1 port map( A1 => n302, A2 => n14108, B1 => n7646, B2 => 
                           n14105, C1 => n294, C2 => n14102, ZN => n3061);
   U6529 : AOI221_X1 port map( B1 => n13896, B2 => n8760, C1 => n13893, C2 => 
                           n8728, A => n4323, ZN => n4318);
   U6530 : OAI222_X1 port map( A1 => n1725, A2 => n13890, B1 => n6899, B2 => 
                           n13889, C1 => n58, C2 => n13884, ZN => n4323);
   U6531 : AOI221_X1 port map( B1 => n13720, B2 => n8442, C1 => n13717, C2 => 
                           n8410, A => n5636, ZN => n5631);
   U6532 : OAI222_X1 port map( A1 => n1751, A2 => n13714, B1 => n6905, B2 => 
                           n13711, C1 => n189, C2 => n13708, ZN => n5636);
   U6533 : AOI221_X1 port map( B1 => n13666, B2 => n8760, C1 => n13663, C2 => 
                           n8728, A => n5644, ZN => n5639);
   U6534 : OAI222_X1 port map( A1 => n1725, A2 => n13660, B1 => n6899, B2 => 
                           n13657, C1 => n58, C2 => n13654, ZN => n5644);
   U6535 : AOI221_X1 port map( B1 => n13897, B2 => n8759, C1 => n13894, C2 => 
                           n8727, A => n4360, ZN => n4355);
   U6536 : OAI222_X1 port map( A1 => n2028, A2 => n13891, B1 => n6923, B2 => 
                           n13888, C1 => n1144, C2 => n13885, ZN => n4360);
   U6537 : AOI221_X1 port map( B1 => n13665, B2 => n8759, C1 => n13662, C2 => 
                           n8727, A => n5681, ZN => n5676);
   U6538 : OAI222_X1 port map( A1 => n2028, A2 => n13659, B1 => n6923, B2 => 
                           n13656, C1 => n1144, C2 => n13653, ZN => n5681);
   U6539 : AOI221_X1 port map( B1 => n13896, B2 => n8758, C1 => n13893, C2 => 
                           n8726, A => n4397, ZN => n4392);
   U6540 : OAI222_X1 port map( A1 => n2027, A2 => n13890, B1 => n6947, B2 => 
                           n13888, C1 => n1143, C2 => n13884, ZN => n4397);
   U6541 : AOI221_X1 port map( B1 => n14113, B2 => n2428, C1 => n14110, C2 => 
                           n852, A => n3209, ZN => n3204);
   U6542 : OAI222_X1 port map( A1 => n808, A2 => n14107, B1 => n7622, B2 => 
                           n14104, C1 => n505, C2 => n14101, ZN => n3209);
   U6543 : AOI221_X1 port map( B1 => n13896, B2 => n8756, C1 => n13893, C2 => 
                           n8724, A => n4471, ZN => n4466);
   U6544 : OAI222_X1 port map( A1 => n2025, A2 => n13890, B1 => n6995, B2 => 
                           n13888, C1 => n1141, C2 => n13884, ZN => n4471);
   U6545 : AOI221_X1 port map( B1 => n13719, B2 => n8438, C1 => n13716, C2 => 
                           n8406, A => n5784, ZN => n5779);
   U6546 : OAI222_X1 port map( A1 => n2134, A2 => n13713, B1 => n7001, B2 => 
                           n13710, C1 => n1459, C2 => n13707, ZN => n5784);
   U6547 : AOI221_X1 port map( B1 => n13665, B2 => n8756, C1 => n13662, C2 => 
                           n8724, A => n5792, ZN => n5787);
   U6548 : OAI222_X1 port map( A1 => n2025, A2 => n13659, B1 => n6995, B2 => 
                           n13656, C1 => n1141, C2 => n13653, ZN => n5792);
   U6549 : AOI221_X1 port map( B1 => n14113, B2 => n2427, C1 => n14110, C2 => 
                           n854, A => n3246, ZN => n3241);
   U6550 : OAI222_X1 port map( A1 => n804, A2 => n14107, B1 => n7616, B2 => 
                           n14104, C1 => n504, C2 => n14101, ZN => n3246);
   U6551 : AOI221_X1 port map( B1 => n13896, B2 => n8755, C1 => n13894, C2 => 
                           n8723, A => n4508, ZN => n4503);
   U6552 : OAI222_X1 port map( A1 => n2024, A2 => n13891, B1 => n7019, B2 => 
                           n13888, C1 => n1140, C2 => n13885, ZN => n4508);
   U6553 : AOI221_X1 port map( B1 => n13719, B2 => n8437, C1 => n13716, C2 => 
                           n8405, A => n5821, ZN => n5816);
   U6554 : OAI222_X1 port map( A1 => n2133, A2 => n13713, B1 => n7025, B2 => 
                           n13710, C1 => n1458, C2 => n13707, ZN => n5821);
   U6555 : AOI221_X1 port map( B1 => n13665, B2 => n8755, C1 => n13662, C2 => 
                           n8723, A => n5829, ZN => n5824);
   U6556 : OAI222_X1 port map( A1 => n2024, A2 => n13659, B1 => n7019, B2 => 
                           n13656, C1 => n1140, C2 => n13653, ZN => n5829);
   U6557 : AOI221_X1 port map( B1 => n14113, B2 => n2426, C1 => n14110, C2 => 
                           n856, A => n3283, ZN => n3278);
   U6558 : OAI222_X1 port map( A1 => n797, A2 => n14107, B1 => n7610, B2 => 
                           n14104, C1 => n503, C2 => n14101, ZN => n3283);
   U6559 : AOI221_X1 port map( B1 => n13896, B2 => n8754, C1 => n13894, C2 => 
                           n8722, A => n4545, ZN => n4540);
   U6560 : OAI222_X1 port map( A1 => n1134, A2 => n13891, B1 => n7043, B2 => 
                           n13888, C1 => n1139, C2 => n13885, ZN => n4545);
   U6561 : AOI221_X1 port map( B1 => n13719, B2 => n8436, C1 => n13716, C2 => 
                           n8404, A => n5858, ZN => n5853);
   U6562 : OAI222_X1 port map( A1 => n1452, A2 => n13713, B1 => n7049, B2 => 
                           n13710, C1 => n1457, C2 => n13707, ZN => n5858);
   U6563 : AOI221_X1 port map( B1 => n13665, B2 => n8754, C1 => n13662, C2 => 
                           n8722, A => n5866, ZN => n5861);
   U6564 : OAI222_X1 port map( A1 => n1134, A2 => n13659, B1 => n7043, B2 => 
                           n13656, C1 => n1139, C2 => n13653, ZN => n5866);
   U6565 : AOI221_X1 port map( B1 => n14113, B2 => n2425, C1 => n14110, C2 => 
                           n858, A => n3322, ZN => n3317);
   U6566 : OAI222_X1 port map( A1 => n796, A2 => n14107, B1 => n7604, B2 => 
                           n14104, C1 => n502, C2 => n14101, ZN => n3322);
   U6567 : AOI221_X1 port map( B1 => n13897, B2 => n8753, C1 => n13894, C2 => 
                           n8721, A => n4582, ZN => n4577);
   U6568 : OAI222_X1 port map( A1 => n1133, A2 => n13891, B1 => n7067, B2 => 
                           n13888, C1 => n1138, C2 => n13885, ZN => n4582);
   U6569 : AOI221_X1 port map( B1 => n13719, B2 => n8435, C1 => n13716, C2 => 
                           n8403, A => n5895, ZN => n5890);
   U6570 : OAI222_X1 port map( A1 => n1451, A2 => n13713, B1 => n7073, B2 => 
                           n13710, C1 => n1456, C2 => n13707, ZN => n5895);
   U6571 : AOI221_X1 port map( B1 => n13665, B2 => n8753, C1 => n13662, C2 => 
                           n8721, A => n5903, ZN => n5898);
   U6572 : OAI222_X1 port map( A1 => n1133, A2 => n13659, B1 => n7067, B2 => 
                           n13656, C1 => n1138, C2 => n13653, ZN => n5903);
   U6573 : AOI221_X1 port map( B1 => n14113, B2 => n2424, C1 => n14110, C2 => 
                           n860, A => n3359, ZN => n3354);
   U6574 : OAI222_X1 port map( A1 => n794, A2 => n14107, B1 => n7598, B2 => 
                           n14104, C1 => n501, C2 => n14101, ZN => n3359);
   U6575 : AOI221_X1 port map( B1 => n13897, B2 => n8752, C1 => n13894, C2 => 
                           n8720, A => n4619, ZN => n4614);
   U6576 : OAI222_X1 port map( A1 => n1132, A2 => n13891, B1 => n7091, B2 => 
                           n13888, C1 => n1137, C2 => n13885, ZN => n4619);
   U6577 : AOI221_X1 port map( B1 => n13719, B2 => n8434, C1 => n13716, C2 => 
                           n8402, A => n5932, ZN => n5927);
   U6578 : OAI222_X1 port map( A1 => n1450, A2 => n13713, B1 => n7097, B2 => 
                           n13710, C1 => n1455, C2 => n13707, ZN => n5932);
   U6579 : AOI221_X1 port map( B1 => n13665, B2 => n8752, C1 => n13662, C2 => 
                           n8720, A => n5940, ZN => n5935);
   U6580 : OAI222_X1 port map( A1 => n1132, A2 => n13659, B1 => n7091, B2 => 
                           n13656, C1 => n1137, C2 => n13653, ZN => n5940);
   U6581 : AOI221_X1 port map( B1 => n14113, B2 => n2423, C1 => n14110, C2 => 
                           n862, A => n3396, ZN => n3391);
   U6582 : OAI222_X1 port map( A1 => n793, A2 => n14107, B1 => n7592, B2 => 
                           n14104, C1 => n500, C2 => n14101, ZN => n3396);
   U6583 : AOI221_X1 port map( B1 => n13897, B2 => n8751, C1 => n13894, C2 => 
                           n8719, A => n4656, ZN => n4651);
   U6584 : OAI222_X1 port map( A1 => n1131, A2 => n13891, B1 => n7115, B2 => 
                           n13888, C1 => n1136, C2 => n13885, ZN => n4656);
   U6585 : AOI221_X1 port map( B1 => n13719, B2 => n8433, C1 => n13716, C2 => 
                           n8401, A => n5969, ZN => n5964);
   U6586 : OAI222_X1 port map( A1 => n1449, A2 => n13713, B1 => n7121, B2 => 
                           n13710, C1 => n1454, C2 => n13707, ZN => n5969);
   U6587 : AOI221_X1 port map( B1 => n13665, B2 => n8751, C1 => n13662, C2 => 
                           n8719, A => n5977, ZN => n5972);
   U6588 : OAI222_X1 port map( A1 => n1131, A2 => n13659, B1 => n7115, B2 => 
                           n13656, C1 => n1136, C2 => n13653, ZN => n5977);
   U6589 : AOI221_X1 port map( B1 => n14113, B2 => n2422, C1 => n14110, C2 => 
                           n864, A => n3433, ZN => n3428);
   U6590 : OAI222_X1 port map( A1 => n792, A2 => n14107, B1 => n7586, B2 => 
                           n14104, C1 => n499, C2 => n14101, ZN => n3433);
   U6591 : AOI221_X1 port map( B1 => n13897, B2 => n8750, C1 => n13894, C2 => 
                           n8718, A => n4693, ZN => n4688);
   U6592 : OAI222_X1 port map( A1 => n1130, A2 => n13891, B1 => n7139, B2 => 
                           n13888, C1 => n1135, C2 => n13885, ZN => n4693);
   U6593 : AOI221_X1 port map( B1 => n13719, B2 => n8432, C1 => n13716, C2 => 
                           n8400, A => n6006, ZN => n6001);
   U6594 : OAI222_X1 port map( A1 => n1448, A2 => n13713, B1 => n7145, B2 => 
                           n13710, C1 => n1453, C2 => n13707, ZN => n6006);
   U6595 : AOI221_X1 port map( B1 => n13665, B2 => n8750, C1 => n13662, C2 => 
                           n8718, A => n6014, ZN => n6009);
   U6596 : OAI222_X1 port map( A1 => n1130, A2 => n13659, B1 => n7139, B2 => 
                           n13656, C1 => n1135, C2 => n13653, ZN => n6014);
   U6597 : AOI221_X1 port map( B1 => n14113, B2 => n2421, C1 => n14110, C2 => 
                           n866, A => n3470, ZN => n3465);
   U6598 : OAI222_X1 port map( A1 => n790, A2 => n14107, B1 => n7580, B2 => 
                           n14104, C1 => n498, C2 => n14101, ZN => n3470);
   U6599 : AOI221_X1 port map( B1 => n14113, B2 => n2420, C1 => n14110, C2 => 
                           n868, A => n3507, ZN => n3502);
   U6600 : OAI222_X1 port map( A1 => n789, A2 => n14107, B1 => n7574, B2 => 
                           n14104, C1 => n497, C2 => n14101, ZN => n3507);
   U6601 : AOI221_X1 port map( B1 => n14113, B2 => n816, C1 => n14110, C2 => 
                           n870, A => n3544, ZN => n3539);
   U6602 : OAI222_X1 port map( A1 => n810, A2 => n14107, B1 => n1868, B2 => 
                           n14104, C1 => n811, C2 => n14101, ZN => n3544);
   U6603 : AOI221_X1 port map( B1 => n770, B2 => n14145, C1 => n14141, C2 => 
                           n1976, A => n3573, ZN => n3568);
   U6604 : OAI222_X1 port map( A1 => n14138, A2 => n1073, B1 => n7848, B2 => 
                           n14134, C1 => n14132, C2 => n1094, ZN => n3573);
   U6605 : AOI221_X1 port map( B1 => n14113, B2 => n752, C1 => n14110, C2 => 
                           n872, A => n3581, ZN => n3576);
   U6606 : OAI222_X1 port map( A1 => n787, A2 => n14107, B1 => n7562, B2 => 
                           n14104, C1 => n495, C2 => n14101, ZN => n3581);
   U6607 : AOI221_X1 port map( B1 => n14143, B2 => n1791, C1 => n14140, C2 => 
                           n1806, A => n6593, ZN => n6587);
   U6608 : OAI222_X1 port map( A1 => n14137, A2 => n260, B1 => n14134, B2 => 
                           n252, C1 => n14131, C2 => n268, ZN => n6593);
   U6609 : AOI221_X1 port map( B1 => n14144, B2 => n1790, C1 => n14142, C2 => 
                           n1805, A => n2850, ZN => n2836);
   U6610 : OAI222_X1 port map( A1 => n14138, A2 => n259, B1 => n7905, B2 => 
                           n14136, C1 => n14132, C2 => n267, ZN => n2850);
   U6611 : AOI221_X1 port map( B1 => n14143, B2 => n1789, C1 => n14142, C2 => 
                           n1804, A => n2905, ZN => n2900);
   U6612 : OAI222_X1 port map( A1 => n14137, A2 => n258, B1 => n7902, B2 => 
                           n14136, C1 => n14131, C2 => n266, ZN => n2905);
   U6613 : AOI221_X1 port map( B1 => n14143, B2 => n1788, C1 => n14142, C2 => 
                           n1803, A => n2942, ZN => n2937);
   U6614 : OAI222_X1 port map( A1 => n14137, A2 => n257, B1 => n7899, B2 => 
                           n14136, C1 => n14131, C2 => n265, ZN => n2942);
   U6615 : AOI221_X1 port map( B1 => n14143, B2 => n1787, C1 => n14142, C2 => 
                           n1802, A => n2979, ZN => n2974);
   U6616 : OAI222_X1 port map( A1 => n14137, A2 => n256, B1 => n7896, B2 => 
                           n14136, C1 => n14131, C2 => n264, ZN => n2979);
   U6617 : AOI221_X1 port map( B1 => n14143, B2 => n1786, C1 => n14142, C2 => 
                           n1801, A => n3016, ZN => n3011);
   U6618 : OAI222_X1 port map( A1 => n14137, A2 => n255, B1 => n7893, B2 => 
                           n14136, C1 => n14131, C2 => n263, ZN => n3016);
   U6619 : AOI221_X1 port map( B1 => n14143, B2 => n1785, C1 => n14142, C2 => 
                           n1800, A => n3053, ZN => n3048);
   U6620 : OAI222_X1 port map( A1 => n14137, A2 => n254, B1 => n7890, B2 => 
                           n14136, C1 => n14131, C2 => n262, ZN => n3053);
   U6621 : AOI221_X1 port map( B1 => n14143, B2 => n1784, C1 => n14142, C2 => 
                           n1799, A => n3090, ZN => n3085);
   U6622 : OAI222_X1 port map( A1 => n14137, A2 => n253, B1 => n7887, B2 => 
                           n14135, C1 => n14131, C2 => n261, ZN => n3090);
   U6623 : AOI221_X1 port map( B1 => n14114, B2 => n1847, C1 => n14111, C2 => 
                           n846, A => n3098, ZN => n3093);
   U6624 : OAI222_X1 port map( A1 => n301, A2 => n14108, B1 => n7640, B2 => 
                           n14105, C1 => n293, C2 => n14102, ZN => n3098);
   U6625 : AOI221_X1 port map( B1 => n13719, B2 => n8441, C1 => n13716, C2 => 
                           n8409, A => n5673, ZN => n5668);
   U6626 : OAI222_X1 port map( A1 => n2137, A2 => n13713, B1 => n6929, B2 => 
                           n13710, C1 => n1462, C2 => n13707, ZN => n5673);
   U6627 : AOI221_X1 port map( B1 => n14143, B2 => n2402, C1 => n14142, C2 => 
                           n1988, A => n3127, ZN => n3122);
   U6628 : OAI222_X1 port map( A1 => n14137, A2 => n1084, B1 => n7884, B2 => 
                           n14135, C1 => n14131, C2 => n1105, ZN => n3127);
   U6629 : AOI221_X1 port map( B1 => n14114, B2 => n2430, C1 => n14111, C2 => 
                           n848, A => n3135, ZN => n3130);
   U6630 : OAI222_X1 port map( A1 => n813, A2 => n14108, B1 => n7634, B2 => 
                           n14105, C1 => n507, C2 => n14102, ZN => n3135);
   U6631 : AOI221_X1 port map( B1 => n13719, B2 => n8440, C1 => n13716, C2 => 
                           n8408, A => n5710, ZN => n5705);
   U6632 : OAI222_X1 port map( A1 => n2136, A2 => n13713, B1 => n6953, B2 => 
                           n13710, C1 => n1461, C2 => n13707, ZN => n5710);
   U6633 : AOI221_X1 port map( B1 => n13665, B2 => n8758, C1 => n13662, C2 => 
                           n8726, A => n5718, ZN => n5713);
   U6634 : OAI222_X1 port map( A1 => n2027, A2 => n13659, B1 => n6947, B2 => 
                           n13656, C1 => n1143, C2 => n13653, ZN => n5718);
   U6635 : AOI221_X1 port map( B1 => n14113, B2 => n2429, C1 => n14110, C2 => 
                           n850, A => n3172, ZN => n3167);
   U6636 : OAI222_X1 port map( A1 => n809, A2 => n14107, B1 => n7628, B2 => 
                           n14104, C1 => n506, C2 => n14101, ZN => n3172);
   U6637 : AOI221_X1 port map( B1 => n13896, B2 => n8757, C1 => n13893, C2 => 
                           n8725, A => n4434, ZN => n4429);
   U6638 : OAI222_X1 port map( A1 => n2026, A2 => n13890, B1 => n6971, B2 => 
                           n13888, C1 => n1142, C2 => n13884, ZN => n4434);
   U6639 : AOI221_X1 port map( B1 => n13719, B2 => n8439, C1 => n13716, C2 => 
                           n8407, A => n5747, ZN => n5742);
   U6640 : OAI222_X1 port map( A1 => n2135, A2 => n13713, B1 => n6977, B2 => 
                           n13710, C1 => n1460, C2 => n13707, ZN => n5747);
   U6641 : AOI221_X1 port map( B1 => n13665, B2 => n8757, C1 => n13662, C2 => 
                           n8725, A => n5755, ZN => n5750);
   U6642 : OAI222_X1 port map( A1 => n2026, A2 => n13659, B1 => n6971, B2 => 
                           n13656, C1 => n1142, C2 => n13653, ZN => n5755);
   U6643 : AOI221_X1 port map( B1 => n14144, B2 => n2389, C1 => n14140, C2 => 
                           n1975, A => n3610, ZN => n3605);
   U6644 : OAI222_X1 port map( A1 => n14138, A2 => n1072, B1 => n7845, B2 => 
                           n14134, C1 => n14132, C2 => n1093, ZN => n3610);
   U6645 : AOI221_X1 port map( B1 => n14112, B2 => n2417, C1 => n14109, C2 => 
                           n874, A => n3618, ZN => n3613);
   U6646 : OAI222_X1 port map( A1 => n785, A2 => n14106, B1 => n7556, B2 => 
                           n14103, C1 => n494, C2 => n14100, ZN => n3618);
   U6647 : AOI221_X1 port map( B1 => n14144, B2 => n2388, C1 => n14140, C2 => 
                           n1974, A => n3647, ZN => n3642);
   U6648 : OAI222_X1 port map( A1 => n14138, A2 => n1071, B1 => n7842, B2 => 
                           n14134, C1 => n14132, C2 => n1092, ZN => n3647);
   U6649 : AOI221_X1 port map( B1 => n14112, B2 => n2416, C1 => n14109, C2 => 
                           n876, A => n3655, ZN => n3650);
   U6650 : OAI222_X1 port map( A1 => n783, A2 => n14106, B1 => n7550, B2 => 
                           n14103, C1 => n493, C2 => n14100, ZN => n3655);
   U6651 : AOI221_X1 port map( B1 => n14144, B2 => n2387, C1 => n14140, C2 => 
                           n1973, A => n3684, ZN => n3679);
   U6652 : OAI222_X1 port map( A1 => n14138, A2 => n1070, B1 => n7839, B2 => 
                           n14134, C1 => n14132, C2 => n1091, ZN => n3684);
   U6653 : AOI221_X1 port map( B1 => n14112, B2 => n2415, C1 => n14109, C2 => 
                           n878, A => n3692, ZN => n3687);
   U6654 : OAI222_X1 port map( A1 => n782, A2 => n14106, B1 => n7544, B2 => 
                           n14103, C1 => n492, C2 => n14100, ZN => n3692);
   U6655 : AOI221_X1 port map( B1 => n14144, B2 => n2386, C1 => n14140, C2 => 
                           n1972, A => n3721, ZN => n3716);
   U6656 : OAI222_X1 port map( A1 => n14139, A2 => n1069, B1 => n7836, B2 => 
                           n14134, C1 => n14133, C2 => n1090, ZN => n3721);
   U6657 : AOI221_X1 port map( B1 => n14112, B2 => n2414, C1 => n14109, C2 => 
                           n880, A => n3729, ZN => n3724);
   U6658 : OAI222_X1 port map( A1 => n781, A2 => n14106, B1 => n7538, B2 => 
                           n14103, C1 => n491, C2 => n14100, ZN => n3729);
   U6659 : AOI221_X1 port map( B1 => n14145, B2 => n2385, C1 => n14140, C2 => 
                           n1971, A => n3758, ZN => n3753);
   U6660 : OAI222_X1 port map( A1 => n14138, A2 => n1068, B1 => n7833, B2 => 
                           n14134, C1 => n14132, C2 => n1089, ZN => n3758);
   U6661 : AOI221_X1 port map( B1 => n14112, B2 => n2413, C1 => n14109, C2 => 
                           n882, A => n3766, ZN => n3761);
   U6662 : OAI222_X1 port map( A1 => n780, A2 => n14106, B1 => n7532, B2 => 
                           n14103, C1 => n490, C2 => n14100, ZN => n3766);
   U6663 : AOI221_X1 port map( B1 => n14145, B2 => n2384, C1 => n14140, C2 => 
                           n1970, A => n3795, ZN => n3790);
   U6664 : OAI222_X1 port map( A1 => n14139, A2 => n1067, B1 => n7830, B2 => 
                           n14134, C1 => n14133, C2 => n1088, ZN => n3795);
   U6665 : AOI221_X1 port map( B1 => n14112, B2 => n2412, C1 => n14109, C2 => 
                           n884, A => n3803, ZN => n3798);
   U6666 : OAI222_X1 port map( A1 => n779, A2 => n14106, B1 => n7526, B2 => 
                           n14103, C1 => n489, C2 => n14100, ZN => n3803);
   U6667 : AOI221_X1 port map( B1 => n14145, B2 => n2383, C1 => n14140, C2 => 
                           n1969, A => n3832, ZN => n3827);
   U6668 : OAI222_X1 port map( A1 => n14139, A2 => n1066, B1 => n7827, B2 => 
                           n14134, C1 => n14133, C2 => n1087, ZN => n3832);
   U6669 : AOI221_X1 port map( B1 => n14112, B2 => n2411, C1 => n14109, C2 => 
                           n886, A => n3840, ZN => n3835);
   U6670 : OAI222_X1 port map( A1 => n778, A2 => n14106, B1 => n7520, B2 => 
                           n14103, C1 => n488, C2 => n14100, ZN => n3840);
   U6671 : AOI221_X1 port map( B1 => n14145, B2 => n2382, C1 => n14140, C2 => 
                           n1968, A => n3869, ZN => n3864);
   U6672 : OAI222_X1 port map( A1 => n14139, A2 => n1065, B1 => n7824, B2 => 
                           n14134, C1 => n14133, C2 => n1707, ZN => n3869);
   U6673 : AOI221_X1 port map( B1 => n14112, B2 => n2484, C1 => n14109, C2 => 
                           n888, A => n3877, ZN => n3872);
   U6674 : OAI222_X1 port map( A1 => n776, A2 => n14106, B1 => n7514, B2 => 
                           n14103, C1 => n487, C2 => n14100, ZN => n3877);
   U6675 : AOI221_X1 port map( B1 => n14145, B2 => n2381, C1 => n14140, C2 => 
                           n1967, A => n3906, ZN => n3901);
   U6676 : OAI222_X1 port map( A1 => n14139, A2 => n1064, B1 => n7821, B2 => 
                           n14134, C1 => n14133, C2 => n1086, ZN => n3906);
   U6677 : AOI221_X1 port map( B1 => n14112, B2 => n2404, C1 => n14109, C2 => 
                           n890, A => n3914, ZN => n3909);
   U6678 : OAI222_X1 port map( A1 => n775, A2 => n14106, B1 => n7508, B2 => 
                           n14103, C1 => n486, C2 => n14100, ZN => n3914);
   U6679 : AOI221_X1 port map( B1 => n14145, B2 => n2380, C1 => n14140, C2 => 
                           n1966, A => n3943, ZN => n3938);
   U6680 : OAI222_X1 port map( A1 => n14139, A2 => n1063, B1 => n7818, B2 => 
                           n14134, C1 => n14133, C2 => n1085, ZN => n3943);
   U6681 : AOI221_X1 port map( B1 => n14112, B2 => n2403, C1 => n14109, C2 => 
                           n892, A => n3951, ZN => n3946);
   U6682 : OAI222_X1 port map( A1 => n773, A2 => n14106, B1 => n7502, B2 => 
                           n14103, C1 => n485, C2 => n14100, ZN => n3951);
   U6683 : AOI221_X1 port map( B1 => n14112, B2 => n1855, C1 => n14109, C2 => 
                           n894, A => n5273, ZN => n5268);
   U6684 : OAI222_X1 port map( A1 => n772, A2 => n14106, B1 => n7496, B2 => 
                           n14103, C1 => n484, C2 => n14100, ZN => n5273);
   U6685 : AOI221_X1 port map( B1 => n14145, B2 => n2379, C1 => n14140, C2 => 
                           n1965, A => n5265, ZN => n5260);
   U6686 : OAI222_X1 port map( A1 => n14139, A2 => n1062, B1 => n14134, B2 => 
                           n1061, C1 => n14133, C2 => n1607, ZN => n5265);
   U6687 : AOI221_X1 port map( B1 => n8672, B2 => n13883, C1 => n8640, C2 => 
                           n13878, A => n5228, ZN => n5220);
   U6688 : OAI22_X1 port map( A1 => n13877, A2 => n1265, B1 => n13874, B2 => 
                           n1241, ZN => n5228);
   U6689 : AOI221_X1 port map( B1 => n8703, B2 => n13883, C1 => n8671, C2 => 
                           n13878, A => n4061, ZN => n4038);
   U6690 : OAI22_X1 port map( A1 => n13877, A2 => n131, B1 => n13874, B2 => 
                           n123, ZN => n4061);
   U6691 : AOI221_X1 port map( B1 => n14738, B2 => n2338, C1 => n14741, C2 => 
                           n774, A => n4797, ZN => n4790);
   U6692 : OAI22_X1 port map( A1 => n1523, A2 => n13870, B1 => n1547, B2 => 
                           n13868, ZN => n4797);
   U6693 : AOI221_X1 port map( B1 => n14097, B2 => n8099, C1 => n14094, C2 => 
                           n8131, A => n6603, ZN => n6595);
   U6694 : OAI22_X1 port map( A1 => n6745, A2 => n14091, B1 => n6744, B2 => 
                           n14088, ZN => n6603);
   U6695 : AOI221_X1 port map( B1 => n14099, B2 => n8098, C1 => n14096, C2 => 
                           n8130, A => n2875, ZN => n2859);
   U6696 : OAI22_X1 port map( A1 => n411, A2 => n14093, B1 => n6768, B2 => 
                           n14090, ZN => n2875);
   U6697 : AOI221_X1 port map( B1 => n14099, B2 => n8097, C1 => n14096, C2 => 
                           n8129, A => n2914, ZN => n2907);
   U6698 : OAI22_X1 port map( A1 => n410, A2 => n14093, B1 => n6792, B2 => 
                           n14090, ZN => n2914);
   U6699 : AOI221_X1 port map( B1 => n14099, B2 => n8096, C1 => n14096, C2 => 
                           n8128, A => n2951, ZN => n2944);
   U6700 : OAI22_X1 port map( A1 => n409, A2 => n14093, B1 => n6816, B2 => 
                           n14090, ZN => n2951);
   U6701 : AOI221_X1 port map( B1 => n14099, B2 => n8095, C1 => n14096, C2 => 
                           n8127, A => n2988, ZN => n2981);
   U6702 : OAI22_X1 port map( A1 => n408, A2 => n14093, B1 => n6840, B2 => 
                           n14090, ZN => n2988);
   U6703 : AOI221_X1 port map( B1 => n14099, B2 => n8094, C1 => n14096, C2 => 
                           n8126, A => n3025, ZN => n3018);
   U6704 : OAI22_X1 port map( A1 => n407, A2 => n14093, B1 => n6864, B2 => 
                           n14090, ZN => n3025);
   U6705 : AOI221_X1 port map( B1 => n14099, B2 => n8093, C1 => n14096, C2 => 
                           n8125, A => n3062, ZN => n3055);
   U6706 : OAI22_X1 port map( A1 => n406, A2 => n14093, B1 => n6888, B2 => 
                           n14090, ZN => n3062);
   U6707 : AOI221_X1 port map( B1 => n14099, B2 => n8092, C1 => n14096, C2 => 
                           n8124, A => n3099, ZN => n3092);
   U6708 : OAI22_X1 port map( A1 => n405, A2 => n14093, B1 => n6912, B2 => 
                           n14090, ZN => n3099);
   U6709 : AOI221_X1 port map( B1 => n14099, B2 => n8091, C1 => n14096, C2 => 
                           n8123, A => n3136, ZN => n3129);
   U6710 : OAI22_X1 port map( A1 => n1706, A2 => n14093, B1 => n6936, B2 => 
                           n14090, ZN => n3136);
   U6711 : AOI221_X1 port map( B1 => n14098, B2 => n8089, C1 => n14095, C2 => 
                           n8121, A => n3210, ZN => n3203);
   U6712 : OAI22_X1 port map( A1 => n1704, A2 => n14092, B1 => n6984, B2 => 
                           n14089, ZN => n3210);
   U6713 : AOI221_X1 port map( B1 => n14098, B2 => n8084, C1 => n14095, C2 => 
                           n8116, A => n3397, ZN => n3390);
   U6714 : OAI22_X1 port map( A1 => n1699, A2 => n14092, B1 => n1693, B2 => 
                           n14089, ZN => n3397);
   U6715 : AOI221_X1 port map( B1 => n13881, B2 => n8697, C1 => n13878, C2 => 
                           n8665, A => n4287, ZN => n4280);
   U6716 : OAI22_X1 port map( A1 => n125, A2 => n13875, B1 => n117, B2 => 
                           n13872, ZN => n4287);
   U6717 : AOI221_X1 port map( B1 => n13882, B2 => n8683, C1 => n13879, C2 => 
                           n8651, A => n4805, ZN => n4798);
   U6718 : OAI22_X1 port map( A1 => n1276, A2 => n13876, B1 => n786, B2 => 
                           n13873, ZN => n4805);
   U6719 : AOI221_X1 port map( B1 => n13882, B2 => n8682, C1 => n13879, C2 => 
                           n8650, A => n4842, ZN => n4835);
   U6720 : OAI22_X1 port map( A1 => n1275, A2 => n13876, B1 => n1251, B2 => 
                           n13873, ZN => n4842);
   U6721 : AOI221_X1 port map( B1 => n13882, B2 => n8681, C1 => n13879, C2 => 
                           n8649, A => n4879, ZN => n4872);
   U6722 : OAI22_X1 port map( A1 => n1274, A2 => n13876, B1 => n1250, B2 => 
                           n13873, ZN => n4879);
   U6723 : AOI221_X1 port map( B1 => n13882, B2 => n8680, C1 => n13879, C2 => 
                           n8648, A => n4916, ZN => n4909);
   U6724 : OAI22_X1 port map( A1 => n1273, A2 => n13876, B1 => n1249, B2 => 
                           n13873, ZN => n4916);
   U6725 : AOI221_X1 port map( B1 => n13882, B2 => n8679, C1 => n13880, C2 => 
                           n8647, A => n4953, ZN => n4946);
   U6726 : OAI22_X1 port map( A1 => n1272, A2 => n13876, B1 => n1248, B2 => 
                           n13873, ZN => n4953);
   U6727 : AOI221_X1 port map( B1 => n13882, B2 => n8685, C1 => n13879, C2 => 
                           n8653, A => n4731, ZN => n4724);
   U6728 : OAI22_X1 port map( A1 => n1278, A2 => n13876, B1 => n1254, B2 => 
                           n13873, ZN => n4731);
   U6729 : AOI221_X1 port map( B1 => n13882, B2 => n8684, C1 => n13879, C2 => 
                           n8652, A => n4768, ZN => n4761);
   U6730 : OAI22_X1 port map( A1 => n1277, A2 => n13876, B1 => n1253, B2 => 
                           n13873, ZN => n4768);
   U6731 : AOI221_X1 port map( B1 => n13650, B2 => n8653, C1 => n13647, C2 => 
                           n8685, A => n6052, ZN => n6045);
   U6732 : OAI22_X1 port map( A1 => n1254, A2 => n13644, B1 => n1278, B2 => 
                           n13641, ZN => n6052);
   U6733 : AOI221_X1 port map( B1 => n13650, B2 => n8652, C1 => n13647, C2 => 
                           n8684, A => n6089, ZN => n6082);
   U6734 : OAI22_X1 port map( A1 => n1253, A2 => n13644, B1 => n1277, B2 => 
                           n13641, ZN => n6089);
   U6735 : AOI221_X1 port map( B1 => n13649, B2 => n8640, C1 => n13646, C2 => 
                           n8672, A => n6549, ZN => n6541);
   U6736 : OAI22_X1 port map( A1 => n1241, A2 => n13643, B1 => n1265, B2 => 
                           n13640, ZN => n6549);
   U6737 : AOI221_X1 port map( B1 => n13651, B2 => n8671, C1 => n13648, C2 => 
                           n8703, A => n5384, ZN => n5361);
   U6738 : OAI22_X1 port map( A1 => n123, A2 => n13645, B1 => n131, B2 => 
                           n13642, ZN => n5384);
   U6739 : AOI221_X1 port map( B1 => n13881, B2 => n8702, C1 => n13878, C2 => 
                           n8670, A => n4102, ZN => n4095);
   U6740 : OAI22_X1 port map( A1 => n130, A2 => n13875, B1 => n122, B2 => 
                           n13872, ZN => n4102);
   U6741 : AOI221_X1 port map( B1 => n13881, B2 => n8701, C1 => n13878, C2 => 
                           n8669, A => n4139, ZN => n4132);
   U6742 : OAI22_X1 port map( A1 => n129, A2 => n13875, B1 => n121, B2 => 
                           n13872, ZN => n4139);
   U6743 : AOI221_X1 port map( B1 => n13881, B2 => n8700, C1 => n13878, C2 => 
                           n8668, A => n4176, ZN => n4169);
   U6744 : OAI22_X1 port map( A1 => n128, A2 => n13875, B1 => n120, B2 => 
                           n13872, ZN => n4176);
   U6745 : AOI221_X1 port map( B1 => n13881, B2 => n8699, C1 => n13878, C2 => 
                           n8667, A => n4213, ZN => n4206);
   U6746 : OAI22_X1 port map( A1 => n127, A2 => n13875, B1 => n119, B2 => 
                           n13872, ZN => n4213);
   U6747 : AOI221_X1 port map( B1 => n14098, B2 => n8090, C1 => n14095, C2 => 
                           n8122, A => n3173, ZN => n3166);
   U6748 : OAI22_X1 port map( A1 => n1705, A2 => n14092, B1 => n6960, B2 => 
                           n14089, ZN => n3173);
   U6749 : AOI221_X1 port map( B1 => n14098, B2 => n8088, C1 => n14095, C2 => 
                           n8120, A => n3247, ZN => n3240);
   U6750 : OAI22_X1 port map( A1 => n1703, A2 => n14092, B1 => n7008, B2 => 
                           n14089, ZN => n3247);
   U6751 : AOI221_X1 port map( B1 => n14098, B2 => n8087, C1 => n14095, C2 => 
                           n8119, A => n3284, ZN => n3277);
   U6752 : OAI22_X1 port map( A1 => n1702, A2 => n14092, B1 => n1696, B2 => 
                           n14089, ZN => n3284);
   U6753 : AOI221_X1 port map( B1 => n14098, B2 => n8086, C1 => n14095, C2 => 
                           n8118, A => n3323, ZN => n3316);
   U6754 : OAI22_X1 port map( A1 => n1701, A2 => n14092, B1 => n1695, B2 => 
                           n14089, ZN => n3323);
   U6755 : AOI221_X1 port map( B1 => n14098, B2 => n8085, C1 => n14095, C2 => 
                           n8117, A => n3360, ZN => n3353);
   U6756 : OAI22_X1 port map( A1 => n1700, A2 => n14092, B1 => n1694, B2 => 
                           n14089, ZN => n3360);
   U6757 : AOI221_X1 port map( B1 => n14098, B2 => n8083, C1 => n14095, C2 => 
                           n8115, A => n3434, ZN => n3427);
   U6758 : OAI22_X1 port map( A1 => n1698, A2 => n14092, B1 => n1692, B2 => 
                           n14089, ZN => n3434);
   U6759 : AOI221_X1 port map( B1 => n14098, B2 => n8082, C1 => n14095, C2 => 
                           n8114, A => n3471, ZN => n3464);
   U6760 : OAI22_X1 port map( A1 => n1697, A2 => n14092, B1 => n7152, B2 => 
                           n14089, ZN => n3471);
   U6761 : AOI221_X1 port map( B1 => n14098, B2 => n8081, C1 => n14095, C2 => 
                           n8113, A => n3508, ZN => n3501);
   U6762 : OAI22_X1 port map( A1 => n7177, A2 => n14092, B1 => n7176, B2 => 
                           n14089, ZN => n3508);
   U6763 : AOI221_X1 port map( B1 => n14098, B2 => n8079, C1 => n14095, C2 => 
                           n8111, A => n3582, ZN => n3575);
   U6764 : OAI22_X1 port map( A1 => n2482, A2 => n14092, B1 => n2480, B2 => 
                           n14089, ZN => n3582);
   U6765 : AOI221_X1 port map( B1 => n14097, B2 => n8078, C1 => n14094, C2 => 
                           n8110, A => n3619, ZN => n3612);
   U6766 : OAI22_X1 port map( A1 => n7249, A2 => n14091, B1 => n7248, B2 => 
                           n14088, ZN => n3619);
   U6767 : AOI221_X1 port map( B1 => n14097, B2 => n8077, C1 => n14094, C2 => 
                           n8109, A => n3656, ZN => n3649);
   U6768 : OAI22_X1 port map( A1 => n7273, A2 => n14091, B1 => n7272, B2 => 
                           n14088, ZN => n3656);
   U6769 : AOI221_X1 port map( B1 => n14097, B2 => n8076, C1 => n14094, C2 => 
                           n8108, A => n3693, ZN => n3686);
   U6770 : OAI22_X1 port map( A1 => n7297, A2 => n14091, B1 => n7296, B2 => 
                           n14088, ZN => n3693);
   U6771 : AOI221_X1 port map( B1 => n14097, B2 => n8075, C1 => n14094, C2 => 
                           n8107, A => n3730, ZN => n3723);
   U6772 : OAI22_X1 port map( A1 => n7321, A2 => n14091, B1 => n7320, B2 => 
                           n14088, ZN => n3730);
   U6773 : AOI221_X1 port map( B1 => n14097, B2 => n8074, C1 => n14094, C2 => 
                           n8106, A => n3767, ZN => n3760);
   U6774 : OAI22_X1 port map( A1 => n7345, A2 => n14091, B1 => n7344, B2 => 
                           n14088, ZN => n3767);
   U6775 : AOI221_X1 port map( B1 => n14097, B2 => n8073, C1 => n14094, C2 => 
                           n8105, A => n3804, ZN => n3797);
   U6776 : OAI22_X1 port map( A1 => n7369, A2 => n14091, B1 => n7368, B2 => 
                           n14088, ZN => n3804);
   U6777 : AOI221_X1 port map( B1 => n14097, B2 => n8072, C1 => n14094, C2 => 
                           n8104, A => n3841, ZN => n3834);
   U6778 : OAI22_X1 port map( A1 => n7393, A2 => n14091, B1 => n7392, B2 => 
                           n14088, ZN => n3841);
   U6779 : AOI221_X1 port map( B1 => n14097, B2 => n8071, C1 => n14094, C2 => 
                           n8103, A => n3878, ZN => n3871);
   U6780 : OAI22_X1 port map( A1 => n7417, A2 => n14091, B1 => n7416, B2 => 
                           n14088, ZN => n3878);
   U6781 : AOI221_X1 port map( B1 => n14097, B2 => n8070, C1 => n14094, C2 => 
                           n8102, A => n3915, ZN => n3908);
   U6782 : OAI22_X1 port map( A1 => n7441, A2 => n14091, B1 => n7440, B2 => 
                           n14088, ZN => n3915);
   U6783 : AOI221_X1 port map( B1 => n14097, B2 => n8069, C1 => n14094, C2 => 
                           n8101, A => n3952, ZN => n3945);
   U6784 : OAI22_X1 port map( A1 => n7465, A2 => n14091, B1 => n7464, B2 => 
                           n14088, ZN => n3952);
   U6785 : AOI221_X1 port map( B1 => n14097, B2 => n8068, C1 => n14094, C2 => 
                           n8100, A => n5274, ZN => n5267);
   U6786 : OAI22_X1 port map( A1 => n7489, A2 => n14091, B1 => n7488, B2 => 
                           n14088, ZN => n5274);
   U6787 : AOI221_X1 port map( B1 => n13881, B2 => n8698, C1 => n13878, C2 => 
                           n8666, A => n4250, ZN => n4243);
   U6788 : OAI22_X1 port map( A1 => n126, A2 => n13875, B1 => n118, B2 => 
                           n13872, ZN => n4250);
   U6789 : AOI221_X1 port map( B1 => n13881, B2 => n8696, C1 => n13878, C2 => 
                           n8664, A => n4324, ZN => n4317);
   U6790 : OAI22_X1 port map( A1 => n124, A2 => n13875, B1 => n116, B2 => 
                           n13872, ZN => n4324);
   U6791 : AOI221_X1 port map( B1 => n13651, B2 => n8664, C1 => n13648, C2 => 
                           n8696, A => n5645, ZN => n5638);
   U6792 : OAI22_X1 port map( A1 => n116, A2 => n13645, B1 => n124, B2 => 
                           n13642, ZN => n5645);
   U6793 : AOI221_X1 port map( B1 => n13882, B2 => n8695, C1 => n13879, C2 => 
                           n8663, A => n4361, ZN => n4354);
   U6794 : OAI22_X1 port map( A1 => n1288, A2 => n13876, B1 => n1264, B2 => 
                           n13873, ZN => n4361);
   U6795 : AOI221_X1 port map( B1 => n13650, B2 => n8663, C1 => n13647, C2 => 
                           n8695, A => n5682, ZN => n5675);
   U6796 : OAI22_X1 port map( A1 => n1264, A2 => n13644, B1 => n1288, B2 => 
                           n13641, ZN => n5682);
   U6797 : AOI221_X1 port map( B1 => n13881, B2 => n8694, C1 => n13878, C2 => 
                           n8662, A => n4398, ZN => n4391);
   U6798 : OAI22_X1 port map( A1 => n1287, A2 => n13875, B1 => n1263, B2 => 
                           n13872, ZN => n4398);
   U6799 : AOI221_X1 port map( B1 => n13650, B2 => n8662, C1 => n13647, C2 => 
                           n8694, A => n5719, ZN => n5712);
   U6800 : OAI22_X1 port map( A1 => n1263, A2 => n13644, B1 => n1287, B2 => 
                           n13641, ZN => n5719);
   U6801 : AOI221_X1 port map( B1 => n13881, B2 => n8693, C1 => n13878, C2 => 
                           n8661, A => n4435, ZN => n4428);
   U6802 : OAI22_X1 port map( A1 => n1286, A2 => n13875, B1 => n1262, B2 => 
                           n13872, ZN => n4435);
   U6803 : AOI221_X1 port map( B1 => n13650, B2 => n8661, C1 => n13647, C2 => 
                           n8693, A => n5756, ZN => n5749);
   U6804 : OAI22_X1 port map( A1 => n1262, A2 => n13644, B1 => n1286, B2 => 
                           n13641, ZN => n5756);
   U6805 : AOI221_X1 port map( B1 => n13881, B2 => n8692, C1 => n13878, C2 => 
                           n8660, A => n4472, ZN => n4465);
   U6806 : OAI22_X1 port map( A1 => n1285, A2 => n13875, B1 => n1261, B2 => 
                           n13872, ZN => n4472);
   U6807 : AOI221_X1 port map( B1 => n13650, B2 => n8660, C1 => n13647, C2 => 
                           n8692, A => n5793, ZN => n5786);
   U6808 : OAI22_X1 port map( A1 => n1261, A2 => n13644, B1 => n1285, B2 => 
                           n13641, ZN => n5793);
   U6809 : AOI221_X1 port map( B1 => n13881, B2 => n8691, C1 => n13879, C2 => 
                           n8659, A => n4509, ZN => n4502);
   U6810 : OAI22_X1 port map( A1 => n1284, A2 => n13875, B1 => n1260, B2 => 
                           n13872, ZN => n4509);
   U6811 : AOI221_X1 port map( B1 => n13650, B2 => n8659, C1 => n13647, C2 => 
                           n8691, A => n5830, ZN => n5823);
   U6812 : OAI22_X1 port map( A1 => n1260, A2 => n13644, B1 => n1284, B2 => 
                           n13641, ZN => n5830);
   U6813 : AOI221_X1 port map( B1 => n13881, B2 => n8690, C1 => n13879, C2 => 
                           n8658, A => n4546, ZN => n4539);
   U6814 : OAI22_X1 port map( A1 => n1283, A2 => n13875, B1 => n1259, B2 => 
                           n13872, ZN => n4546);
   U6815 : AOI221_X1 port map( B1 => n13650, B2 => n8658, C1 => n13647, C2 => 
                           n8690, A => n5867, ZN => n5860);
   U6816 : OAI22_X1 port map( A1 => n1259, A2 => n13644, B1 => n1283, B2 => 
                           n13641, ZN => n5867);
   U6817 : AOI221_X1 port map( B1 => n13882, B2 => n8689, C1 => n13879, C2 => 
                           n8657, A => n4583, ZN => n4576);
   U6818 : OAI22_X1 port map( A1 => n1282, A2 => n13876, B1 => n1258, B2 => 
                           n13873, ZN => n4583);
   U6819 : AOI221_X1 port map( B1 => n13650, B2 => n8657, C1 => n13647, C2 => 
                           n8689, A => n5904, ZN => n5897);
   U6820 : OAI22_X1 port map( A1 => n1258, A2 => n13644, B1 => n1282, B2 => 
                           n13641, ZN => n5904);
   U6821 : AOI221_X1 port map( B1 => n13882, B2 => n8688, C1 => n13879, C2 => 
                           n8656, A => n4620, ZN => n4613);
   U6822 : OAI22_X1 port map( A1 => n1281, A2 => n13876, B1 => n1257, B2 => 
                           n13873, ZN => n4620);
   U6823 : AOI221_X1 port map( B1 => n13650, B2 => n8656, C1 => n13647, C2 => 
                           n8688, A => n5941, ZN => n5934);
   U6824 : OAI22_X1 port map( A1 => n1257, A2 => n13644, B1 => n1281, B2 => 
                           n13641, ZN => n5941);
   U6825 : AOI221_X1 port map( B1 => n13882, B2 => n8687, C1 => n13879, C2 => 
                           n8655, A => n4657, ZN => n4650);
   U6826 : OAI22_X1 port map( A1 => n1280, A2 => n13876, B1 => n1256, B2 => 
                           n13873, ZN => n4657);
   U6827 : AOI221_X1 port map( B1 => n13650, B2 => n8655, C1 => n13647, C2 => 
                           n8687, A => n5978, ZN => n5971);
   U6828 : OAI22_X1 port map( A1 => n1256, A2 => n13644, B1 => n1280, B2 => 
                           n13641, ZN => n5978);
   U6829 : AOI221_X1 port map( B1 => n13882, B2 => n8686, C1 => n13879, C2 => 
                           n8654, A => n4694, ZN => n4687);
   U6830 : OAI22_X1 port map( A1 => n1279, A2 => n13876, B1 => n1255, B2 => 
                           n13873, ZN => n4694);
   U6831 : AOI221_X1 port map( B1 => n13650, B2 => n8654, C1 => n13647, C2 => 
                           n8686, A => n6015, ZN => n6008);
   U6832 : OAI22_X1 port map( A1 => n1255, A2 => n13644, B1 => n1279, B2 => 
                           n13641, ZN => n6015);
   U6833 : AOI221_X1 port map( B1 => n8322, B2 => n13220, C1 => n8354, C2 => 
                           n13871, A => n5219, ZN => n5210);
   U6834 : OAI22_X1 port map( A1 => n4036, A2 => n1511, B1 => n7688, B2 => 
                           n4037, ZN => n5219);
   U6835 : AOI221_X1 port map( B1 => n13703, B2 => n2338, C1 => n13700, C2 => 
                           n774, A => n6118, ZN => n6111);
   U6836 : OAI22_X1 port map( A1 => n1523, A2 => n13697, B1 => n1547, B2 => 
                           n13694, ZN => n6118);
   U6837 : AOI221_X1 port map( B1 => n8353, B2 => n13220, C1 => n8385, C2 => 
                           n13871, A => n4035, ZN => n4014);
   U6838 : OAI22_X1 port map( A1 => n4036, A2 => n212, B1 => n7812, B2 => n4037
                           , ZN => n4035);
   U6839 : AOI221_X1 port map( B1 => n13705, B2 => n1781, C1 => n13702, C2 => 
                           n830, A => n5358, ZN => n5335);
   U6840 : OAI22_X1 port map( A1 => n220, A2 => n13699, B1 => n228, B2 => 
                           n13696, ZN => n5358);
   U6841 : BUF_X1 port map( A => n7627, Z => n14761);
   U6842 : BUF_X1 port map( A => n7629, Z => n14755);
   U6843 : BUF_X1 port map( A => n7596, Z => n14887);
   U6844 : BUF_X1 port map( A => n7597, Z => n14881);
   U6845 : BUF_X1 port map( A => n7599, Z => n14875);
   U6846 : BUF_X1 port map( A => n7601, Z => n14869);
   U6847 : BUF_X1 port map( A => n7602, Z => n14863);
   U6848 : BUF_X1 port map( A => n7603, Z => n14857);
   U6849 : BUF_X1 port map( A => n7605, Z => n14851);
   U6850 : BUF_X1 port map( A => n7607, Z => n14845);
   U6851 : BUF_X1 port map( A => n7608, Z => n14839);
   U6852 : BUF_X1 port map( A => n7609, Z => n14833);
   U6853 : BUF_X1 port map( A => n7611, Z => n14827);
   U6854 : BUF_X1 port map( A => n7613, Z => n14821);
   U6855 : BUF_X1 port map( A => n7614, Z => n14815);
   U6856 : BUF_X1 port map( A => n7615, Z => n14809);
   U6857 : BUF_X1 port map( A => n7617, Z => n14803);
   U6858 : BUF_X1 port map( A => n7619, Z => n14797);
   U6859 : BUF_X1 port map( A => n7620, Z => n14791);
   U6860 : BUF_X1 port map( A => n7621, Z => n14785);
   U6861 : BUF_X1 port map( A => n7623, Z => n14779);
   U6862 : BUF_X1 port map( A => n7625, Z => n14773);
   U6863 : BUF_X1 port map( A => n7631, Z => n14749);
   U6864 : BUF_X1 port map( A => n7584, Z => n14935);
   U6865 : BUF_X1 port map( A => n7585, Z => n14929);
   U6866 : BUF_X1 port map( A => n7587, Z => n14923);
   U6867 : BUF_X1 port map( A => n7589, Z => n14917);
   U6868 : BUF_X1 port map( A => n7590, Z => n14911);
   U6869 : BUF_X1 port map( A => n7591, Z => n14905);
   U6870 : BUF_X1 port map( A => n7593, Z => n14899);
   U6871 : BUF_X1 port map( A => n7595, Z => n14893);
   U6872 : BUF_X1 port map( A => n7626, Z => n14767);
   U6873 : BUF_X1 port map( A => n7626, Z => n14771);
   U6874 : BUF_X1 port map( A => n7596, Z => n14891);
   U6875 : BUF_X1 port map( A => n7597, Z => n14885);
   U6876 : BUF_X1 port map( A => n7599, Z => n14879);
   U6877 : BUF_X1 port map( A => n7601, Z => n14873);
   U6878 : BUF_X1 port map( A => n7602, Z => n14867);
   U6879 : BUF_X1 port map( A => n7603, Z => n14861);
   U6880 : BUF_X1 port map( A => n7605, Z => n14855);
   U6881 : BUF_X1 port map( A => n7607, Z => n14849);
   U6882 : BUF_X1 port map( A => n7608, Z => n14843);
   U6883 : BUF_X1 port map( A => n7609, Z => n14837);
   U6884 : BUF_X1 port map( A => n7611, Z => n14831);
   U6885 : BUF_X1 port map( A => n7613, Z => n14825);
   U6886 : BUF_X1 port map( A => n7614, Z => n14819);
   U6887 : BUF_X1 port map( A => n7615, Z => n14813);
   U6888 : BUF_X1 port map( A => n7617, Z => n14807);
   U6889 : BUF_X1 port map( A => n7619, Z => n14801);
   U6890 : BUF_X1 port map( A => n7620, Z => n14795);
   U6891 : BUF_X1 port map( A => n7621, Z => n14789);
   U6892 : BUF_X1 port map( A => n7623, Z => n14783);
   U6893 : BUF_X1 port map( A => n7625, Z => n14777);
   U6894 : BUF_X1 port map( A => n7627, Z => n14765);
   U6895 : BUF_X1 port map( A => n7629, Z => n14759);
   U6896 : BUF_X1 port map( A => n7631, Z => n14753);
   U6897 : BUF_X1 port map( A => n7611, Z => n14830);
   U6898 : BUF_X1 port map( A => n7613, Z => n14824);
   U6899 : BUF_X1 port map( A => n7614, Z => n14818);
   U6900 : BUF_X1 port map( A => n7615, Z => n14812);
   U6901 : BUF_X1 port map( A => n7617, Z => n14806);
   U6902 : BUF_X1 port map( A => n7619, Z => n14800);
   U6903 : BUF_X1 port map( A => n7620, Z => n14794);
   U6904 : BUF_X1 port map( A => n7621, Z => n14788);
   U6905 : BUF_X1 port map( A => n7623, Z => n14782);
   U6906 : BUF_X1 port map( A => n7625, Z => n14776);
   U6907 : BUF_X1 port map( A => n7626, Z => n14770);
   U6908 : BUF_X1 port map( A => n7596, Z => n14890);
   U6909 : BUF_X1 port map( A => n7597, Z => n14884);
   U6910 : BUF_X1 port map( A => n7599, Z => n14878);
   U6911 : BUF_X1 port map( A => n7601, Z => n14872);
   U6912 : BUF_X1 port map( A => n7602, Z => n14866);
   U6913 : BUF_X1 port map( A => n7603, Z => n14860);
   U6914 : BUF_X1 port map( A => n7605, Z => n14854);
   U6915 : BUF_X1 port map( A => n7607, Z => n14848);
   U6916 : BUF_X1 port map( A => n7608, Z => n14842);
   U6917 : BUF_X1 port map( A => n7609, Z => n14836);
   U6918 : BUF_X1 port map( A => n7596, Z => n14892);
   U6919 : BUF_X1 port map( A => n7597, Z => n14886);
   U6920 : BUF_X1 port map( A => n7599, Z => n14880);
   U6921 : BUF_X1 port map( A => n7601, Z => n14874);
   U6922 : BUF_X1 port map( A => n7602, Z => n14868);
   U6923 : BUF_X1 port map( A => n7603, Z => n14862);
   U6924 : BUF_X1 port map( A => n7605, Z => n14856);
   U6925 : BUF_X1 port map( A => n7607, Z => n14850);
   U6926 : BUF_X1 port map( A => n7608, Z => n14844);
   U6927 : BUF_X1 port map( A => n7609, Z => n14838);
   U6928 : BUF_X1 port map( A => n7611, Z => n14832);
   U6929 : BUF_X1 port map( A => n7613, Z => n14826);
   U6930 : BUF_X1 port map( A => n7614, Z => n14820);
   U6931 : BUF_X1 port map( A => n7615, Z => n14814);
   U6932 : BUF_X1 port map( A => n7617, Z => n14808);
   U6933 : BUF_X1 port map( A => n7619, Z => n14802);
   U6934 : BUF_X1 port map( A => n7620, Z => n14796);
   U6935 : BUF_X1 port map( A => n7621, Z => n14790);
   U6936 : BUF_X1 port map( A => n7623, Z => n14784);
   U6937 : BUF_X1 port map( A => n7625, Z => n14778);
   U6938 : BUF_X1 port map( A => n7626, Z => n14772);
   U6939 : BUF_X1 port map( A => n7627, Z => n14766);
   U6940 : BUF_X1 port map( A => n7629, Z => n14760);
   U6941 : BUF_X1 port map( A => n7631, Z => n14754);
   U6942 : BUF_X1 port map( A => n7596, Z => n14889);
   U6943 : BUF_X1 port map( A => n7597, Z => n14883);
   U6944 : BUF_X1 port map( A => n7599, Z => n14877);
   U6945 : BUF_X1 port map( A => n7601, Z => n14871);
   U6946 : BUF_X1 port map( A => n7602, Z => n14865);
   U6947 : BUF_X1 port map( A => n7603, Z => n14859);
   U6948 : BUF_X1 port map( A => n7605, Z => n14853);
   U6949 : BUF_X1 port map( A => n7607, Z => n14847);
   U6950 : BUF_X1 port map( A => n7608, Z => n14841);
   U6951 : BUF_X1 port map( A => n7609, Z => n14835);
   U6952 : BUF_X1 port map( A => n7611, Z => n14829);
   U6953 : BUF_X1 port map( A => n7613, Z => n14823);
   U6954 : BUF_X1 port map( A => n7614, Z => n14817);
   U6955 : BUF_X1 port map( A => n7615, Z => n14811);
   U6956 : BUF_X1 port map( A => n7617, Z => n14805);
   U6957 : BUF_X1 port map( A => n7619, Z => n14799);
   U6958 : BUF_X1 port map( A => n7620, Z => n14793);
   U6959 : BUF_X1 port map( A => n7621, Z => n14787);
   U6960 : BUF_X1 port map( A => n7623, Z => n14781);
   U6961 : BUF_X1 port map( A => n7625, Z => n14775);
   U6962 : BUF_X1 port map( A => n7626, Z => n14769);
   U6963 : BUF_X1 port map( A => n7631, Z => n14751);
   U6964 : BUF_X1 port map( A => n7627, Z => n14763);
   U6965 : BUF_X1 port map( A => n7629, Z => n14757);
   U6966 : BUF_X1 port map( A => n7627, Z => n14764);
   U6967 : BUF_X1 port map( A => n7629, Z => n14758);
   U6968 : BUF_X1 port map( A => n7631, Z => n14752);
   U6969 : BUF_X1 port map( A => n7626, Z => n14768);
   U6970 : BUF_X1 port map( A => n7596, Z => n14888);
   U6971 : BUF_X1 port map( A => n7597, Z => n14882);
   U6972 : BUF_X1 port map( A => n7599, Z => n14876);
   U6973 : BUF_X1 port map( A => n7601, Z => n14870);
   U6974 : BUF_X1 port map( A => n7602, Z => n14864);
   U6975 : BUF_X1 port map( A => n7603, Z => n14858);
   U6976 : BUF_X1 port map( A => n7605, Z => n14852);
   U6977 : BUF_X1 port map( A => n7607, Z => n14846);
   U6978 : BUF_X1 port map( A => n7608, Z => n14840);
   U6979 : BUF_X1 port map( A => n7609, Z => n14834);
   U6980 : BUF_X1 port map( A => n7611, Z => n14828);
   U6981 : BUF_X1 port map( A => n7613, Z => n14822);
   U6982 : BUF_X1 port map( A => n7614, Z => n14816);
   U6983 : BUF_X1 port map( A => n7615, Z => n14810);
   U6984 : BUF_X1 port map( A => n7617, Z => n14804);
   U6985 : BUF_X1 port map( A => n7619, Z => n14798);
   U6986 : BUF_X1 port map( A => n7620, Z => n14792);
   U6987 : BUF_X1 port map( A => n7621, Z => n14786);
   U6988 : BUF_X1 port map( A => n7623, Z => n14780);
   U6989 : BUF_X1 port map( A => n7625, Z => n14774);
   U6990 : BUF_X1 port map( A => n7627, Z => n14762);
   U6991 : BUF_X1 port map( A => n7629, Z => n14756);
   U6992 : BUF_X1 port map( A => n7631, Z => n14750);
   U6993 : BUF_X1 port map( A => n7584, Z => n14936);
   U6994 : BUF_X1 port map( A => n7585, Z => n14930);
   U6995 : BUF_X1 port map( A => n7587, Z => n14924);
   U6996 : BUF_X1 port map( A => n7589, Z => n14918);
   U6997 : BUF_X1 port map( A => n7590, Z => n14912);
   U6998 : BUF_X1 port map( A => n7591, Z => n14906);
   U6999 : BUF_X1 port map( A => n7593, Z => n14900);
   U7000 : BUF_X1 port map( A => n7595, Z => n14894);
   U7001 : BUF_X1 port map( A => n7584, Z => n14940);
   U7002 : BUF_X1 port map( A => n7585, Z => n14934);
   U7003 : BUF_X1 port map( A => n7587, Z => n14928);
   U7004 : BUF_X1 port map( A => n7589, Z => n14922);
   U7005 : BUF_X1 port map( A => n7590, Z => n14916);
   U7006 : BUF_X1 port map( A => n7591, Z => n14910);
   U7007 : BUF_X1 port map( A => n7593, Z => n14904);
   U7008 : BUF_X1 port map( A => n7595, Z => n14898);
   U7009 : BUF_X1 port map( A => n7584, Z => n14939);
   U7010 : BUF_X1 port map( A => n7585, Z => n14933);
   U7011 : BUF_X1 port map( A => n7587, Z => n14927);
   U7012 : BUF_X1 port map( A => n7589, Z => n14921);
   U7013 : BUF_X1 port map( A => n7590, Z => n14915);
   U7014 : BUF_X1 port map( A => n7591, Z => n14909);
   U7015 : BUF_X1 port map( A => n7593, Z => n14903);
   U7016 : BUF_X1 port map( A => n7595, Z => n14897);
   U7017 : BUF_X1 port map( A => n7584, Z => n14938);
   U7018 : BUF_X1 port map( A => n7585, Z => n14932);
   U7019 : BUF_X1 port map( A => n7587, Z => n14926);
   U7020 : BUF_X1 port map( A => n7589, Z => n14920);
   U7021 : BUF_X1 port map( A => n7590, Z => n14914);
   U7022 : BUF_X1 port map( A => n7591, Z => n14908);
   U7023 : BUF_X1 port map( A => n7593, Z => n14902);
   U7024 : BUF_X1 port map( A => n7595, Z => n14896);
   U7025 : BUF_X1 port map( A => n7584, Z => n14937);
   U7026 : BUF_X1 port map( A => n7585, Z => n14931);
   U7027 : BUF_X1 port map( A => n7587, Z => n14925);
   U7028 : BUF_X1 port map( A => n7589, Z => n14919);
   U7029 : BUF_X1 port map( A => n7590, Z => n14913);
   U7030 : BUF_X1 port map( A => n7591, Z => n14907);
   U7031 : BUF_X1 port map( A => n7593, Z => n14901);
   U7032 : BUF_X1 port map( A => n7595, Z => n14895);
   U7033 : AOI221_X1 port map( B1 => n8799, B2 => n13910, C1 => n8768, C2 => 
                           n13905, A => n5225, ZN => n5222);
   U7034 : OAI22_X1 port map( A1 => n13904, A2 => n710, B1 => n13901, B2 => 
                           n686, ZN => n5225);
   U7035 : AOI221_X1 port map( B1 => n8894, B2 => n13910, C1 => n8895, C2 => 
                           n13905, A => n4050, ZN => n4040);
   U7036 : OAI22_X1 port map( A1 => n13904, A2 => n40, B1 => n13901, B2 => n32,
                           ZN => n4050);
   U7037 : OAI22_X1 port map( A1 => n824, A2 => n3312, B1 => n823, B2 => n3313,
                           ZN => n3535);
   U7038 : OAI22_X1 port map( A1 => n6756, A2 => n14168, B1 => n14167, B2 => 
                           n139, ZN => n2832);
   U7039 : OAI22_X1 port map( A1 => n6762, A2 => n14122, B1 => n14121, B2 => 
                           n235, ZN => n2856);
   U7040 : OAI22_X1 port map( A1 => n6786, A2 => n14122, B1 => n14121, B2 => 
                           n234, ZN => n2906);
   U7041 : OAI22_X1 port map( A1 => n6804, A2 => n14168, B1 => n14167, B2 => 
                           n137, ZN => n2935);
   U7042 : OAI22_X1 port map( A1 => n6810, A2 => n14122, B1 => n14121, B2 => 
                           n233, ZN => n2943);
   U7043 : OAI22_X1 port map( A1 => n6828, A2 => n14168, B1 => n14167, B2 => 
                           n136, ZN => n2972);
   U7044 : OAI22_X1 port map( A1 => n6834, A2 => n14122, B1 => n14121, B2 => 
                           n232, ZN => n2980);
   U7045 : OAI22_X1 port map( A1 => n6852, A2 => n14168, B1 => n14167, B2 => 
                           n135, ZN => n3009);
   U7046 : OAI22_X1 port map( A1 => n6858, A2 => n14122, B1 => n14121, B2 => 
                           n231, ZN => n3017);
   U7047 : OAI22_X1 port map( A1 => n6876, A2 => n14168, B1 => n14167, B2 => 
                           n134, ZN => n3046);
   U7048 : OAI22_X1 port map( A1 => n6882, A2 => n14122, B1 => n14121, B2 => 
                           n230, ZN => n3054);
   U7049 : OAI22_X1 port map( A1 => n6900, A2 => n14168, B1 => n14167, B2 => 
                           n133, ZN => n3083);
   U7050 : OAI22_X1 port map( A1 => n6906, A2 => n14122, B1 => n14121, B2 => 
                           n229, ZN => n3091);
   U7051 : OAI22_X1 port map( A1 => n6924, A2 => n14168, B1 => n14167, B2 => 
                           n1303, ZN => n3120);
   U7052 : OAI22_X1 port map( A1 => n6930, A2 => n14122, B1 => n14121, B2 => 
                           n1574, ZN => n3128);
   U7053 : OAI22_X1 port map( A1 => n829, A2 => n13779, B1 => n828, B2 => 
                           n13776, ZN => n6071);
   U7054 : OAI22_X1 port map( A1 => n811, A2 => n13833, B1 => n810, B2 => 
                           n13830, ZN => n6063);
   U7055 : OAI22_X1 port map( A1 => n802, A2 => n13806, B1 => n801, B2 => 
                           n13803, ZN => n6065);
   U7056 : OAI22_X1 port map( A1 => n6742, A2 => n2846, B1 => n6741, B2 => 
                           n2847, ZN => n6592);
   U7057 : OAI22_X1 port map( A1 => n6766, A2 => n2846, B1 => n6765, B2 => 
                           n2847, ZN => n2845);
   U7058 : OAI22_X1 port map( A1 => n6790, A2 => n2846, B1 => n6789, B2 => 
                           n2847, ZN => n2904);
   U7059 : OAI22_X1 port map( A1 => n6814, A2 => n14148, B1 => n6813, B2 => 
                           n14146, ZN => n2941);
   U7060 : OAI22_X1 port map( A1 => n6838, A2 => n14148, B1 => n6837, B2 => 
                           n14146, ZN => n2978);
   U7061 : OAI22_X1 port map( A1 => n6862, A2 => n14148, B1 => n6861, B2 => 
                           n14146, ZN => n3015);
   U7062 : OAI22_X1 port map( A1 => n6886, A2 => n14148, B1 => n6885, B2 => 
                           n14146, ZN => n3052);
   U7063 : OAI22_X1 port map( A1 => n6910, A2 => n14148, B1 => n6909, B2 => 
                           n14146, ZN => n3089);
   U7064 : OAI22_X1 port map( A1 => n6934, A2 => n14148, B1 => n6933, B2 => 
                           n14146, ZN => n3126);
   U7065 : OAI22_X1 port map( A1 => n6958, A2 => n14148, B1 => n6957, B2 => 
                           n14146, ZN => n3163);
   U7066 : OAI22_X1 port map( A1 => n6982, A2 => n14148, B1 => n6981, B2 => 
                           n14146, ZN => n3200);
   U7067 : OAI22_X1 port map( A1 => n7006, A2 => n14148, B1 => n7005, B2 => 
                           n14146, ZN => n3237);
   U7068 : OAI22_X1 port map( A1 => n7030, A2 => n14148, B1 => n7029, B2 => 
                           n14146, ZN => n3274);
   U7069 : OAI22_X1 port map( A1 => n7150, A2 => n14148, B1 => n7149, B2 => 
                           n14146, ZN => n3461);
   U7070 : OAI22_X1 port map( A1 => n7174, A2 => n14148, B1 => n7173, B2 => 
                           n14146, ZN => n3498);
   U7071 : OAI22_X1 port map( A1 => n7246, A2 => n2846, B1 => n7245, B2 => 
                           n2847, ZN => n3609);
   U7072 : OAI22_X1 port map( A1 => n7270, A2 => n2846, B1 => n7269, B2 => 
                           n2847, ZN => n3646);
   U7073 : OAI22_X1 port map( A1 => n7294, A2 => n2846, B1 => n7293, B2 => 
                           n2847, ZN => n3683);
   U7074 : OAI22_X1 port map( A1 => n7318, A2 => n2846, B1 => n7317, B2 => 
                           n2847, ZN => n3720);
   U7075 : OAI22_X1 port map( A1 => n7342, A2 => n2846, B1 => n7341, B2 => 
                           n2847, ZN => n3757);
   U7076 : OAI22_X1 port map( A1 => n7366, A2 => n2846, B1 => n7365, B2 => 
                           n2847, ZN => n3794);
   U7077 : OAI22_X1 port map( A1 => n7390, A2 => n2846, B1 => n7389, B2 => 
                           n2847, ZN => n3831);
   U7078 : OAI22_X1 port map( A1 => n7414, A2 => n14148, B1 => n7413, B2 => 
                           n2847, ZN => n3868);
   U7079 : OAI22_X1 port map( A1 => n7486, A2 => n2846, B1 => n7485, B2 => 
                           n14146, ZN => n5264);
   U7080 : OAI22_X1 port map( A1 => n7438, A2 => n14148, B1 => n7437, B2 => 
                           n2847, ZN => n3905);
   U7081 : OAI22_X1 port map( A1 => n7462, A2 => n2846, B1 => n7461, B2 => 
                           n14146, ZN => n3942);
   U7082 : OAI22_X1 port map( A1 => n828, A2 => n13999, B1 => n829, B2 => 
                           n13996, ZN => n4750);
   U7083 : OAI22_X1 port map( A1 => n7648, A2 => n14027, B1 => n350, B2 => 
                           n14024, ZN => n4263);
   U7084 : OAI22_X1 port map( A1 => n7684, A2 => n14027, B1 => n356, B2 => 
                           n14024, ZN => n3985);
   U7085 : OAI22_X1 port map( A1 => n7678, A2 => n14027, B1 => n355, B2 => 
                           n14024, ZN => n4076);
   U7086 : OAI22_X1 port map( A1 => n7672, A2 => n14027, B1 => n354, B2 => 
                           n14024, ZN => n4115);
   U7087 : OAI22_X1 port map( A1 => n7666, A2 => n14027, B1 => n353, B2 => 
                           n14024, ZN => n4152);
   U7088 : OAI22_X1 port map( A1 => n7660, A2 => n14027, B1 => n352, B2 => 
                           n14024, ZN => n4189);
   U7089 : OAI22_X1 port map( A1 => n7654, A2 => n14027, B1 => n351, B2 => 
                           n14024, ZN => n4226);
   U7090 : OAI22_X1 port map( A1 => n7642, A2 => n14027, B1 => n349, B2 => 
                           n14024, ZN => n4300);
   U7091 : OAI22_X1 port map( A1 => n7646, A2 => n14054, B1 => n286, B2 => 
                           n14051, ZN => n4261);
   U7092 : OAI22_X1 port map( A1 => n7682, A2 => n14054, B1 => n292, B2 => 
                           n14051, ZN => n3974);
   U7093 : OAI22_X1 port map( A1 => n7676, A2 => n14054, B1 => n291, B2 => 
                           n14051, ZN => n4074);
   U7094 : OAI22_X1 port map( A1 => n7670, A2 => n14054, B1 => n290, B2 => 
                           n14051, ZN => n4113);
   U7095 : OAI22_X1 port map( A1 => n7664, A2 => n14054, B1 => n289, B2 => 
                           n14051, ZN => n4150);
   U7096 : OAI22_X1 port map( A1 => n7658, A2 => n14054, B1 => n288, B2 => 
                           n14051, ZN => n4187);
   U7097 : OAI22_X1 port map( A1 => n7652, A2 => n14054, B1 => n287, B2 => 
                           n14051, ZN => n4224);
   U7098 : OAI22_X1 port map( A1 => n7640, A2 => n14054, B1 => n285, B2 => 
                           n14051, ZN => n4298);
   U7099 : AOI221_X1 port map( B1 => n13651, B2 => n8670, C1 => n13648, C2 => 
                           n8702, A => n5423, ZN => n5416);
   U7100 : OAI22_X1 port map( A1 => n122, A2 => n13645, B1 => n130, B2 => 
                           n13642, ZN => n5423);
   U7101 : AOI221_X1 port map( B1 => n13651, B2 => n8668, C1 => n13648, C2 => 
                           n8700, A => n5497, ZN => n5490);
   U7102 : OAI22_X1 port map( A1 => n120, A2 => n13645, B1 => n128, B2 => 
                           n13642, ZN => n5497);
   U7103 : AOI221_X1 port map( B1 => n13651, B2 => n8667, C1 => n13648, C2 => 
                           n8699, A => n5534, ZN => n5527);
   U7104 : OAI22_X1 port map( A1 => n119, A2 => n13645, B1 => n127, B2 => 
                           n13642, ZN => n5534);
   U7105 : AOI221_X1 port map( B1 => n13651, B2 => n8666, C1 => n13648, C2 => 
                           n8698, A => n5571, ZN => n5564);
   U7106 : OAI22_X1 port map( A1 => n118, A2 => n13645, B1 => n126, B2 => 
                           n13642, ZN => n5571);
   U7107 : AOI221_X1 port map( B1 => n13651, B2 => n8665, C1 => n13648, C2 => 
                           n8697, A => n5608, ZN => n5601);
   U7108 : OAI22_X1 port map( A1 => n117, A2 => n13645, B1 => n125, B2 => 
                           n13642, ZN => n5608);
   U7109 : AOI221_X1 port map( B1 => n13651, B2 => n8669, C1 => n13648, C2 => 
                           n8701, A => n5460, ZN => n5453);
   U7110 : OAI22_X1 port map( A1 => n121, A2 => n13645, B1 => n129, B2 => 
                           n13642, ZN => n5460);
   U7111 : AOI221_X1 port map( B1 => n13883, B2 => n8678, C1 => n13880, C2 => 
                           n8646, A => n4990, ZN => n4983);
   U7112 : OAI22_X1 port map( A1 => n1271, A2 => n13877, B1 => n1247, B2 => 
                           n13874, ZN => n4990);
   U7113 : AOI221_X1 port map( B1 => n13883, B2 => n8677, C1 => n13880, C2 => 
                           n8645, A => n5027, ZN => n5020);
   U7114 : OAI22_X1 port map( A1 => n1270, A2 => n13877, B1 => n1246, B2 => 
                           n13874, ZN => n5027);
   U7115 : AOI221_X1 port map( B1 => n13883, B2 => n8676, C1 => n13880, C2 => 
                           n8644, A => n5064, ZN => n5057);
   U7116 : OAI22_X1 port map( A1 => n1269, A2 => n13877, B1 => n1245, B2 => 
                           n13874, ZN => n5064);
   U7117 : AOI221_X1 port map( B1 => n13883, B2 => n8675, C1 => n13880, C2 => 
                           n8643, A => n5101, ZN => n5094);
   U7118 : OAI22_X1 port map( A1 => n1268, A2 => n13877, B1 => n1244, B2 => 
                           n13874, ZN => n5101);
   U7119 : AOI221_X1 port map( B1 => n13883, B2 => n8674, C1 => n13880, C2 => 
                           n8642, A => n5138, ZN => n5131);
   U7120 : OAI22_X1 port map( A1 => n1267, A2 => n13877, B1 => n1243, B2 => 
                           n13874, ZN => n5138);
   U7121 : AOI221_X1 port map( B1 => n13883, B2 => n8673, C1 => n13878, C2 => 
                           n8641, A => n5175, ZN => n5168);
   U7122 : OAI22_X1 port map( A1 => n1266, A2 => n13877, B1 => n1242, B2 => 
                           n13874, ZN => n5175);
   U7123 : OAI22_X1 port map( A1 => n7496, A2 => n14052, B1 => n460, B2 => 
                           n14049, ZN => n5193);
   U7124 : OAI22_X1 port map( A1 => n7498, A2 => n14025, B1 => n556, B2 => 
                           n14022, ZN => n5199);
   U7125 : OAI22_X1 port map( A1 => n7562, A2 => n14052, B1 => n471, B2 => 
                           n14049, ZN => n4779);
   U7126 : OAI22_X1 port map( A1 => n7564, A2 => n14025, B1 => n567, B2 => 
                           n14022, ZN => n4781);
   U7127 : OAI22_X1 port map( A1 => n756, A2 => n13971, B1 => n1679, B2 => 
                           n13968, ZN => n4789);
   U7128 : OAI22_X1 port map( A1 => n7556, A2 => n14052, B1 => n470, B2 => 
                           n14049, ZN => n4816);
   U7129 : OAI22_X1 port map( A1 => n7558, A2 => n14025, B1 => n566, B2 => 
                           n14022, ZN => n4818);
   U7130 : OAI22_X1 port map( A1 => n7550, A2 => n14052, B1 => n469, B2 => 
                           n14049, ZN => n4853);
   U7131 : OAI22_X1 port map( A1 => n7552, A2 => n14025, B1 => n565, B2 => 
                           n14022, ZN => n4855);
   U7132 : OAI22_X1 port map( A1 => n7544, A2 => n14052, B1 => n468, B2 => 
                           n14049, ZN => n4890);
   U7133 : OAI22_X1 port map( A1 => n7546, A2 => n14025, B1 => n564, B2 => 
                           n14022, ZN => n4892);
   U7134 : OAI22_X1 port map( A1 => n7538, A2 => n14052, B1 => n467, B2 => 
                           n14049, ZN => n4927);
   U7135 : OAI22_X1 port map( A1 => n7540, A2 => n14025, B1 => n563, B2 => 
                           n14022, ZN => n4929);
   U7136 : OAI22_X1 port map( A1 => n756, A2 => n13751, B1 => n1679, B2 => 
                           n13748, ZN => n6110);
   U7137 : OAI22_X1 port map( A1 => n7574, A2 => n14053, B1 => n473, B2 => 
                           n14050, ZN => n4705);
   U7138 : OAI22_X1 port map( A1 => n7576, A2 => n14026, B1 => n569, B2 => 
                           n14023, ZN => n4707);
   U7139 : OAI22_X1 port map( A1 => n820, A2 => n13972, B1 => n1680, B2 => 
                           n13969, ZN => n4752);
   U7140 : OAI22_X1 port map( A1 => n820, A2 => n13752, B1 => n1680, B2 => 
                           n13749, ZN => n6073);
   U7141 : OAI22_X1 port map( A1 => n7532, A2 => n14052, B1 => n466, B2 => 
                           n14049, ZN => n4964);
   U7142 : OAI22_X1 port map( A1 => n7534, A2 => n14025, B1 => n562, B2 => 
                           n14022, ZN => n4966);
   U7143 : OAI22_X1 port map( A1 => n7526, A2 => n14052, B1 => n465, B2 => 
                           n14049, ZN => n5001);
   U7144 : OAI22_X1 port map( A1 => n7528, A2 => n14025, B1 => n561, B2 => 
                           n14022, ZN => n5003);
   U7145 : OAI22_X1 port map( A1 => n7520, A2 => n14052, B1 => n464, B2 => 
                           n14049, ZN => n5038);
   U7146 : OAI22_X1 port map( A1 => n7522, A2 => n14025, B1 => n560, B2 => 
                           n14022, ZN => n5040);
   U7147 : OAI22_X1 port map( A1 => n7514, A2 => n14052, B1 => n463, B2 => 
                           n14049, ZN => n5075);
   U7148 : OAI22_X1 port map( A1 => n7516, A2 => n14025, B1 => n559, B2 => 
                           n14022, ZN => n5077);
   U7149 : OAI22_X1 port map( A1 => n7508, A2 => n14052, B1 => n462, B2 => 
                           n14049, ZN => n5112);
   U7150 : OAI22_X1 port map( A1 => n7510, A2 => n14025, B1 => n558, B2 => 
                           n14022, ZN => n5114);
   U7151 : OAI22_X1 port map( A1 => n7502, A2 => n14052, B1 => n461, B2 => 
                           n14049, ZN => n5149);
   U7152 : OAI22_X1 port map( A1 => n7504, A2 => n14025, B1 => n557, B2 => 
                           n14022, ZN => n5151);
   U7153 : OAI22_X1 port map( A1 => n7634, A2 => n14053, B1 => n483, B2 => 
                           n14050, ZN => n4335);
   U7154 : OAI22_X1 port map( A1 => n7636, A2 => n14026, B1 => n579, B2 => 
                           n14023, ZN => n4337);
   U7155 : OAI22_X1 port map( A1 => n7628, A2 => n14053, B1 => n482, B2 => 
                           n14050, ZN => n4372);
   U7156 : OAI22_X1 port map( A1 => n7630, A2 => n14026, B1 => n578, B2 => 
                           n14023, ZN => n4374);
   U7157 : OAI22_X1 port map( A1 => n6948, A2 => n14168, B1 => n14166, B2 => 
                           n1302, ZN => n3157);
   U7158 : OAI22_X1 port map( A1 => n6954, A2 => n14122, B1 => n14120, B2 => 
                           n1573, ZN => n3165);
   U7159 : OAI22_X1 port map( A1 => n7622, A2 => n14053, B1 => n481, B2 => 
                           n14050, ZN => n4409);
   U7160 : OAI22_X1 port map( A1 => n7624, A2 => n14026, B1 => n577, B2 => 
                           n14023, ZN => n4411);
   U7161 : OAI22_X1 port map( A1 => n6972, A2 => n14168, B1 => n14166, B2 => 
                           n1301, ZN => n3194);
   U7162 : OAI22_X1 port map( A1 => n6978, A2 => n14122, B1 => n14120, B2 => 
                           n1572, ZN => n3202);
   U7163 : OAI22_X1 port map( A1 => n7616, A2 => n14053, B1 => n480, B2 => 
                           n14050, ZN => n4446);
   U7164 : OAI22_X1 port map( A1 => n7618, A2 => n14026, B1 => n576, B2 => 
                           n14023, ZN => n4448);
   U7165 : OAI22_X1 port map( A1 => n6996, A2 => n14168, B1 => n14166, B2 => 
                           n1300, ZN => n3231);
   U7166 : OAI22_X1 port map( A1 => n7002, A2 => n14122, B1 => n14120, B2 => 
                           n1571, ZN => n3239);
   U7167 : OAI22_X1 port map( A1 => n7610, A2 => n14053, B1 => n479, B2 => 
                           n14050, ZN => n4483);
   U7168 : OAI22_X1 port map( A1 => n7612, A2 => n14026, B1 => n575, B2 => 
                           n14023, ZN => n4485);
   U7169 : OAI22_X1 port map( A1 => n7020, A2 => n14168, B1 => n14166, B2 => 
                           n1299, ZN => n3268);
   U7170 : OAI22_X1 port map( A1 => n7604, A2 => n14053, B1 => n478, B2 => 
                           n14050, ZN => n4520);
   U7171 : OAI22_X1 port map( A1 => n7606, A2 => n14026, B1 => n574, B2 => 
                           n14023, ZN => n4522);
   U7172 : OAI22_X1 port map( A1 => n7598, A2 => n14053, B1 => n477, B2 => 
                           n14050, ZN => n4557);
   U7173 : OAI22_X1 port map( A1 => n7600, A2 => n14026, B1 => n573, B2 => 
                           n14023, ZN => n4559);
   U7174 : OAI22_X1 port map( A1 => n7592, A2 => n14053, B1 => n476, B2 => 
                           n14050, ZN => n4594);
   U7175 : OAI22_X1 port map( A1 => n7594, A2 => n14026, B1 => n572, B2 => 
                           n14023, ZN => n4596);
   U7176 : OAI22_X1 port map( A1 => n7586, A2 => n14053, B1 => n475, B2 => 
                           n14050, ZN => n4631);
   U7177 : OAI22_X1 port map( A1 => n7588, A2 => n14026, B1 => n571, B2 => 
                           n14023, ZN => n4633);
   U7178 : OAI22_X1 port map( A1 => n7580, A2 => n14053, B1 => n474, B2 => 
                           n14050, ZN => n4668);
   U7179 : OAI22_X1 port map( A1 => n7582, A2 => n14026, B1 => n570, B2 => 
                           n14023, ZN => n4670);
   U7180 : OAI22_X1 port map( A1 => n7146, A2 => n14122, B1 => n14120, B2 => 
                           n1565, ZN => n3463);
   U7181 : AOI221_X1 port map( B1 => n13649, B2 => n8651, C1 => n13646, C2 => 
                           n8683, A => n6126, ZN => n6119);
   U7182 : OAI22_X1 port map( A1 => n786, A2 => n13643, B1 => n1276, B2 => 
                           n13640, ZN => n6126);
   U7183 : AOI221_X1 port map( B1 => n13649, B2 => n8650, C1 => n13646, C2 => 
                           n8682, A => n6163, ZN => n6156);
   U7184 : OAI22_X1 port map( A1 => n1251, A2 => n13643, B1 => n1275, B2 => 
                           n13640, ZN => n6163);
   U7185 : AOI221_X1 port map( B1 => n13649, B2 => n8649, C1 => n13646, C2 => 
                           n8681, A => n6200, ZN => n6193);
   U7186 : OAI22_X1 port map( A1 => n1250, A2 => n13643, B1 => n1274, B2 => 
                           n13640, ZN => n6200);
   U7187 : AOI221_X1 port map( B1 => n13649, B2 => n8648, C1 => n13646, C2 => 
                           n8680, A => n6237, ZN => n6230);
   U7188 : OAI22_X1 port map( A1 => n1249, A2 => n13643, B1 => n1273, B2 => 
                           n13640, ZN => n6237);
   U7189 : AOI221_X1 port map( B1 => n13649, B2 => n8647, C1 => n13646, C2 => 
                           n8679, A => n6274, ZN => n6267);
   U7190 : OAI22_X1 port map( A1 => n1248, A2 => n13643, B1 => n1272, B2 => 
                           n13640, ZN => n6274);
   U7191 : AOI221_X1 port map( B1 => n13649, B2 => n8646, C1 => n13646, C2 => 
                           n8678, A => n6311, ZN => n6304);
   U7192 : OAI22_X1 port map( A1 => n1247, A2 => n13643, B1 => n1271, B2 => 
                           n13640, ZN => n6311);
   U7193 : AOI221_X1 port map( B1 => n13649, B2 => n8645, C1 => n13646, C2 => 
                           n8677, A => n6348, ZN => n6341);
   U7194 : OAI22_X1 port map( A1 => n1246, A2 => n13643, B1 => n1270, B2 => 
                           n13640, ZN => n6348);
   U7195 : AOI221_X1 port map( B1 => n13649, B2 => n8644, C1 => n13646, C2 => 
                           n8676, A => n6385, ZN => n6378);
   U7196 : OAI22_X1 port map( A1 => n1245, A2 => n13643, B1 => n1269, B2 => 
                           n13640, ZN => n6385);
   U7197 : AOI221_X1 port map( B1 => n13649, B2 => n8643, C1 => n13646, C2 => 
                           n8675, A => n6422, ZN => n6415);
   U7198 : OAI22_X1 port map( A1 => n1244, A2 => n13643, B1 => n1268, B2 => 
                           n13640, ZN => n6422);
   U7199 : AOI221_X1 port map( B1 => n13649, B2 => n8642, C1 => n13646, C2 => 
                           n8674, A => n6459, ZN => n6452);
   U7200 : OAI22_X1 port map( A1 => n1243, A2 => n13643, B1 => n1267, B2 => 
                           n13640, ZN => n6459);
   U7201 : AOI221_X1 port map( B1 => n13649, B2 => n8641, C1 => n13646, C2 => 
                           n8673, A => n6496, ZN => n6489);
   U7202 : OAI22_X1 port map( A1 => n1242, A2 => n13643, B1 => n1266, B2 => 
                           n13640, ZN => n6496);
   U7203 : AOI221_X1 port map( B1 => n13703, B2 => n2327, C1 => n13700, C2 => 
                           n831, A => n6540, ZN => n6531);
   U7204 : OAI22_X1 port map( A1 => n1512, A2 => n13697, B1 => n1536, B2 => 
                           n13694, ZN => n6540);
   U7205 : OAI22_X1 port map( A1 => n14936, A2 => n14276, B1 => n6559, B2 => 
                           n14285, ZN => n11501);
   U7206 : NOR4_X1 port map( A1 => n6560, A2 => n6561, A3 => n6562, A4 => n6563
                           , ZN => n6559);
   U7207 : NAND4_X1 port map( A1 => n6595, A2 => n6596, A3 => n6597, A4 => 
                           n6598, ZN => n6560);
   U7208 : OAI22_X1 port map( A1 => n14930, A2 => n14276, B1 => n2777, B2 => 
                           n14278, ZN => n9226);
   U7209 : NOR4_X1 port map( A1 => n2779, A2 => n2780, A3 => n2781, A4 => n2782
                           , ZN => n2777);
   U7210 : NAND4_X1 port map( A1 => n2859, A2 => n2860, A3 => n2861, A4 => 
                           n2862, ZN => n2779);
   U7211 : OAI22_X1 port map( A1 => n14924, A2 => n14276, B1 => n2878, B2 => 
                           n14278, ZN => n9224);
   U7212 : NOR4_X1 port map( A1 => n2879, A2 => n2880, A3 => n2881, A4 => n2882
                           , ZN => n2878);
   U7213 : NAND4_X1 port map( A1 => n2907, A2 => n2908, A3 => n2909, A4 => 
                           n2910, ZN => n2879);
   U7214 : OAI22_X1 port map( A1 => n14918, A2 => n14276, B1 => n2915, B2 => 
                           n14278, ZN => n9222);
   U7215 : NOR4_X1 port map( A1 => n2916, A2 => n2917, A3 => n2918, A4 => n2919
                           , ZN => n2915);
   U7216 : NAND4_X1 port map( A1 => n2944, A2 => n2945, A3 => n2946, A4 => 
                           n2947, ZN => n2916);
   U7217 : OAI22_X1 port map( A1 => n14912, A2 => n14276, B1 => n2952, B2 => 
                           n14278, ZN => n9220);
   U7218 : NOR4_X1 port map( A1 => n2953, A2 => n2954, A3 => n2955, A4 => n2956
                           , ZN => n2952);
   U7219 : NAND4_X1 port map( A1 => n2981, A2 => n2982, A3 => n2983, A4 => 
                           n2984, ZN => n2953);
   U7220 : OAI22_X1 port map( A1 => n14906, A2 => n14276, B1 => n2989, B2 => 
                           n14279, ZN => n9218);
   U7221 : NOR4_X1 port map( A1 => n2990, A2 => n2991, A3 => n2992, A4 => n2993
                           , ZN => n2989);
   U7222 : NAND4_X1 port map( A1 => n3018, A2 => n3019, A3 => n3020, A4 => 
                           n3021, ZN => n2990);
   U7223 : OAI22_X1 port map( A1 => n14900, A2 => n14276, B1 => n3026, B2 => 
                           n14279, ZN => n9216);
   U7224 : NOR4_X1 port map( A1 => n3027, A2 => n3028, A3 => n3029, A4 => n3030
                           , ZN => n3026);
   U7225 : NAND4_X1 port map( A1 => n3055, A2 => n3056, A3 => n3057, A4 => 
                           n3058, ZN => n3027);
   U7226 : OAI22_X1 port map( A1 => n14894, A2 => n14276, B1 => n3063, B2 => 
                           n14279, ZN => n9214);
   U7227 : NOR4_X1 port map( A1 => n3064, A2 => n3065, A3 => n3066, A4 => n3067
                           , ZN => n3063);
   U7228 : NAND4_X1 port map( A1 => n3092, A2 => n3093, A3 => n3094, A4 => 
                           n3095, ZN => n3064);
   U7229 : OAI22_X1 port map( A1 => n14891, A2 => n14276, B1 => n3100, B2 => 
                           n14279, ZN => n9212);
   U7230 : NOR4_X1 port map( A1 => n3101, A2 => n3102, A3 => n3103, A4 => n3104
                           , ZN => n3100);
   U7231 : NAND4_X1 port map( A1 => n3129, A2 => n3130, A3 => n3131, A4 => 
                           n3132, ZN => n3101);
   U7232 : OAI22_X1 port map( A1 => n14885, A2 => n14276, B1 => n3137, B2 => 
                           n14280, ZN => n9210);
   U7233 : NOR4_X1 port map( A1 => n3138, A2 => n3139, A3 => n3140, A4 => n3141
                           , ZN => n3137);
   U7234 : NAND4_X1 port map( A1 => n3166, A2 => n3167, A3 => n3168, A4 => 
                           n3169, ZN => n3138);
   U7235 : OAI22_X1 port map( A1 => n14879, A2 => n14276, B1 => n3174, B2 => 
                           n14280, ZN => n9208);
   U7236 : NOR4_X1 port map( A1 => n3175, A2 => n3176, A3 => n3177, A4 => n3178
                           , ZN => n3174);
   U7237 : NAND4_X1 port map( A1 => n3203, A2 => n3204, A3 => n3205, A4 => 
                           n3206, ZN => n3175);
   U7238 : OAI22_X1 port map( A1 => n14873, A2 => n14276, B1 => n3211, B2 => 
                           n14280, ZN => n9206);
   U7239 : NOR4_X1 port map( A1 => n3212, A2 => n3213, A3 => n3214, A4 => n3215
                           , ZN => n3211);
   U7240 : NAND4_X1 port map( A1 => n3240, A2 => n3241, A3 => n3242, A4 => 
                           n3243, ZN => n3212);
   U7241 : OAI22_X1 port map( A1 => n14867, A2 => n14276, B1 => n3248, B2 => 
                           n14280, ZN => n9204);
   U7242 : NOR4_X1 port map( A1 => n3249, A2 => n3250, A3 => n3251, A4 => n3252
                           , ZN => n3248);
   U7243 : NAND4_X1 port map( A1 => n3277, A2 => n3278, A3 => n3279, A4 => 
                           n3280, ZN => n3249);
   U7244 : OAI22_X1 port map( A1 => n14861, A2 => n14277, B1 => n3285, B2 => 
                           n14281, ZN => n9202);
   U7245 : NOR4_X1 port map( A1 => n3286, A2 => n3287, A3 => n3288, A4 => n3289
                           , ZN => n3285);
   U7246 : NAND4_X1 port map( A1 => n3316, A2 => n3317, A3 => n3318, A4 => 
                           n3319, ZN => n3286);
   U7247 : OAI22_X1 port map( A1 => n14855, A2 => n14277, B1 => n3324, B2 => 
                           n14281, ZN => n9200);
   U7248 : NOR4_X1 port map( A1 => n3325, A2 => n3326, A3 => n3327, A4 => n3328
                           , ZN => n3324);
   U7249 : NAND4_X1 port map( A1 => n3353, A2 => n3354, A3 => n3355, A4 => 
                           n3356, ZN => n3325);
   U7250 : OAI22_X1 port map( A1 => n14849, A2 => n14277, B1 => n3361, B2 => 
                           n14281, ZN => n9198);
   U7251 : NOR4_X1 port map( A1 => n3362, A2 => n3363, A3 => n3364, A4 => n3365
                           , ZN => n3361);
   U7252 : NAND4_X1 port map( A1 => n3390, A2 => n3391, A3 => n3392, A4 => 
                           n3393, ZN => n3362);
   U7253 : OAI22_X1 port map( A1 => n14843, A2 => n14277, B1 => n3398, B2 => 
                           n14281, ZN => n9196);
   U7254 : NOR4_X1 port map( A1 => n3399, A2 => n3400, A3 => n3401, A4 => n3402
                           , ZN => n3398);
   U7255 : NAND4_X1 port map( A1 => n3427, A2 => n3428, A3 => n3429, A4 => 
                           n3430, ZN => n3399);
   U7256 : OAI22_X1 port map( A1 => n14837, A2 => n14277, B1 => n3435, B2 => 
                           n14282, ZN => n9194);
   U7257 : NOR4_X1 port map( A1 => n3436, A2 => n3437, A3 => n3438, A4 => n3439
                           , ZN => n3435);
   U7258 : NAND4_X1 port map( A1 => n3464, A2 => n3465, A3 => n3466, A4 => 
                           n3467, ZN => n3436);
   U7259 : OAI22_X1 port map( A1 => n14831, A2 => n14277, B1 => n3472, B2 => 
                           n14282, ZN => n9192);
   U7260 : NOR4_X1 port map( A1 => n3473, A2 => n3474, A3 => n3475, A4 => n3476
                           , ZN => n3472);
   U7261 : NAND4_X1 port map( A1 => n3501, A2 => n3502, A3 => n3503, A4 => 
                           n3504, ZN => n3473);
   U7262 : OAI22_X1 port map( A1 => n14825, A2 => n14277, B1 => n3509, B2 => 
                           n14282, ZN => n9190);
   U7263 : NOR4_X1 port map( A1 => n3510, A2 => n3511, A3 => n3512, A4 => n3513
                           , ZN => n3509);
   U7264 : NAND4_X1 port map( A1 => n3538, A2 => n3539, A3 => n3540, A4 => 
                           n3541, ZN => n3510);
   U7265 : OAI22_X1 port map( A1 => n14819, A2 => n14277, B1 => n3546, B2 => 
                           n14282, ZN => n9188);
   U7266 : NOR4_X1 port map( A1 => n3547, A2 => n3548, A3 => n3549, A4 => n3550
                           , ZN => n3546);
   U7267 : NAND4_X1 port map( A1 => n3575, A2 => n3576, A3 => n3577, A4 => 
                           n3578, ZN => n3547);
   U7268 : OAI22_X1 port map( A1 => n14813, A2 => n14277, B1 => n3583, B2 => 
                           n14283, ZN => n9186);
   U7269 : NOR4_X1 port map( A1 => n3584, A2 => n3585, A3 => n3586, A4 => n3587
                           , ZN => n3583);
   U7270 : NAND4_X1 port map( A1 => n3612, A2 => n3613, A3 => n3614, A4 => 
                           n3615, ZN => n3584);
   U7271 : OAI22_X1 port map( A1 => n14807, A2 => n14277, B1 => n3620, B2 => 
                           n14283, ZN => n9184);
   U7272 : NOR4_X1 port map( A1 => n3621, A2 => n3622, A3 => n3623, A4 => n3624
                           , ZN => n3620);
   U7273 : NAND4_X1 port map( A1 => n3649, A2 => n3650, A3 => n3651, A4 => 
                           n3652, ZN => n3621);
   U7274 : OAI22_X1 port map( A1 => n14801, A2 => n14277, B1 => n3657, B2 => 
                           n14283, ZN => n9182);
   U7275 : NOR4_X1 port map( A1 => n3658, A2 => n3659, A3 => n3660, A4 => n3661
                           , ZN => n3657);
   U7276 : NAND4_X1 port map( A1 => n3686, A2 => n3687, A3 => n3688, A4 => 
                           n3689, ZN => n3658);
   U7277 : OAI22_X1 port map( A1 => n14795, A2 => n14277, B1 => n3694, B2 => 
                           n14283, ZN => n9180);
   U7278 : NOR4_X1 port map( A1 => n3695, A2 => n3696, A3 => n3697, A4 => n3698
                           , ZN => n3694);
   U7279 : NAND4_X1 port map( A1 => n3723, A2 => n3724, A3 => n3725, A4 => 
                           n3726, ZN => n3695);
   U7280 : OAI22_X1 port map( A1 => n14789, A2 => n14277, B1 => n3731, B2 => 
                           n14284, ZN => n9178);
   U7281 : NOR4_X1 port map( A1 => n3732, A2 => n3733, A3 => n3734, A4 => n3735
                           , ZN => n3731);
   U7282 : NAND4_X1 port map( A1 => n3760, A2 => n3761, A3 => n3762, A4 => 
                           n3763, ZN => n3732);
   U7283 : OAI22_X1 port map( A1 => n14783, A2 => n14276, B1 => n3768, B2 => 
                           n14284, ZN => n9176);
   U7284 : NOR4_X1 port map( A1 => n3769, A2 => n3770, A3 => n3771, A4 => n3772
                           , ZN => n3768);
   U7285 : NAND4_X1 port map( A1 => n3797, A2 => n3798, A3 => n3799, A4 => 
                           n3800, ZN => n3769);
   U7286 : OAI22_X1 port map( A1 => n14777, A2 => n14277, B1 => n3805, B2 => 
                           n14284, ZN => n9174);
   U7287 : NOR4_X1 port map( A1 => n3806, A2 => n3807, A3 => n3808, A4 => n3809
                           , ZN => n3805);
   U7288 : NAND4_X1 port map( A1 => n3834, A2 => n3835, A3 => n3836, A4 => 
                           n3837, ZN => n3806);
   U7289 : OAI22_X1 port map( A1 => n14771, A2 => n14276, B1 => n3842, B2 => 
                           n14284, ZN => n9172);
   U7290 : NOR4_X1 port map( A1 => n3843, A2 => n3844, A3 => n3845, A4 => n3846
                           , ZN => n3842);
   U7291 : NAND4_X1 port map( A1 => n3871, A2 => n3872, A3 => n3873, A4 => 
                           n3874, ZN => n3843);
   U7292 : OAI22_X1 port map( A1 => n14766, A2 => n14277, B1 => n3879, B2 => 
                           n14285, ZN => n9170);
   U7293 : NOR4_X1 port map( A1 => n3880, A2 => n3881, A3 => n3882, A4 => n3883
                           , ZN => n3879);
   U7294 : NAND4_X1 port map( A1 => n3908, A2 => n3909, A3 => n3910, A4 => 
                           n3911, ZN => n3880);
   U7295 : OAI22_X1 port map( A1 => n14760, A2 => n14276, B1 => n3916, B2 => 
                           n14285, ZN => n9168);
   U7296 : NOR4_X1 port map( A1 => n3917, A2 => n3918, A3 => n3919, A4 => n3920
                           , ZN => n3916);
   U7297 : NAND4_X1 port map( A1 => n3945, A2 => n3946, A3 => n3947, A4 => 
                           n3948, ZN => n3917);
   U7298 : OAI22_X1 port map( A1 => n14753, A2 => n14277, B1 => n5238, B2 => 
                           n14285, ZN => n9134);
   U7299 : NOR4_X1 port map( A1 => n5239, A2 => n5240, A3 => n5241, A4 => n5242
                           , ZN => n5238);
   U7300 : NAND4_X1 port map( A1 => n5267, A2 => n5268, A3 => n5269, A4 => 
                           n5270, ZN => n5239);
   U7301 : NAND4_X1 port map( A1 => n3551, A2 => n3552, A3 => n3553, A4 => 
                           n3554, ZN => n3550);
   U7302 : AOI221_X1 port map( B1 => n800, B2 => n14230, C1 => n799, C2 => 
                           n14226, A => n3558, ZN => n3551);
   U7303 : AOI221_X1 port map( B1 => n8747, B2 => n14256, C1 => n8715, C2 => 
                           n14253, A => n3556, ZN => n3553);
   U7304 : AOI221_X1 port map( B1 => n798, B2 => n14245, C1 => n14242, C2 => 
                           n697, A => n3557, ZN => n3552);
   U7305 : NAND4_X1 port map( A1 => n3588, A2 => n3589, A3 => n3590, A4 => 
                           n3591, ZN => n3587);
   U7306 : AOI221_X1 port map( B1 => n736, B2 => n14230, C1 => n735, C2 => 
                           n14226, A => n3595, ZN => n3588);
   U7307 : AOI221_X1 port map( B1 => n8746, B2 => n14255, C1 => n8714, C2 => 
                           n14252, A => n3593, ZN => n3590);
   U7308 : AOI221_X1 port map( B1 => n734, B2 => n14245, C1 => n14242, C2 => 
                           n696, A => n3594, ZN => n3589);
   U7309 : NAND4_X1 port map( A1 => n4256, A2 => n4257, A3 => n4258, A4 => 
                           n4259, ZN => n4255);
   U7310 : AOI221_X1 port map( B1 => n14033, B2 => n7933, C1 => n14030, C2 => 
                           n7891, A => n4263, ZN => n4256);
   U7311 : AOI221_X1 port map( B1 => n14060, B2 => n8061, C1 => n14057, C2 => 
                           n8029, A => n4261, ZN => n4258);
   U7312 : AOI221_X1 port map( B1 => n14048, B2 => n7997, C1 => n14045, C2 => 
                           n7965, A => n4262, ZN => n4257);
   U7313 : NAND4_X1 port map( A1 => n5392, A2 => n5393, A3 => n5394, A4 => 
                           n5395, ZN => n5391);
   U7314 : AOI221_X1 port map( B1 => n13813, B2 => n1829, C1 => n13810, C2 => 
                           n835, A => n5399, ZN => n5392);
   U7315 : AOI221_X1 port map( B1 => n13840, B2 => n1821, C1 => n13837, C2 => 
                           n834, A => n5397, ZN => n5394);
   U7316 : AOI221_X1 port map( B1 => n13828, B2 => n8002, C1 => n13825, C2 => 
                           n7970, A => n5398, ZN => n5393);
   U7317 : NAND4_X1 port map( A1 => n5466, A2 => n5467, A3 => n5468, A4 => 
                           n5469, ZN => n5465);
   U7318 : AOI221_X1 port map( B1 => n13813, B2 => n1827, C1 => n13810, C2 => 
                           n839, A => n5473, ZN => n5466);
   U7319 : AOI221_X1 port map( B1 => n13840, B2 => n1819, C1 => n13837, C2 => 
                           n838, A => n5471, ZN => n5468);
   U7320 : AOI221_X1 port map( B1 => n13828, B2 => n8000, C1 => n13825, C2 => 
                           n7968, A => n5472, ZN => n5467);
   U7321 : NAND4_X1 port map( A1 => n5503, A2 => n5504, A3 => n5505, A4 => 
                           n5506, ZN => n5502);
   U7322 : AOI221_X1 port map( B1 => n13813, B2 => n1826, C1 => n13810, C2 => 
                           n841, A => n5510, ZN => n5503);
   U7323 : AOI221_X1 port map( B1 => n13840, B2 => n1818, C1 => n13837, C2 => 
                           n840, A => n5508, ZN => n5505);
   U7324 : AOI221_X1 port map( B1 => n13828, B2 => n7999, C1 => n13825, C2 => 
                           n7967, A => n5509, ZN => n5504);
   U7325 : NAND4_X1 port map( A1 => n5540, A2 => n5541, A3 => n5542, A4 => 
                           n5543, ZN => n5539);
   U7326 : AOI221_X1 port map( B1 => n13813, B2 => n1825, C1 => n13810, C2 => 
                           n843, A => n5547, ZN => n5540);
   U7327 : AOI221_X1 port map( B1 => n13840, B2 => n1817, C1 => n13837, C2 => 
                           n842, A => n5545, ZN => n5542);
   U7328 : AOI221_X1 port map( B1 => n13828, B2 => n7998, C1 => n13825, C2 => 
                           n7966, A => n5546, ZN => n5541);
   U7329 : NAND4_X1 port map( A1 => n5577, A2 => n5578, A3 => n5579, A4 => 
                           n5580, ZN => n5576);
   U7330 : AOI221_X1 port map( B1 => n13813, B2 => n1824, C1 => n13810, C2 => 
                           n845, A => n5584, ZN => n5577);
   U7331 : AOI221_X1 port map( B1 => n13840, B2 => n1816, C1 => n13837, C2 => 
                           n844, A => n5582, ZN => n5579);
   U7332 : AOI221_X1 port map( B1 => n13828, B2 => n7997, C1 => n13825, C2 => 
                           n7965, A => n5583, ZN => n5578);
   U7333 : NAND4_X1 port map( A1 => n5181, A2 => n5182, A3 => n5183, A4 => 
                           n5184, ZN => n5180);
   U7334 : AOI221_X1 port map( B1 => n14073, B2 => n8100, C1 => n14070, C2 => 
                           n8068, A => n5185, ZN => n5184);
   U7335 : AOI221_X1 port map( B1 => n14031, B2 => n7908, C1 => n14028, C2 => 
                           n7816, A => n5199, ZN => n5181);
   U7336 : AOI221_X1 port map( B1 => n14058, B2 => n8036, C1 => n14055, C2 => 
                           n8004, A => n5193, ZN => n5183);
   U7337 : NAND4_X1 port map( A1 => n4774, A2 => n4775, A3 => n4776, A4 => 
                           n4777, ZN => n4773);
   U7338 : AOI221_X1 port map( B1 => n14031, B2 => n7919, C1 => n14028, C2 => 
                           n7849, A => n4781, ZN => n4774);
   U7339 : AOI221_X1 port map( B1 => n14058, B2 => n8047, C1 => n14055, C2 => 
                           n8015, A => n4779, ZN => n4776);
   U7340 : AOI221_X1 port map( B1 => n14046, B2 => n7983, C1 => n14043, C2 => 
                           n7951, A => n4780, ZN => n4775);
   U7341 : NAND4_X1 port map( A1 => n4811, A2 => n4812, A3 => n4813, A4 => 
                           n4814, ZN => n4810);
   U7342 : AOI221_X1 port map( B1 => n14073, B2 => n8110, C1 => n14070, C2 => 
                           n8078, A => n4815, ZN => n4814);
   U7343 : AOI221_X1 port map( B1 => n14031, B2 => n7918, C1 => n14028, C2 => 
                           n7846, A => n4818, ZN => n4811);
   U7344 : AOI221_X1 port map( B1 => n14058, B2 => n8046, C1 => n14055, C2 => 
                           n8014, A => n4816, ZN => n4813);
   U7345 : NAND4_X1 port map( A1 => n4848, A2 => n4849, A3 => n4850, A4 => 
                           n4851, ZN => n4847);
   U7346 : AOI221_X1 port map( B1 => n14073, B2 => n8109, C1 => n14070, C2 => 
                           n8077, A => n4852, ZN => n4851);
   U7347 : AOI221_X1 port map( B1 => n14031, B2 => n7917, C1 => n14028, C2 => 
                           n7843, A => n4855, ZN => n4848);
   U7348 : AOI221_X1 port map( B1 => n14058, B2 => n8045, C1 => n14055, C2 => 
                           n8013, A => n4853, ZN => n4850);
   U7349 : NAND4_X1 port map( A1 => n4885, A2 => n4886, A3 => n4887, A4 => 
                           n4888, ZN => n4884);
   U7350 : AOI221_X1 port map( B1 => n14073, B2 => n8108, C1 => n14070, C2 => 
                           n8076, A => n4889, ZN => n4888);
   U7351 : AOI221_X1 port map( B1 => n14031, B2 => n7916, C1 => n14028, C2 => 
                           n7840, A => n4892, ZN => n4885);
   U7352 : AOI221_X1 port map( B1 => n14058, B2 => n8044, C1 => n14055, C2 => 
                           n8012, A => n4890, ZN => n4887);
   U7353 : NAND4_X1 port map( A1 => n4922, A2 => n4923, A3 => n4924, A4 => 
                           n4925, ZN => n4921);
   U7354 : AOI221_X1 port map( B1 => n14073, B2 => n8107, C1 => n14070, C2 => 
                           n8075, A => n4926, ZN => n4925);
   U7355 : AOI221_X1 port map( B1 => n14031, B2 => n7915, C1 => n14028, C2 => 
                           n7837, A => n4929, ZN => n4922);
   U7356 : AOI221_X1 port map( B1 => n14058, B2 => n8043, C1 => n14055, C2 => 
                           n8011, A => n4927, ZN => n4924);
   U7357 : NAND4_X1 port map( A1 => n6095, A2 => n6096, A3 => n6097, A4 => 
                           n6098, ZN => n6094);
   U7358 : AOI221_X1 port map( B1 => n13811, B2 => n1891, C1 => n13808, C2 => 
                           n873, A => n6102, ZN => n6095);
   U7359 : AOI221_X1 port map( B1 => n13838, B2 => n1867, C1 => n13835, C2 => 
                           n872, A => n6100, ZN => n6097);
   U7360 : AOI221_X1 port map( B1 => n13826, B2 => n7983, C1 => n13823, C2 => 
                           n7951, A => n6101, ZN => n6096);
   U7361 : NAND4_X1 port map( A1 => n6132, A2 => n6133, A3 => n6134, A4 => 
                           n6135, ZN => n6131);
   U7362 : AOI221_X1 port map( B1 => n13853, B2 => n8110, C1 => n13850, C2 => 
                           n8078, A => n6136, ZN => n6135);
   U7363 : AOI221_X1 port map( B1 => n13811, B2 => n1890, C1 => n13808, C2 => 
                           n875, A => n6139, ZN => n6132);
   U7364 : AOI221_X1 port map( B1 => n13838, B2 => n1866, C1 => n13835, C2 => 
                           n874, A => n6137, ZN => n6134);
   U7365 : NAND4_X1 port map( A1 => n6169, A2 => n6170, A3 => n6171, A4 => 
                           n6172, ZN => n6168);
   U7366 : AOI221_X1 port map( B1 => n13853, B2 => n8109, C1 => n13850, C2 => 
                           n8077, A => n6173, ZN => n6172);
   U7367 : AOI221_X1 port map( B1 => n13811, B2 => n1889, C1 => n13808, C2 => 
                           n877, A => n6176, ZN => n6169);
   U7368 : AOI221_X1 port map( B1 => n13838, B2 => n1865, C1 => n13835, C2 => 
                           n876, A => n6174, ZN => n6171);
   U7369 : NAND4_X1 port map( A1 => n6206, A2 => n6207, A3 => n6208, A4 => 
                           n6209, ZN => n6205);
   U7370 : AOI221_X1 port map( B1 => n13853, B2 => n8108, C1 => n13850, C2 => 
                           n8076, A => n6210, ZN => n6209);
   U7371 : AOI221_X1 port map( B1 => n13811, B2 => n1888, C1 => n13808, C2 => 
                           n879, A => n6213, ZN => n6206);
   U7372 : AOI221_X1 port map( B1 => n13838, B2 => n1864, C1 => n13835, C2 => 
                           n878, A => n6211, ZN => n6208);
   U7373 : NAND4_X1 port map( A1 => n6243, A2 => n6244, A3 => n6245, A4 => 
                           n6246, ZN => n6242);
   U7374 : AOI221_X1 port map( B1 => n13853, B2 => n8107, C1 => n13850, C2 => 
                           n8075, A => n6247, ZN => n6246);
   U7375 : AOI221_X1 port map( B1 => n13811, B2 => n1887, C1 => n13808, C2 => 
                           n881, A => n6250, ZN => n6243);
   U7376 : AOI221_X1 port map( B1 => n13838, B2 => n1863, C1 => n13835, C2 => 
                           n880, A => n6248, ZN => n6245);
   U7377 : NAND4_X1 port map( A1 => n6280, A2 => n6281, A3 => n6282, A4 => 
                           n6283, ZN => n6279);
   U7378 : AOI221_X1 port map( B1 => n13853, B2 => n8106, C1 => n13850, C2 => 
                           n8074, A => n6284, ZN => n6283);
   U7379 : AOI221_X1 port map( B1 => n13811, B2 => n1886, C1 => n13808, C2 => 
                           n883, A => n6287, ZN => n6280);
   U7380 : AOI221_X1 port map( B1 => n13838, B2 => n1862, C1 => n13835, C2 => 
                           n882, A => n6285, ZN => n6282);
   U7381 : NAND4_X1 port map( A1 => n6317, A2 => n6318, A3 => n6319, A4 => 
                           n6320, ZN => n6316);
   U7382 : AOI221_X1 port map( B1 => n13853, B2 => n8105, C1 => n13850, C2 => 
                           n8073, A => n6321, ZN => n6320);
   U7383 : AOI221_X1 port map( B1 => n13811, B2 => n1885, C1 => n13808, C2 => 
                           n885, A => n6324, ZN => n6317);
   U7384 : AOI221_X1 port map( B1 => n13838, B2 => n1861, C1 => n13835, C2 => 
                           n884, A => n6322, ZN => n6319);
   U7385 : NAND4_X1 port map( A1 => n6354, A2 => n6355, A3 => n6356, A4 => 
                           n6357, ZN => n6353);
   U7386 : AOI221_X1 port map( B1 => n13853, B2 => n8104, C1 => n13850, C2 => 
                           n8072, A => n6358, ZN => n6357);
   U7387 : AOI221_X1 port map( B1 => n13811, B2 => n1884, C1 => n13808, C2 => 
                           n887, A => n6361, ZN => n6354);
   U7388 : AOI221_X1 port map( B1 => n13838, B2 => n1860, C1 => n13835, C2 => 
                           n886, A => n6359, ZN => n6356);
   U7389 : NAND4_X1 port map( A1 => n6391, A2 => n6392, A3 => n6393, A4 => 
                           n6394, ZN => n6390);
   U7390 : AOI221_X1 port map( B1 => n13853, B2 => n8103, C1 => n13850, C2 => 
                           n8071, A => n6395, ZN => n6394);
   U7391 : AOI221_X1 port map( B1 => n13811, B2 => n1883, C1 => n13808, C2 => 
                           n889, A => n6398, ZN => n6391);
   U7392 : AOI221_X1 port map( B1 => n13838, B2 => n1859, C1 => n13835, C2 => 
                           n888, A => n6396, ZN => n6393);
   U7393 : NAND4_X1 port map( A1 => n6428, A2 => n6429, A3 => n6430, A4 => 
                           n6431, ZN => n6427);
   U7394 : AOI221_X1 port map( B1 => n13853, B2 => n8102, C1 => n13850, C2 => 
                           n8070, A => n6432, ZN => n6431);
   U7395 : AOI221_X1 port map( B1 => n13811, B2 => n1882, C1 => n13808, C2 => 
                           n891, A => n6435, ZN => n6428);
   U7396 : AOI221_X1 port map( B1 => n13838, B2 => n1858, C1 => n13835, C2 => 
                           n890, A => n6433, ZN => n6430);
   U7397 : NAND4_X1 port map( A1 => n6465, A2 => n6466, A3 => n6467, A4 => 
                           n6468, ZN => n6464);
   U7398 : AOI221_X1 port map( B1 => n13853, B2 => n8101, C1 => n13850, C2 => 
                           n8069, A => n6469, ZN => n6468);
   U7399 : AOI221_X1 port map( B1 => n13811, B2 => n1881, C1 => n13808, C2 => 
                           n893, A => n6472, ZN => n6465);
   U7400 : AOI221_X1 port map( B1 => n13838, B2 => n1857, C1 => n13835, C2 => 
                           n892, A => n6470, ZN => n6467);
   U7401 : NAND4_X1 port map( A1 => n4700, A2 => n4701, A3 => n4702, A4 => 
                           n4703, ZN => n4699);
   U7402 : AOI221_X1 port map( B1 => n14074, B2 => n8113, C1 => n14071, C2 => 
                           n8081, A => n4704, ZN => n4703);
   U7403 : AOI221_X1 port map( B1 => n14032, B2 => n7921, C1 => n14029, C2 => 
                           n7855, A => n4707, ZN => n4700);
   U7404 : AOI221_X1 port map( B1 => n14059, B2 => n8049, C1 => n14056, C2 => 
                           n8017, A => n4705, ZN => n4702);
   U7405 : NAND4_X1 port map( A1 => n6021, A2 => n6022, A3 => n6023, A4 => 
                           n6024, ZN => n6020);
   U7406 : AOI221_X1 port map( B1 => n13854, B2 => n8113, C1 => n13851, C2 => 
                           n8081, A => n6025, ZN => n6024);
   U7407 : AOI221_X1 port map( B1 => n13812, B2 => n1893, C1 => n13809, C2 => 
                           n869, A => n6028, ZN => n6021);
   U7408 : AOI221_X1 port map( B1 => n13839, B2 => n1869, C1 => n13836, C2 => 
                           n868, A => n6026, ZN => n6023);
   U7409 : NAND4_X1 port map( A1 => n6058, A2 => n6059, A3 => n6060, A4 => 
                           n6061, ZN => n6057);
   U7410 : AOI221_X1 port map( B1 => n13812, B2 => n803, C1 => n13809, C2 => 
                           n871, A => n6065, ZN => n6058);
   U7411 : AOI221_X1 port map( B1 => n13839, B2 => n812, C1 => n13836, C2 => 
                           n870, A => n6063, ZN => n6060);
   U7412 : AOI221_X1 port map( B1 => n13827, B2 => n1025, C1 => n13824, C2 => 
                           n544, A => n6064, ZN => n6059);
   U7413 : NAND4_X1 port map( A1 => n6502, A2 => n6503, A3 => n6504, A4 => 
                           n6505, ZN => n6501);
   U7414 : AOI221_X1 port map( B1 => n13853, B2 => n8100, C1 => n13850, C2 => 
                           n8068, A => n6506, ZN => n6505);
   U7415 : AOI221_X1 port map( B1 => n13811, B2 => n1880, C1 => n13808, C2 => 
                           n895, A => n6520, ZN => n6502);
   U7416 : AOI221_X1 port map( B1 => n13838, B2 => n1856, C1 => n13835, C2 => 
                           n894, A => n6514, ZN => n6504);
   U7417 : NAND4_X1 port map( A1 => n4959, A2 => n4960, A3 => n4961, A4 => 
                           n4962, ZN => n4958);
   U7418 : AOI221_X1 port map( B1 => n14073, B2 => n8106, C1 => n14070, C2 => 
                           n8074, A => n4963, ZN => n4962);
   U7419 : AOI221_X1 port map( B1 => n14031, B2 => n7914, C1 => n14028, C2 => 
                           n7834, A => n4966, ZN => n4959);
   U7420 : AOI221_X1 port map( B1 => n14058, B2 => n8042, C1 => n14055, C2 => 
                           n8010, A => n4964, ZN => n4961);
   U7421 : NAND4_X1 port map( A1 => n4996, A2 => n4997, A3 => n4998, A4 => 
                           n4999, ZN => n4995);
   U7422 : AOI221_X1 port map( B1 => n14073, B2 => n8105, C1 => n14070, C2 => 
                           n8073, A => n5000, ZN => n4999);
   U7423 : AOI221_X1 port map( B1 => n14031, B2 => n7913, C1 => n14028, C2 => 
                           n7831, A => n5003, ZN => n4996);
   U7424 : AOI221_X1 port map( B1 => n14058, B2 => n8041, C1 => n14055, C2 => 
                           n8009, A => n5001, ZN => n4998);
   U7425 : NAND4_X1 port map( A1 => n5033, A2 => n5034, A3 => n5035, A4 => 
                           n5036, ZN => n5032);
   U7426 : AOI221_X1 port map( B1 => n14073, B2 => n8104, C1 => n14070, C2 => 
                           n8072, A => n5037, ZN => n5036);
   U7427 : AOI221_X1 port map( B1 => n14031, B2 => n7912, C1 => n14028, C2 => 
                           n7828, A => n5040, ZN => n5033);
   U7428 : AOI221_X1 port map( B1 => n14058, B2 => n8040, C1 => n14055, C2 => 
                           n8008, A => n5038, ZN => n5035);
   U7429 : NAND4_X1 port map( A1 => n5070, A2 => n5071, A3 => n5072, A4 => 
                           n5073, ZN => n5069);
   U7430 : AOI221_X1 port map( B1 => n14073, B2 => n8103, C1 => n14070, C2 => 
                           n8071, A => n5074, ZN => n5073);
   U7431 : AOI221_X1 port map( B1 => n14031, B2 => n7911, C1 => n14028, C2 => 
                           n7825, A => n5077, ZN => n5070);
   U7432 : AOI221_X1 port map( B1 => n14058, B2 => n8039, C1 => n14055, C2 => 
                           n8007, A => n5075, ZN => n5072);
   U7433 : NAND4_X1 port map( A1 => n5107, A2 => n5108, A3 => n5109, A4 => 
                           n5110, ZN => n5106);
   U7434 : AOI221_X1 port map( B1 => n14073, B2 => n8102, C1 => n14070, C2 => 
                           n8070, A => n5111, ZN => n5110);
   U7435 : AOI221_X1 port map( B1 => n14031, B2 => n7910, C1 => n14028, C2 => 
                           n7822, A => n5114, ZN => n5107);
   U7436 : AOI221_X1 port map( B1 => n14058, B2 => n8038, C1 => n14055, C2 => 
                           n8006, A => n5112, ZN => n5109);
   U7437 : NAND4_X1 port map( A1 => n5144, A2 => n5145, A3 => n5146, A4 => 
                           n5147, ZN => n5143);
   U7438 : AOI221_X1 port map( B1 => n14073, B2 => n8101, C1 => n14070, C2 => 
                           n8069, A => n5148, ZN => n5147);
   U7439 : AOI221_X1 port map( B1 => n14031, B2 => n7909, C1 => n14028, C2 => 
                           n7819, A => n5151, ZN => n5144);
   U7440 : AOI221_X1 port map( B1 => n14058, B2 => n8037, C1 => n14055, C2 => 
                           n8005, A => n5149, ZN => n5146);
   U7441 : NAND4_X1 port map( A1 => n3962, A2 => n3963, A3 => n3964, A4 => 
                           n3965, ZN => n3961);
   U7442 : AOI221_X1 port map( B1 => n14075, B2 => n8131, C1 => n14072, C2 => 
                           n8099, A => n3968, ZN => n3965);
   U7443 : AOI221_X1 port map( B1 => n14033, B2 => n7939, C1 => n14030, C2 => 
                           n7907, A => n3985, ZN => n3962);
   U7444 : AOI221_X1 port map( B1 => n14060, B2 => n8067, C1 => n14057, C2 => 
                           n8035, A => n3974, ZN => n3964);
   U7445 : NAND4_X1 port map( A1 => n5283, A2 => n5284, A3 => n5285, A4 => 
                           n5286, ZN => n5282);
   U7446 : AOI221_X1 port map( B1 => n13855, B2 => n8131, C1 => n13852, C2 => 
                           n8099, A => n5289, ZN => n5286);
   U7447 : AOI221_X1 port map( B1 => n13813, B2 => n1830, C1 => n13810, C2 => 
                           n833, A => n5306, ZN => n5283);
   U7448 : AOI221_X1 port map( B1 => n13840, B2 => n1822, C1 => n13837, C2 => 
                           n832, A => n5295, ZN => n5285);
   U7449 : NAND4_X1 port map( A1 => n6564, A2 => n6565, A3 => n6566, A4 => 
                           n6567, ZN => n6563);
   U7450 : AOI221_X1 port map( B1 => n14228, B2 => n2494, C1 => n14227, C2 => 
                           n1716, A => n6575, ZN => n6564);
   U7451 : AOI221_X1 port map( B1 => n8767, B2 => n14255, C1 => n8735, C2 => 
                           n14252, A => n6570, ZN => n6566);
   U7452 : AOI221_X1 port map( B1 => n14243, B2 => n1724, C1 => n7113, C2 => 
                           n14240, A => n6571, ZN => n6565);
   U7453 : NAND4_X1 port map( A1 => n4069, A2 => n4070, A3 => n4071, A4 => 
                           n4072, ZN => n4068);
   U7454 : AOI221_X1 port map( B1 => n14033, B2 => n7938, C1 => n14030, C2 => 
                           n7906, A => n4076, ZN => n4069);
   U7455 : AOI221_X1 port map( B1 => n14060, B2 => n8066, C1 => n14057, C2 => 
                           n8034, A => n4074, ZN => n4071);
   U7456 : AOI221_X1 port map( B1 => n14048, B2 => n8002, C1 => n14045, C2 => 
                           n7970, A => n4075, ZN => n4070);
   U7457 : NAND4_X1 port map( A1 => n2783, A2 => n2784, A3 => n2785, A4 => 
                           n2786, ZN => n2782);
   U7458 : AOI221_X1 port map( B1 => n14229, B2 => n2493, C1 => n899, C2 => 
                           n14226, A => n2806, ZN => n2783);
   U7459 : AOI221_X1 port map( B1 => n8766, B2 => n14257, C1 => n8734, C2 => 
                           n14254, A => n2795, ZN => n2785);
   U7460 : AOI221_X1 port map( B1 => n14244, B2 => n1723, C1 => n7114, C2 => 
                           n14241, A => n2800, ZN => n2784);
   U7461 : NAND4_X1 port map( A1 => n4108, A2 => n4109, A3 => n4110, A4 => 
                           n4111, ZN => n4107);
   U7462 : AOI221_X1 port map( B1 => n14033, B2 => n7937, C1 => n14030, C2 => 
                           n7903, A => n4115, ZN => n4108);
   U7463 : AOI221_X1 port map( B1 => n14060, B2 => n8065, C1 => n14057, C2 => 
                           n8033, A => n4113, ZN => n4110);
   U7464 : AOI221_X1 port map( B1 => n14048, B2 => n8001, C1 => n14045, C2 => 
                           n7969, A => n4114, ZN => n4109);
   U7465 : NAND4_X1 port map( A1 => n5429, A2 => n5430, A3 => n5431, A4 => 
                           n5432, ZN => n5428);
   U7466 : AOI221_X1 port map( B1 => n13813, B2 => n1828, C1 => n13810, C2 => 
                           n837, A => n5436, ZN => n5429);
   U7467 : AOI221_X1 port map( B1 => n13840, B2 => n1820, C1 => n13837, C2 => 
                           n836, A => n5434, ZN => n5431);
   U7468 : AOI221_X1 port map( B1 => n13828, B2 => n8001, C1 => n13825, C2 => 
                           n7969, A => n5435, ZN => n5430);
   U7469 : NAND4_X1 port map( A1 => n2883, A2 => n2884, A3 => n2885, A4 => 
                           n2886, ZN => n2882);
   U7470 : AOI221_X1 port map( B1 => n14228, B2 => n2492, C1 => n905, C2 => 
                           n14225, A => n2890, ZN => n2883);
   U7471 : AOI221_X1 port map( B1 => n8765, B2 => n14257, C1 => n8733, C2 => 
                           n14254, A => n2888, ZN => n2885);
   U7472 : AOI221_X1 port map( B1 => n14243, B2 => n1722, C1 => n7116, C2 => 
                           n14240, A => n2889, ZN => n2884);
   U7473 : NAND4_X1 port map( A1 => n4145, A2 => n4146, A3 => n4147, A4 => 
                           n4148, ZN => n4144);
   U7474 : AOI221_X1 port map( B1 => n14033, B2 => n7936, C1 => n14030, C2 => 
                           n7900, A => n4152, ZN => n4145);
   U7475 : AOI221_X1 port map( B1 => n14060, B2 => n8064, C1 => n14057, C2 => 
                           n8032, A => n4150, ZN => n4147);
   U7476 : AOI221_X1 port map( B1 => n14048, B2 => n8000, C1 => n14045, C2 => 
                           n7968, A => n4151, ZN => n4146);
   U7477 : NAND4_X1 port map( A1 => n2920, A2 => n2921, A3 => n2922, A4 => 
                           n2923, ZN => n2919);
   U7478 : AOI221_X1 port map( B1 => n14228, B2 => n2491, C1 => n911, C2 => 
                           n14225, A => n2927, ZN => n2920);
   U7479 : AOI221_X1 port map( B1 => n8764, B2 => n14257, C1 => n8732, C2 => 
                           n14254, A => n2925, ZN => n2922);
   U7480 : AOI221_X1 port map( B1 => n14243, B2 => n1721, C1 => n7117, C2 => 
                           n14240, A => n2926, ZN => n2921);
   U7481 : NAND4_X1 port map( A1 => n4182, A2 => n4183, A3 => n4184, A4 => 
                           n4185, ZN => n4181);
   U7482 : AOI221_X1 port map( B1 => n14033, B2 => n7935, C1 => n14030, C2 => 
                           n7897, A => n4189, ZN => n4182);
   U7483 : AOI221_X1 port map( B1 => n14060, B2 => n8063, C1 => n14057, C2 => 
                           n8031, A => n4187, ZN => n4184);
   U7484 : AOI221_X1 port map( B1 => n14048, B2 => n7999, C1 => n14045, C2 => 
                           n7967, A => n4188, ZN => n4183);
   U7485 : NAND4_X1 port map( A1 => n2957, A2 => n2958, A3 => n2959, A4 => 
                           n2960, ZN => n2956);
   U7486 : AOI221_X1 port map( B1 => n14228, B2 => n2490, C1 => n917, C2 => 
                           n14225, A => n2964, ZN => n2957);
   U7487 : AOI221_X1 port map( B1 => n8763, B2 => n14257, C1 => n8731, C2 => 
                           n14254, A => n2962, ZN => n2959);
   U7488 : AOI221_X1 port map( B1 => n14243, B2 => n1720, C1 => n7119, C2 => 
                           n14240, A => n2963, ZN => n2958);
   U7489 : NAND4_X1 port map( A1 => n4219, A2 => n4220, A3 => n4221, A4 => 
                           n4222, ZN => n4218);
   U7490 : AOI221_X1 port map( B1 => n14033, B2 => n7934, C1 => n14030, C2 => 
                           n7894, A => n4226, ZN => n4219);
   U7491 : AOI221_X1 port map( B1 => n14060, B2 => n8062, C1 => n14057, C2 => 
                           n8030, A => n4224, ZN => n4221);
   U7492 : AOI221_X1 port map( B1 => n14048, B2 => n7998, C1 => n14045, C2 => 
                           n7966, A => n4225, ZN => n4220);
   U7493 : NAND4_X1 port map( A1 => n2994, A2 => n2995, A3 => n2996, A4 => 
                           n2997, ZN => n2993);
   U7494 : AOI221_X1 port map( B1 => n14228, B2 => n2489, C1 => n923, C2 => 
                           n14225, A => n3001, ZN => n2994);
   U7495 : AOI221_X1 port map( B1 => n8762, B2 => n14257, C1 => n8730, C2 => 
                           n14254, A => n2999, ZN => n2996);
   U7496 : AOI221_X1 port map( B1 => n14243, B2 => n1719, C1 => n7120, C2 => 
                           n14240, A => n3000, ZN => n2995);
   U7497 : NAND4_X1 port map( A1 => n3031, A2 => n3032, A3 => n3033, A4 => 
                           n3034, ZN => n3030);
   U7498 : AOI221_X1 port map( B1 => n14228, B2 => n2488, C1 => n929, C2 => 
                           n14225, A => n3038, ZN => n3031);
   U7499 : AOI221_X1 port map( B1 => n8761, B2 => n14257, C1 => n8729, C2 => 
                           n14254, A => n3036, ZN => n3033);
   U7500 : AOI221_X1 port map( B1 => n14243, B2 => n1718, C1 => n7122, C2 => 
                           n14240, A => n3037, ZN => n3032);
   U7501 : NAND4_X1 port map( A1 => n4293, A2 => n4294, A3 => n4295, A4 => 
                           n4296, ZN => n4292);
   U7502 : AOI221_X1 port map( B1 => n14033, B2 => n7932, C1 => n14030, C2 => 
                           n7888, A => n4300, ZN => n4293);
   U7503 : AOI221_X1 port map( B1 => n14060, B2 => n8060, C1 => n14057, C2 => 
                           n8028, A => n4298, ZN => n4295);
   U7504 : AOI221_X1 port map( B1 => n14048, B2 => n7996, C1 => n14045, C2 => 
                           n7964, A => n4299, ZN => n4294);
   U7505 : NAND4_X1 port map( A1 => n5614, A2 => n5615, A3 => n5616, A4 => 
                           n5617, ZN => n5613);
   U7506 : AOI221_X1 port map( B1 => n13813, B2 => n1823, C1 => n13810, C2 => 
                           n847, A => n5621, ZN => n5614);
   U7507 : AOI221_X1 port map( B1 => n13840, B2 => n1815, C1 => n13837, C2 => 
                           n846, A => n5619, ZN => n5616);
   U7508 : AOI221_X1 port map( B1 => n13828, B2 => n7996, C1 => n13825, C2 => 
                           n7964, A => n5620, ZN => n5615);
   U7509 : NAND4_X1 port map( A1 => n3068, A2 => n3069, A3 => n3070, A4 => 
                           n3071, ZN => n3067);
   U7510 : AOI221_X1 port map( B1 => n14228, B2 => n2487, C1 => n935, C2 => 
                           n14225, A => n3075, ZN => n3068);
   U7511 : AOI221_X1 port map( B1 => n8760, B2 => n14257, C1 => n8728, C2 => 
                           n14254, A => n3073, ZN => n3070);
   U7512 : AOI221_X1 port map( B1 => n14243, B2 => n1717, C1 => n7123, C2 => 
                           n14240, A => n3074, ZN => n3069);
   U7513 : NAND4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => 
                           n4333, ZN => n4329);
   U7514 : AOI221_X1 port map( B1 => n14032, B2 => n7931, C1 => n14029, C2 => 
                           n7885, A => n4337, ZN => n4330);
   U7515 : AOI221_X1 port map( B1 => n14059, B2 => n8059, C1 => n14056, C2 => 
                           n8027, A => n4335, ZN => n4332);
   U7516 : AOI221_X1 port map( B1 => n14047, B2 => n7995, C1 => n14044, C2 => 
                           n7963, A => n4336, ZN => n4331);
   U7517 : NAND4_X1 port map( A1 => n5651, A2 => n5652, A3 => n5653, A4 => 
                           n5654, ZN => n5650);
   U7518 : AOI221_X1 port map( B1 => n13812, B2 => n1903, C1 => n13809, C2 => 
                           n849, A => n5658, ZN => n5651);
   U7519 : AOI221_X1 port map( B1 => n13839, B2 => n1879, C1 => n13836, C2 => 
                           n848, A => n5656, ZN => n5653);
   U7520 : AOI221_X1 port map( B1 => n13827, B2 => n7995, C1 => n13824, C2 => 
                           n7963, A => n5657, ZN => n5652);
   U7521 : NAND4_X1 port map( A1 => n3105, A2 => n3106, A3 => n3107, A4 => 
                           n3108, ZN => n3104);
   U7522 : AOI221_X1 port map( B1 => n14228, B2 => n2518, C1 => n941, C2 => 
                           n14225, A => n3112, ZN => n3105);
   U7523 : AOI221_X1 port map( B1 => n8759, B2 => n14257, C1 => n8727, C2 => 
                           n14254, A => n3110, ZN => n3107);
   U7524 : AOI221_X1 port map( B1 => n14243, B2 => n1941, C1 => n7125, C2 => 
                           n14240, A => n3111, ZN => n3106);
   U7525 : NAND4_X1 port map( A1 => n4367, A2 => n4368, A3 => n4369, A4 => 
                           n4370, ZN => n4366);
   U7526 : AOI221_X1 port map( B1 => n14032, B2 => n7930, C1 => n14029, C2 => 
                           n7882, A => n4374, ZN => n4367);
   U7527 : AOI221_X1 port map( B1 => n14059, B2 => n8058, C1 => n14056, C2 => 
                           n8026, A => n4372, ZN => n4369);
   U7528 : AOI221_X1 port map( B1 => n14047, B2 => n7994, C1 => n14044, C2 => 
                           n7962, A => n4373, ZN => n4368);
   U7529 : NAND4_X1 port map( A1 => n5688, A2 => n5689, A3 => n5690, A4 => 
                           n5691, ZN => n5687);
   U7530 : AOI221_X1 port map( B1 => n13812, B2 => n1902, C1 => n13809, C2 => 
                           n851, A => n5695, ZN => n5688);
   U7531 : AOI221_X1 port map( B1 => n13839, B2 => n1878, C1 => n13836, C2 => 
                           n850, A => n5693, ZN => n5690);
   U7532 : AOI221_X1 port map( B1 => n13827, B2 => n7994, C1 => n13824, C2 => 
                           n7962, A => n5694, ZN => n5689);
   U7533 : NAND4_X1 port map( A1 => n3142, A2 => n3143, A3 => n3144, A4 => 
                           n3145, ZN => n3141);
   U7534 : AOI221_X1 port map( B1 => n14228, B2 => n2517, C1 => n947, C2 => 
                           n14225, A => n3149, ZN => n3142);
   U7535 : AOI221_X1 port map( B1 => n8758, B2 => n14256, C1 => n8726, C2 => 
                           n14253, A => n3147, ZN => n3144);
   U7536 : AOI221_X1 port map( B1 => n14243, B2 => n1940, C1 => n7128, C2 => 
                           n14240, A => n3148, ZN => n3143);
   U7537 : NAND4_X1 port map( A1 => n4404, A2 => n4405, A3 => n4406, A4 => 
                           n4407, ZN => n4403);
   U7538 : AOI221_X1 port map( B1 => n14032, B2 => n7929, C1 => n14029, C2 => 
                           n7879, A => n4411, ZN => n4404);
   U7539 : AOI221_X1 port map( B1 => n14059, B2 => n8057, C1 => n14056, C2 => 
                           n8025, A => n4409, ZN => n4406);
   U7540 : AOI221_X1 port map( B1 => n14047, B2 => n7993, C1 => n14044, C2 => 
                           n7961, A => n4410, ZN => n4405);
   U7541 : NAND4_X1 port map( A1 => n5725, A2 => n5726, A3 => n5727, A4 => 
                           n5728, ZN => n5724);
   U7542 : AOI221_X1 port map( B1 => n13812, B2 => n1901, C1 => n13809, C2 => 
                           n853, A => n5732, ZN => n5725);
   U7543 : AOI221_X1 port map( B1 => n13839, B2 => n1877, C1 => n13836, C2 => 
                           n852, A => n5730, ZN => n5727);
   U7544 : AOI221_X1 port map( B1 => n13827, B2 => n7993, C1 => n13824, C2 => 
                           n7961, A => n5731, ZN => n5726);
   U7545 : NAND4_X1 port map( A1 => n3179, A2 => n3180, A3 => n3181, A4 => 
                           n3182, ZN => n3178);
   U7546 : AOI221_X1 port map( B1 => n14228, B2 => n2516, C1 => n953, C2 => 
                           n14225, A => n3186, ZN => n3179);
   U7547 : AOI221_X1 port map( B1 => n8757, B2 => n14256, C1 => n8725, C2 => 
                           n14253, A => n3184, ZN => n3181);
   U7548 : AOI221_X1 port map( B1 => n14243, B2 => n1939, C1 => n7129, C2 => 
                           n14240, A => n3185, ZN => n3180);
   U7549 : NAND4_X1 port map( A1 => n4441, A2 => n4442, A3 => n4443, A4 => 
                           n4444, ZN => n4440);
   U7550 : AOI221_X1 port map( B1 => n14032, B2 => n7928, C1 => n14029, C2 => 
                           n7876, A => n4448, ZN => n4441);
   U7551 : AOI221_X1 port map( B1 => n14059, B2 => n8056, C1 => n14056, C2 => 
                           n8024, A => n4446, ZN => n4443);
   U7552 : AOI221_X1 port map( B1 => n14047, B2 => n7992, C1 => n14044, C2 => 
                           n7960, A => n4447, ZN => n4442);
   U7553 : NAND4_X1 port map( A1 => n5762, A2 => n5763, A3 => n5764, A4 => 
                           n5765, ZN => n5761);
   U7554 : AOI221_X1 port map( B1 => n13812, B2 => n1900, C1 => n13809, C2 => 
                           n855, A => n5769, ZN => n5762);
   U7555 : AOI221_X1 port map( B1 => n13839, B2 => n1876, C1 => n13836, C2 => 
                           n854, A => n5767, ZN => n5764);
   U7556 : AOI221_X1 port map( B1 => n13827, B2 => n7992, C1 => n13824, C2 => 
                           n7960, A => n5768, ZN => n5763);
   U7557 : NAND4_X1 port map( A1 => n3216, A2 => n3217, A3 => n3218, A4 => 
                           n3219, ZN => n3215);
   U7558 : AOI221_X1 port map( B1 => n14228, B2 => n2515, C1 => n959, C2 => 
                           n14225, A => n3223, ZN => n3216);
   U7559 : AOI221_X1 port map( B1 => n8756, B2 => n14256, C1 => n8724, C2 => 
                           n14253, A => n3221, ZN => n3218);
   U7560 : AOI221_X1 port map( B1 => n14243, B2 => n1938, C1 => n7131, C2 => 
                           n14240, A => n3222, ZN => n3217);
   U7561 : NAND4_X1 port map( A1 => n4478, A2 => n4479, A3 => n4480, A4 => 
                           n4481, ZN => n4477);
   U7562 : AOI221_X1 port map( B1 => n14032, B2 => n7927, C1 => n14029, C2 => 
                           n7873, A => n4485, ZN => n4478);
   U7563 : AOI221_X1 port map( B1 => n14059, B2 => n8055, C1 => n14056, C2 => 
                           n8023, A => n4483, ZN => n4480);
   U7564 : AOI221_X1 port map( B1 => n14047, B2 => n7991, C1 => n14044, C2 => 
                           n7959, A => n4484, ZN => n4479);
   U7565 : NAND4_X1 port map( A1 => n5799, A2 => n5800, A3 => n5801, A4 => 
                           n5802, ZN => n5798);
   U7566 : AOI221_X1 port map( B1 => n13812, B2 => n1899, C1 => n13809, C2 => 
                           n857, A => n5806, ZN => n5799);
   U7567 : AOI221_X1 port map( B1 => n13839, B2 => n1875, C1 => n13836, C2 => 
                           n856, A => n5804, ZN => n5801);
   U7568 : AOI221_X1 port map( B1 => n13827, B2 => n7991, C1 => n13824, C2 => 
                           n7959, A => n5805, ZN => n5800);
   U7569 : NAND4_X1 port map( A1 => n3253, A2 => n3254, A3 => n3255, A4 => 
                           n3256, ZN => n3252);
   U7570 : AOI221_X1 port map( B1 => n14228, B2 => n2514, C1 => n965, C2 => 
                           n14225, A => n3260, ZN => n3253);
   U7571 : AOI221_X1 port map( B1 => n8755, B2 => n14256, C1 => n8723, C2 => 
                           n14253, A => n3258, ZN => n3255);
   U7572 : AOI221_X1 port map( B1 => n14243, B2 => n1937, C1 => n7132, C2 => 
                           n14240, A => n3259, ZN => n3254);
   U7573 : NAND4_X1 port map( A1 => n4515, A2 => n4516, A3 => n4517, A4 => 
                           n4518, ZN => n4514);
   U7574 : AOI221_X1 port map( B1 => n14032, B2 => n7926, C1 => n14029, C2 => 
                           n7870, A => n4522, ZN => n4515);
   U7575 : AOI221_X1 port map( B1 => n14059, B2 => n8054, C1 => n14056, C2 => 
                           n8022, A => n4520, ZN => n4517);
   U7576 : AOI221_X1 port map( B1 => n14047, B2 => n7990, C1 => n14044, C2 => 
                           n7958, A => n4521, ZN => n4516);
   U7577 : NAND4_X1 port map( A1 => n5836, A2 => n5837, A3 => n5838, A4 => 
                           n5839, ZN => n5835);
   U7578 : AOI221_X1 port map( B1 => n13812, B2 => n1898, C1 => n13809, C2 => 
                           n859, A => n5843, ZN => n5836);
   U7579 : AOI221_X1 port map( B1 => n13839, B2 => n1874, C1 => n13836, C2 => 
                           n858, A => n5841, ZN => n5838);
   U7580 : AOI221_X1 port map( B1 => n13827, B2 => n7990, C1 => n13824, C2 => 
                           n7958, A => n5842, ZN => n5837);
   U7581 : NAND4_X1 port map( A1 => n3290, A2 => n3291, A3 => n3292, A4 => 
                           n3293, ZN => n3289);
   U7582 : AOI221_X1 port map( B1 => n14229, B2 => n2513, C1 => n971, C2 => 
                           n14225, A => n3297, ZN => n3290);
   U7583 : AOI221_X1 port map( B1 => n8754, B2 => n14256, C1 => n8722, C2 => 
                           n14253, A => n3295, ZN => n3292);
   U7584 : AOI221_X1 port map( B1 => n14244, B2 => n1936, C1 => n7133, C2 => 
                           n14241, A => n3296, ZN => n3291);
   U7585 : NAND4_X1 port map( A1 => n4552, A2 => n4553, A3 => n4554, A4 => 
                           n4555, ZN => n4551);
   U7586 : AOI221_X1 port map( B1 => n14032, B2 => n7925, C1 => n14029, C2 => 
                           n7867, A => n4559, ZN => n4552);
   U7587 : AOI221_X1 port map( B1 => n14059, B2 => n8053, C1 => n14056, C2 => 
                           n8021, A => n4557, ZN => n4554);
   U7588 : AOI221_X1 port map( B1 => n14047, B2 => n7989, C1 => n14044, C2 => 
                           n7957, A => n4558, ZN => n4553);
   U7589 : NAND4_X1 port map( A1 => n5873, A2 => n5874, A3 => n5875, A4 => 
                           n5876, ZN => n5872);
   U7590 : AOI221_X1 port map( B1 => n13812, B2 => n1897, C1 => n13809, C2 => 
                           n861, A => n5880, ZN => n5873);
   U7591 : AOI221_X1 port map( B1 => n13839, B2 => n1873, C1 => n13836, C2 => 
                           n860, A => n5878, ZN => n5875);
   U7592 : AOI221_X1 port map( B1 => n13827, B2 => n7989, C1 => n13824, C2 => 
                           n7957, A => n5879, ZN => n5874);
   U7593 : NAND4_X1 port map( A1 => n3329, A2 => n3330, A3 => n3331, A4 => 
                           n3332, ZN => n3328);
   U7594 : AOI221_X1 port map( B1 => n14229, B2 => n2512, C1 => n977, C2 => 
                           n14226, A => n3336, ZN => n3329);
   U7595 : AOI221_X1 port map( B1 => n8753, B2 => n14256, C1 => n8721, C2 => 
                           n14253, A => n3334, ZN => n3331);
   U7596 : AOI221_X1 port map( B1 => n14244, B2 => n1935, C1 => n7135, C2 => 
                           n14241, A => n3335, ZN => n3330);
   U7597 : NAND4_X1 port map( A1 => n4589, A2 => n4590, A3 => n4591, A4 => 
                           n4592, ZN => n4588);
   U7598 : AOI221_X1 port map( B1 => n14032, B2 => n7924, C1 => n14029, C2 => 
                           n7864, A => n4596, ZN => n4589);
   U7599 : AOI221_X1 port map( B1 => n14059, B2 => n8052, C1 => n14056, C2 => 
                           n8020, A => n4594, ZN => n4591);
   U7600 : AOI221_X1 port map( B1 => n14047, B2 => n7988, C1 => n14044, C2 => 
                           n7956, A => n4595, ZN => n4590);
   U7601 : NAND4_X1 port map( A1 => n5910, A2 => n5911, A3 => n5912, A4 => 
                           n5913, ZN => n5909);
   U7602 : AOI221_X1 port map( B1 => n13812, B2 => n1896, C1 => n13809, C2 => 
                           n863, A => n5917, ZN => n5910);
   U7603 : AOI221_X1 port map( B1 => n13839, B2 => n1872, C1 => n13836, C2 => 
                           n862, A => n5915, ZN => n5912);
   U7604 : AOI221_X1 port map( B1 => n13827, B2 => n7988, C1 => n13824, C2 => 
                           n7956, A => n5916, ZN => n5911);
   U7605 : NAND4_X1 port map( A1 => n3366, A2 => n3367, A3 => n3368, A4 => 
                           n3369, ZN => n3365);
   U7606 : AOI221_X1 port map( B1 => n14229, B2 => n2511, C1 => n983, C2 => 
                           n14226, A => n3373, ZN => n3366);
   U7607 : AOI221_X1 port map( B1 => n8752, B2 => n14256, C1 => n8720, C2 => 
                           n14253, A => n3371, ZN => n3368);
   U7608 : AOI221_X1 port map( B1 => n14244, B2 => n1934, C1 => n7137, C2 => 
                           n14241, A => n3372, ZN => n3367);
   U7609 : NAND4_X1 port map( A1 => n4626, A2 => n4627, A3 => n4628, A4 => 
                           n4629, ZN => n4625);
   U7610 : AOI221_X1 port map( B1 => n14032, B2 => n7923, C1 => n14029, C2 => 
                           n7861, A => n4633, ZN => n4626);
   U7611 : AOI221_X1 port map( B1 => n14059, B2 => n8051, C1 => n14056, C2 => 
                           n8019, A => n4631, ZN => n4628);
   U7612 : AOI221_X1 port map( B1 => n14047, B2 => n7987, C1 => n14044, C2 => 
                           n7955, A => n4632, ZN => n4627);
   U7613 : NAND4_X1 port map( A1 => n5947, A2 => n5948, A3 => n5949, A4 => 
                           n5950, ZN => n5946);
   U7614 : AOI221_X1 port map( B1 => n13812, B2 => n1895, C1 => n13809, C2 => 
                           n865, A => n5954, ZN => n5947);
   U7615 : AOI221_X1 port map( B1 => n13839, B2 => n1871, C1 => n13836, C2 => 
                           n864, A => n5952, ZN => n5949);
   U7616 : AOI221_X1 port map( B1 => n13827, B2 => n7987, C1 => n13824, C2 => 
                           n7955, A => n5953, ZN => n5948);
   U7617 : NAND4_X1 port map( A1 => n3403, A2 => n3404, A3 => n3405, A4 => 
                           n3406, ZN => n3402);
   U7618 : AOI221_X1 port map( B1 => n14229, B2 => n2510, C1 => n989, C2 => 
                           n14226, A => n3410, ZN => n3403);
   U7619 : AOI221_X1 port map( B1 => n8751, B2 => n14256, C1 => n8719, C2 => 
                           n14253, A => n3408, ZN => n3405);
   U7620 : AOI221_X1 port map( B1 => n14244, B2 => n1933, C1 => n7138, C2 => 
                           n14241, A => n3409, ZN => n3404);
   U7621 : NAND4_X1 port map( A1 => n4663, A2 => n4664, A3 => n4665, A4 => 
                           n4666, ZN => n4662);
   U7622 : AOI221_X1 port map( B1 => n14032, B2 => n7922, C1 => n14029, C2 => 
                           n7858, A => n4670, ZN => n4663);
   U7623 : AOI221_X1 port map( B1 => n14059, B2 => n8050, C1 => n14056, C2 => 
                           n8018, A => n4668, ZN => n4665);
   U7624 : AOI221_X1 port map( B1 => n14047, B2 => n7986, C1 => n14044, C2 => 
                           n7954, A => n4669, ZN => n4664);
   U7625 : NAND4_X1 port map( A1 => n5984, A2 => n5985, A3 => n5986, A4 => 
                           n5987, ZN => n5983);
   U7626 : AOI221_X1 port map( B1 => n13812, B2 => n1894, C1 => n13809, C2 => 
                           n867, A => n5991, ZN => n5984);
   U7627 : AOI221_X1 port map( B1 => n13839, B2 => n1870, C1 => n13836, C2 => 
                           n866, A => n5989, ZN => n5986);
   U7628 : AOI221_X1 port map( B1 => n13827, B2 => n7986, C1 => n13824, C2 => 
                           n7954, A => n5990, ZN => n5985);
   U7629 : NAND4_X1 port map( A1 => n3440, A2 => n3441, A3 => n3442, A4 => 
                           n3443, ZN => n3439);
   U7630 : AOI221_X1 port map( B1 => n14229, B2 => n2509, C1 => n995, C2 => 
                           n14226, A => n3447, ZN => n3440);
   U7631 : AOI221_X1 port map( B1 => n8750, B2 => n14256, C1 => n8718, C2 => 
                           n14253, A => n3445, ZN => n3442);
   U7632 : AOI221_X1 port map( B1 => n14244, B2 => n1932, C1 => n7140, C2 => 
                           n14241, A => n3446, ZN => n3441);
   U7633 : NAND4_X1 port map( A1 => n3477, A2 => n3478, A3 => n3479, A4 => 
                           n3480, ZN => n3476);
   U7634 : AOI221_X1 port map( B1 => n14229, B2 => n2508, C1 => n14226, C2 => 
                           n1917, A => n3484, ZN => n3477);
   U7635 : AOI221_X1 port map( B1 => n8749, B2 => n14256, C1 => n8717, C2 => 
                           n14253, A => n3482, ZN => n3479);
   U7636 : AOI221_X1 port map( B1 => n14244, B2 => n1931, C1 => n7141, C2 => 
                           n14241, A => n3483, ZN => n3478);
   U7637 : NAND4_X1 port map( A1 => n3514, A2 => n3515, A3 => n3516, A4 => 
                           n3517, ZN => n3513);
   U7638 : AOI221_X1 port map( B1 => n14229, B2 => n2507, C1 => n14226, C2 => 
                           n1916, A => n3521, ZN => n3514);
   U7639 : AOI221_X1 port map( B1 => n8748, B2 => n14256, C1 => n8716, C2 => 
                           n14253, A => n3519, ZN => n3516);
   U7640 : AOI221_X1 port map( B1 => n14244, B2 => n1930, C1 => n7143, C2 => 
                           n14241, A => n3520, ZN => n3515);
   U7641 : NAND4_X1 port map( A1 => n3625, A2 => n3626, A3 => n3627, A4 => 
                           n3628, ZN => n3624);
   U7642 : AOI221_X1 port map( B1 => n14229, B2 => n2504, C1 => n14226, C2 => 
                           n1913, A => n3632, ZN => n3625);
   U7643 : AOI221_X1 port map( B1 => n8745, B2 => n14255, C1 => n8713, C2 => 
                           n14252, A => n3630, ZN => n3627);
   U7644 : AOI221_X1 port map( B1 => n14244, B2 => n1927, C1 => n7153, C2 => 
                           n14241, A => n3631, ZN => n3626);
   U7645 : NAND4_X1 port map( A1 => n3662, A2 => n3663, A3 => n3664, A4 => 
                           n3665, ZN => n3661);
   U7646 : AOI221_X1 port map( B1 => n14229, B2 => n2503, C1 => n14226, C2 => 
                           n1912, A => n3669, ZN => n3662);
   U7647 : AOI221_X1 port map( B1 => n8744, B2 => n14255, C1 => n8712, C2 => 
                           n14252, A => n3667, ZN => n3664);
   U7648 : AOI221_X1 port map( B1 => n14244, B2 => n1926, C1 => n7155, C2 => 
                           n14241, A => n3668, ZN => n3663);
   U7649 : NAND4_X1 port map( A1 => n3699, A2 => n3700, A3 => n3701, A4 => 
                           n3702, ZN => n3698);
   U7650 : AOI221_X1 port map( B1 => n14229, B2 => n2502, C1 => n14226, C2 => 
                           n1911, A => n3706, ZN => n3699);
   U7651 : AOI221_X1 port map( B1 => n8743, B2 => n14255, C1 => n8711, C2 => 
                           n14252, A => n3704, ZN => n3701);
   U7652 : AOI221_X1 port map( B1 => n14244, B2 => n1925, C1 => n7156, C2 => 
                           n14241, A => n3705, ZN => n3700);
   U7653 : NAND4_X1 port map( A1 => n3736, A2 => n3737, A3 => n3738, A4 => 
                           n3739, ZN => n3735);
   U7654 : AOI221_X1 port map( B1 => n14229, B2 => n2501, C1 => n14227, C2 => 
                           n1910, A => n3743, ZN => n3736);
   U7655 : AOI221_X1 port map( B1 => n8742, B2 => n14255, C1 => n8710, C2 => 
                           n14252, A => n3741, ZN => n3738);
   U7656 : AOI221_X1 port map( B1 => n14244, B2 => n1924, C1 => n7157, C2 => 
                           n14241, A => n3742, ZN => n3737);
   U7657 : NAND4_X1 port map( A1 => n3773, A2 => n3774, A3 => n3775, A4 => 
                           n3776, ZN => n3772);
   U7658 : AOI221_X1 port map( B1 => n14230, B2 => n2500, C1 => n14227, C2 => 
                           n1909, A => n3780, ZN => n3773);
   U7659 : AOI221_X1 port map( B1 => n8741, B2 => n14255, C1 => n8709, C2 => 
                           n14252, A => n3778, ZN => n3775);
   U7660 : AOI221_X1 port map( B1 => n14245, B2 => n1923, C1 => n7179, C2 => 
                           n14242, A => n3779, ZN => n3774);
   U7661 : NAND4_X1 port map( A1 => n3810, A2 => n3811, A3 => n3812, A4 => 
                           n3813, ZN => n3809);
   U7662 : AOI221_X1 port map( B1 => n14230, B2 => n2499, C1 => n14227, C2 => 
                           n1908, A => n3817, ZN => n3810);
   U7663 : AOI221_X1 port map( B1 => n8740, B2 => n14255, C1 => n8708, C2 => 
                           n14252, A => n3815, ZN => n3812);
   U7664 : AOI221_X1 port map( B1 => n14245, B2 => n1922, C1 => n7180, C2 => 
                           n14242, A => n3816, ZN => n3811);
   U7665 : NAND4_X1 port map( A1 => n3847, A2 => n3848, A3 => n3849, A4 => 
                           n3850, ZN => n3846);
   U7666 : AOI221_X1 port map( B1 => n14230, B2 => n2520, C1 => n14227, C2 => 
                           n1907, A => n3854, ZN => n3847);
   U7667 : AOI221_X1 port map( B1 => n8739, B2 => n14255, C1 => n8707, C2 => 
                           n14252, A => n3852, ZN => n3849);
   U7668 : AOI221_X1 port map( B1 => n14245, B2 => n1921, C1 => n7181, C2 => 
                           n14242, A => n3853, ZN => n3848);
   U7669 : NAND4_X1 port map( A1 => n3884, A2 => n3885, A3 => n3886, A4 => 
                           n3887, ZN => n3883);
   U7670 : AOI221_X1 port map( B1 => n14230, B2 => n2496, C1 => n14227, C2 => 
                           n1906, A => n3891, ZN => n3884);
   U7671 : AOI221_X1 port map( B1 => n8738, B2 => n14255, C1 => n8706, C2 => 
                           n14252, A => n3889, ZN => n3886);
   U7672 : AOI221_X1 port map( B1 => n14245, B2 => n1920, C1 => n7203, C2 => 
                           n14242, A => n3890, ZN => n3885);
   U7673 : NAND4_X1 port map( A1 => n3921, A2 => n3922, A3 => n3923, A4 => 
                           n3924, ZN => n3920);
   U7674 : AOI221_X1 port map( B1 => n14230, B2 => n2495, C1 => n14227, C2 => 
                           n1905, A => n3928, ZN => n3921);
   U7675 : AOI221_X1 port map( B1 => n8737, B2 => n14255, C1 => n8705, C2 => 
                           n14252, A => n3926, ZN => n3923);
   U7676 : AOI221_X1 port map( B1 => n14245, B2 => n1919, C1 => n7204, C2 => 
                           n14242, A => n3927, ZN => n3922);
   U7677 : NAND4_X1 port map( A1 => n5243, A2 => n5244, A3 => n5245, A4 => 
                           n5246, ZN => n5242);
   U7678 : AOI221_X1 port map( B1 => n14230, B2 => n2498, C1 => n14227, C2 => 
                           n1904, A => n5250, ZN => n5243);
   U7679 : AOI221_X1 port map( B1 => n8736, B2 => n14255, C1 => n8704, C2 => 
                           n14252, A => n5248, ZN => n5245);
   U7680 : AOI221_X1 port map( B1 => n14245, B2 => n1918, C1 => n7205, C2 => 
                           n14242, A => n5249, ZN => n5244);
   U7681 : NAND4_X1 port map( A1 => n2809, A2 => n2810, A3 => n2811, A4 => 
                           n2812, ZN => n2781);
   U7682 : AOI221_X1 port map( B1 => n8638, B2 => n14176, C1 => n8606, C2 => 
                           n14173, A => n2832, ZN => n2809);
   U7683 : AOI221_X1 port map( B1 => n8448, B2 => n14203, C1 => n8416, C2 => 
                           n14200, A => n2821, ZN => n2811);
   U7684 : AOI221_X1 port map( B1 => n14190, B2 => n1749, C1 => n8480, C2 => 
                           n14188, A => n2826, ZN => n2810);
   U7685 : NAND4_X1 port map( A1 => n2891, A2 => n2892, A3 => n2893, A4 => 
                           n2894, ZN => n2881);
   U7686 : AOI221_X1 port map( B1 => n8637, B2 => n14176, C1 => n8605, C2 => 
                           n14173, A => n2898, ZN => n2891);
   U7687 : AOI221_X1 port map( B1 => n8447, B2 => n14203, C1 => n8415, C2 => 
                           n14200, A => n2896, ZN => n2893);
   U7688 : AOI221_X1 port map( B1 => n14189, B2 => n1748, C1 => n8479, C2 => 
                           n14188, A => n2897, ZN => n2892);
   U7689 : NAND4_X1 port map( A1 => n2928, A2 => n2929, A3 => n2930, A4 => 
                           n2931, ZN => n2918);
   U7690 : AOI221_X1 port map( B1 => n8636, B2 => n14176, C1 => n8604, C2 => 
                           n14173, A => n2935, ZN => n2928);
   U7691 : AOI221_X1 port map( B1 => n8446, B2 => n14203, C1 => n8414, C2 => 
                           n14200, A => n2933, ZN => n2930);
   U7692 : AOI221_X1 port map( B1 => n14189, B2 => n1747, C1 => n8478, C2 => 
                           n14188, A => n2934, ZN => n2929);
   U7693 : NAND4_X1 port map( A1 => n2965, A2 => n2966, A3 => n2967, A4 => 
                           n2968, ZN => n2955);
   U7694 : AOI221_X1 port map( B1 => n8635, B2 => n14176, C1 => n8603, C2 => 
                           n14173, A => n2972, ZN => n2965);
   U7695 : AOI221_X1 port map( B1 => n8445, B2 => n14203, C1 => n8413, C2 => 
                           n14200, A => n2970, ZN => n2967);
   U7696 : AOI221_X1 port map( B1 => n14189, B2 => n1746, C1 => n8477, C2 => 
                           n14188, A => n2971, ZN => n2966);
   U7697 : NAND4_X1 port map( A1 => n3002, A2 => n3003, A3 => n3004, A4 => 
                           n3005, ZN => n2992);
   U7698 : AOI221_X1 port map( B1 => n8634, B2 => n14176, C1 => n8602, C2 => 
                           n14173, A => n3009, ZN => n3002);
   U7699 : AOI221_X1 port map( B1 => n8444, B2 => n14203, C1 => n8412, C2 => 
                           n14200, A => n3007, ZN => n3004);
   U7700 : AOI221_X1 port map( B1 => n14189, B2 => n1745, C1 => n8476, C2 => 
                           n14188, A => n3008, ZN => n3003);
   U7701 : NAND4_X1 port map( A1 => n3039, A2 => n3040, A3 => n3041, A4 => 
                           n3042, ZN => n3029);
   U7702 : AOI221_X1 port map( B1 => n8633, B2 => n14176, C1 => n8601, C2 => 
                           n14173, A => n3046, ZN => n3039);
   U7703 : AOI221_X1 port map( B1 => n8443, B2 => n14203, C1 => n8411, C2 => 
                           n14200, A => n3044, ZN => n3041);
   U7704 : AOI221_X1 port map( B1 => n14189, B2 => n1744, C1 => n8475, C2 => 
                           n14188, A => n3045, ZN => n3040);
   U7705 : NAND4_X1 port map( A1 => n3076, A2 => n3077, A3 => n3078, A4 => 
                           n3079, ZN => n3066);
   U7706 : AOI221_X1 port map( B1 => n8632, B2 => n14176, C1 => n8600, C2 => 
                           n14173, A => n3083, ZN => n3076);
   U7707 : AOI221_X1 port map( B1 => n8442, B2 => n14203, C1 => n8410, C2 => 
                           n14200, A => n3081, ZN => n3078);
   U7708 : AOI221_X1 port map( B1 => n14189, B2 => n1743, C1 => n8474, C2 => 
                           n14188, A => n3082, ZN => n3077);
   U7709 : NAND4_X1 port map( A1 => n3113, A2 => n3114, A3 => n3115, A4 => 
                           n3116, ZN => n3103);
   U7710 : AOI221_X1 port map( B1 => n8631, B2 => n14176, C1 => n8599, C2 => 
                           n14173, A => n3120, ZN => n3113);
   U7711 : AOI221_X1 port map( B1 => n8441, B2 => n14203, C1 => n8409, C2 => 
                           n14200, A => n3118, ZN => n3115);
   U7712 : AOI221_X1 port map( B1 => n14189, B2 => n2118, C1 => n8473, C2 => 
                           n14188, A => n3119, ZN => n3114);
   U7713 : NAND4_X1 port map( A1 => n4264, A2 => n4265, A3 => n4266, A4 => 
                           n4267, ZN => n4254);
   U7714 : AOI221_X1 port map( B1 => n13994, B2 => n8189, C1 => n13991, C2 => 
                           n8157, A => n4270, ZN => n4265);
   U7715 : AOI221_X1 port map( B1 => n13979, B2 => n1840, C1 => n13976, C2 => 
                           n1832, A => n4271, ZN => n4264);
   U7716 : AOI221_X1 port map( B1 => n14004, B2 => n1793, C1 => n14003, C2 => 
                           n1800, A => n4269, ZN => n4266);
   U7717 : NAND4_X1 port map( A1 => n5400, A2 => n5401, A3 => n5402, A4 => 
                           n5403, ZN => n5390);
   U7718 : AOI221_X1 port map( B1 => n13774, B2 => n8194, C1 => n13771, C2 => 
                           n8162, A => n5406, ZN => n5401);
   U7719 : AOI221_X1 port map( B1 => n13759, B2 => n1845, C1 => n13756, C2 => 
                           n1837, A => n5407, ZN => n5400);
   U7720 : AOI221_X1 port map( B1 => n13786, B2 => n1805, C1 => n13783, C2 => 
                           n1798, A => n5405, ZN => n5402);
   U7721 : NAND4_X1 port map( A1 => n5474, A2 => n5475, A3 => n5476, A4 => 
                           n5477, ZN => n5464);
   U7722 : AOI221_X1 port map( B1 => n13774, B2 => n8192, C1 => n13771, C2 => 
                           n8160, A => n5480, ZN => n5475);
   U7723 : AOI221_X1 port map( B1 => n13759, B2 => n1843, C1 => n13756, C2 => 
                           n1835, A => n5481, ZN => n5474);
   U7724 : AOI221_X1 port map( B1 => n13786, B2 => n1803, C1 => n13783, C2 => 
                           n1796, A => n5479, ZN => n5476);
   U7725 : NAND4_X1 port map( A1 => n5511, A2 => n5512, A3 => n5513, A4 => 
                           n5514, ZN => n5501);
   U7726 : AOI221_X1 port map( B1 => n13774, B2 => n8191, C1 => n13771, C2 => 
                           n8159, A => n5517, ZN => n5512);
   U7727 : AOI221_X1 port map( B1 => n13759, B2 => n1842, C1 => n13756, C2 => 
                           n1834, A => n5518, ZN => n5511);
   U7728 : AOI221_X1 port map( B1 => n13786, B2 => n1802, C1 => n13783, C2 => 
                           n1795, A => n5516, ZN => n5513);
   U7729 : NAND4_X1 port map( A1 => n5548, A2 => n5549, A3 => n5550, A4 => 
                           n5551, ZN => n5538);
   U7730 : AOI221_X1 port map( B1 => n13774, B2 => n8190, C1 => n13771, C2 => 
                           n8158, A => n5554, ZN => n5549);
   U7731 : AOI221_X1 port map( B1 => n13759, B2 => n1841, C1 => n13756, C2 => 
                           n1833, A => n5555, ZN => n5548);
   U7732 : AOI221_X1 port map( B1 => n13786, B2 => n1801, C1 => n13783, C2 => 
                           n1794, A => n5553, ZN => n5550);
   U7733 : NAND4_X1 port map( A1 => n5585, A2 => n5586, A3 => n5587, A4 => 
                           n5588, ZN => n5575);
   U7734 : AOI221_X1 port map( B1 => n13774, B2 => n8189, C1 => n13771, C2 => 
                           n8157, A => n5591, ZN => n5586);
   U7735 : AOI221_X1 port map( B1 => n13759, B2 => n1840, C1 => n13756, C2 => 
                           n1832, A => n5592, ZN => n5585);
   U7736 : AOI221_X1 port map( B1 => n13786, B2 => n1800, C1 => n13783, C2 => 
                           n1793, A => n5590, ZN => n5587);
   U7737 : NAND4_X1 port map( A1 => n5200, A2 => n5201, A3 => n5202, A4 => 
                           n5203, ZN => n5179);
   U7738 : AOI221_X1 port map( B1 => n13992, B2 => n8164, C1 => n13989, C2 => 
                           n8132, A => n5208, ZN => n5201);
   U7739 : AOI221_X1 port map( B1 => n13977, B2 => n2459, C1 => n13974, C2 => 
                           n2438, A => n5209, ZN => n5200);
   U7740 : AOI221_X1 port map( B1 => n897, B2 => n14006, C1 => n14001, C2 => 
                           n1965, A => n5207, ZN => n5202);
   U7741 : NAND4_X1 port map( A1 => n4782, A2 => n4783, A3 => n4784, A4 => 
                           n4785, ZN => n4772);
   U7742 : AOI221_X1 port map( B1 => n13977, B2 => n2467, C1 => n13974, C2 => 
                           n2446, A => n4789, ZN => n4782);
   U7743 : AOI221_X1 port map( B1 => n14005, B2 => n1952, C1 => n14001, C2 => 
                           n1976, A => n4787, ZN => n4784);
   U7744 : AOI221_X1 port map( B1 => n13992, B2 => n8175, C1 => n13989, C2 => 
                           n8143, A => n4788, ZN => n4783);
   U7745 : NAND4_X1 port map( A1 => n4819, A2 => n4820, A3 => n4821, A4 => 
                           n4822, ZN => n4809);
   U7746 : AOI221_X1 port map( B1 => n13992, B2 => n8174, C1 => n13989, C2 => 
                           n8142, A => n4825, ZN => n4820);
   U7747 : AOI221_X1 port map( B1 => n13977, B2 => n2466, C1 => n13974, C2 => 
                           n2445, A => n4826, ZN => n4819);
   U7748 : AOI221_X1 port map( B1 => n14005, B2 => n1951, C1 => n14001, C2 => 
                           n1975, A => n4824, ZN => n4821);
   U7749 : NAND4_X1 port map( A1 => n4856, A2 => n4857, A3 => n4858, A4 => 
                           n4859, ZN => n4846);
   U7750 : AOI221_X1 port map( B1 => n13992, B2 => n8173, C1 => n13989, C2 => 
                           n8141, A => n4862, ZN => n4857);
   U7751 : AOI221_X1 port map( B1 => n13977, B2 => n2465, C1 => n13974, C2 => 
                           n2444, A => n4863, ZN => n4856);
   U7752 : AOI221_X1 port map( B1 => n14005, B2 => n1950, C1 => n14001, C2 => 
                           n1974, A => n4861, ZN => n4858);
   U7753 : NAND4_X1 port map( A1 => n4893, A2 => n4894, A3 => n4895, A4 => 
                           n4896, ZN => n4883);
   U7754 : AOI221_X1 port map( B1 => n13992, B2 => n8172, C1 => n13989, C2 => 
                           n8140, A => n4899, ZN => n4894);
   U7755 : AOI221_X1 port map( B1 => n13977, B2 => n2464, C1 => n13974, C2 => 
                           n2443, A => n4900, ZN => n4893);
   U7756 : AOI221_X1 port map( B1 => n14005, B2 => n1949, C1 => n14001, C2 => 
                           n1973, A => n4898, ZN => n4895);
   U7757 : NAND4_X1 port map( A1 => n4930, A2 => n4931, A3 => n4932, A4 => 
                           n4933, ZN => n4920);
   U7758 : AOI221_X1 port map( B1 => n13992, B2 => n8171, C1 => n13989, C2 => 
                           n8139, A => n4936, ZN => n4931);
   U7759 : AOI221_X1 port map( B1 => n13977, B2 => n2463, C1 => n13974, C2 => 
                           n2442, A => n4937, ZN => n4930);
   U7760 : AOI221_X1 port map( B1 => n14005, B2 => n1948, C1 => n14001, C2 => 
                           n1972, A => n4935, ZN => n4932);
   U7761 : NAND4_X1 port map( A1 => n6103, A2 => n6104, A3 => n6105, A4 => 
                           n6106, ZN => n6093);
   U7762 : AOI221_X1 port map( B1 => n13757, B2 => n2467, C1 => n13754, C2 => 
                           n2446, A => n6110, ZN => n6103);
   U7763 : AOI221_X1 port map( B1 => n13784, B2 => n1976, C1 => n13781, C2 => 
                           n1952, A => n6108, ZN => n6105);
   U7764 : AOI221_X1 port map( B1 => n13772, B2 => n8175, C1 => n13769, C2 => 
                           n8143, A => n6109, ZN => n6104);
   U7765 : NAND4_X1 port map( A1 => n6140, A2 => n6141, A3 => n6142, A4 => 
                           n6143, ZN => n6130);
   U7766 : AOI221_X1 port map( B1 => n13772, B2 => n8174, C1 => n13769, C2 => 
                           n8142, A => n6146, ZN => n6141);
   U7767 : AOI221_X1 port map( B1 => n13757, B2 => n2466, C1 => n13754, C2 => 
                           n2445, A => n6147, ZN => n6140);
   U7768 : AOI221_X1 port map( B1 => n13784, B2 => n1975, C1 => n13781, C2 => 
                           n1951, A => n6145, ZN => n6142);
   U7769 : NAND4_X1 port map( A1 => n6177, A2 => n6178, A3 => n6179, A4 => 
                           n6180, ZN => n6167);
   U7770 : AOI221_X1 port map( B1 => n13772, B2 => n8173, C1 => n13769, C2 => 
                           n8141, A => n6183, ZN => n6178);
   U7771 : AOI221_X1 port map( B1 => n13757, B2 => n2465, C1 => n13754, C2 => 
                           n2444, A => n6184, ZN => n6177);
   U7772 : AOI221_X1 port map( B1 => n13784, B2 => n1974, C1 => n13781, C2 => 
                           n1950, A => n6182, ZN => n6179);
   U7773 : NAND4_X1 port map( A1 => n6214, A2 => n6215, A3 => n6216, A4 => 
                           n6217, ZN => n6204);
   U7774 : AOI221_X1 port map( B1 => n13772, B2 => n8172, C1 => n13769, C2 => 
                           n8140, A => n6220, ZN => n6215);
   U7775 : AOI221_X1 port map( B1 => n13757, B2 => n2464, C1 => n13754, C2 => 
                           n2443, A => n6221, ZN => n6214);
   U7776 : AOI221_X1 port map( B1 => n13784, B2 => n1973, C1 => n13781, C2 => 
                           n1949, A => n6219, ZN => n6216);
   U7777 : NAND4_X1 port map( A1 => n6251, A2 => n6252, A3 => n6253, A4 => 
                           n6254, ZN => n6241);
   U7778 : AOI221_X1 port map( B1 => n13772, B2 => n8171, C1 => n13769, C2 => 
                           n8139, A => n6257, ZN => n6252);
   U7779 : AOI221_X1 port map( B1 => n13757, B2 => n2463, C1 => n13754, C2 => 
                           n2442, A => n6258, ZN => n6251);
   U7780 : AOI221_X1 port map( B1 => n13784, B2 => n1972, C1 => n13781, C2 => 
                           n1948, A => n6256, ZN => n6253);
   U7781 : NAND4_X1 port map( A1 => n6288, A2 => n6289, A3 => n6290, A4 => 
                           n6291, ZN => n6278);
   U7782 : AOI221_X1 port map( B1 => n13772, B2 => n8170, C1 => n13769, C2 => 
                           n8138, A => n6294, ZN => n6289);
   U7783 : AOI221_X1 port map( B1 => n13757, B2 => n2462, C1 => n13754, C2 => 
                           n2441, A => n6295, ZN => n6288);
   U7784 : AOI221_X1 port map( B1 => n13784, B2 => n1971, C1 => n13781, C2 => 
                           n1947, A => n6293, ZN => n6290);
   U7785 : NAND4_X1 port map( A1 => n6325, A2 => n6326, A3 => n6327, A4 => 
                           n6328, ZN => n6315);
   U7786 : AOI221_X1 port map( B1 => n13772, B2 => n8169, C1 => n13769, C2 => 
                           n8137, A => n6331, ZN => n6326);
   U7787 : AOI221_X1 port map( B1 => n13757, B2 => n2461, C1 => n13754, C2 => 
                           n2440, A => n6332, ZN => n6325);
   U7788 : AOI221_X1 port map( B1 => n13784, B2 => n1970, C1 => n13781, C2 => 
                           n1946, A => n6330, ZN => n6327);
   U7789 : NAND4_X1 port map( A1 => n6362, A2 => n6363, A3 => n6364, A4 => 
                           n6365, ZN => n6352);
   U7790 : AOI221_X1 port map( B1 => n13772, B2 => n8168, C1 => n13769, C2 => 
                           n8136, A => n6368, ZN => n6363);
   U7791 : AOI221_X1 port map( B1 => n13757, B2 => n2460, C1 => n13754, C2 => 
                           n2439, A => n6369, ZN => n6362);
   U7792 : AOI221_X1 port map( B1 => n13784, B2 => n1969, C1 => n13781, C2 => 
                           n1945, A => n6367, ZN => n6364);
   U7793 : NAND4_X1 port map( A1 => n6399, A2 => n6400, A3 => n6401, A4 => 
                           n6402, ZN => n6389);
   U7794 : AOI221_X1 port map( B1 => n13772, B2 => n8167, C1 => n13769, C2 => 
                           n8135, A => n6405, ZN => n6400);
   U7795 : AOI221_X1 port map( B1 => n13757, B2 => n2486, C1 => n13754, C2 => 
                           n2485, A => n6406, ZN => n6399);
   U7796 : AOI221_X1 port map( B1 => n13784, B2 => n1968, C1 => n13781, C2 => 
                           n1944, A => n6404, ZN => n6401);
   U7797 : NAND4_X1 port map( A1 => n6436, A2 => n6437, A3 => n6438, A4 => 
                           n6439, ZN => n6426);
   U7798 : AOI221_X1 port map( B1 => n13772, B2 => n8166, C1 => n13769, C2 => 
                           n8134, A => n6442, ZN => n6437);
   U7799 : AOI221_X1 port map( B1 => n13757, B2 => n2410, C1 => n13754, C2 => 
                           n2408, A => n6443, ZN => n6436);
   U7800 : AOI221_X1 port map( B1 => n13784, B2 => n1967, C1 => n13781, C2 => 
                           n1943, A => n6441, ZN => n6438);
   U7801 : NAND4_X1 port map( A1 => n6473, A2 => n6474, A3 => n6475, A4 => 
                           n6476, ZN => n6463);
   U7802 : AOI221_X1 port map( B1 => n13772, B2 => n8165, C1 => n13769, C2 => 
                           n8133, A => n6479, ZN => n6474);
   U7803 : AOI221_X1 port map( B1 => n13757, B2 => n2409, C1 => n13754, C2 => 
                           n2407, A => n6480, ZN => n6473);
   U7804 : AOI221_X1 port map( B1 => n13784, B2 => n1966, C1 => n13781, C2 => 
                           n1942, A => n6478, ZN => n6475);
   U7805 : NAND4_X1 port map( A1 => n4708, A2 => n4709, A3 => n4710, A4 => 
                           n4711, ZN => n4698);
   U7806 : AOI221_X1 port map( B1 => n13993, B2 => n8177, C1 => n13990, C2 => 
                           n8145, A => n4714, ZN => n4709);
   U7807 : AOI221_X1 port map( B1 => n13978, B2 => n2469, C1 => n13975, C2 => 
                           n2448, A => n4715, ZN => n4708);
   U7808 : AOI221_X1 port map( B1 => n14005, B2 => n1954, C1 => n14002, C2 => 
                           n1978, A => n4713, ZN => n4710);
   U7809 : NAND4_X1 port map( A1 => n4745, A2 => n4746, A3 => n4747, A4 => 
                           n4748, ZN => n4735);
   U7810 : AOI221_X1 port map( B1 => n14005, B2 => n1953, C1 => n14002, C2 => 
                           n1977, A => n4750, ZN => n4747);
   U7811 : AOI221_X1 port map( B1 => n13978, B2 => n821, C1 => n13975, C2 => 
                           n822, A => n4752, ZN => n4745);
   U7812 : AOI221_X1 port map( B1 => n13993, B2 => n1617, C1 => n13990, C2 => 
                           n1638, A => n4751, ZN => n4746);
   U7813 : NAND4_X1 port map( A1 => n6029, A2 => n6030, A3 => n6031, A4 => 
                           n6032, ZN => n6019);
   U7814 : AOI221_X1 port map( B1 => n13773, B2 => n8177, C1 => n13770, C2 => 
                           n8145, A => n6035, ZN => n6030);
   U7815 : AOI221_X1 port map( B1 => n13758, B2 => n2469, C1 => n13755, C2 => 
                           n2448, A => n6036, ZN => n6029);
   U7816 : AOI221_X1 port map( B1 => n13785, B2 => n1978, C1 => n13782, C2 => 
                           n1954, A => n6034, ZN => n6031);
   U7817 : NAND4_X1 port map( A1 => n6066, A2 => n6067, A3 => n6068, A4 => 
                           n6069, ZN => n6056);
   U7818 : AOI221_X1 port map( B1 => n13785, B2 => n1977, C1 => n13782, C2 => 
                           n1953, A => n6071, ZN => n6068);
   U7819 : AOI221_X1 port map( B1 => n13758, B2 => n821, C1 => n13755, C2 => 
                           n822, A => n6073, ZN => n6066);
   U7820 : AOI221_X1 port map( B1 => n13773, B2 => n1617, C1 => n13770, C2 => 
                           n1638, A => n6072, ZN => n6067);
   U7821 : NAND4_X1 port map( A1 => n6521, A2 => n6522, A3 => n6523, A4 => 
                           n6524, ZN => n6500);
   U7822 : AOI221_X1 port map( B1 => n13772, B2 => n8164, C1 => n13769, C2 => 
                           n8132, A => n6529, ZN => n6522);
   U7823 : AOI221_X1 port map( B1 => n13757, B2 => n2459, C1 => n13754, C2 => 
                           n2438, A => n6530, ZN => n6521);
   U7824 : AOI221_X1 port map( B1 => n13784, B2 => n1965, C1 => n13781, C2 => 
                           n897, A => n6528, ZN => n6523);
   U7825 : NAND4_X1 port map( A1 => n4967, A2 => n4968, A3 => n4969, A4 => 
                           n4970, ZN => n4957);
   U7826 : AOI221_X1 port map( B1 => n13992, B2 => n8170, C1 => n13989, C2 => 
                           n8138, A => n4973, ZN => n4968);
   U7827 : AOI221_X1 port map( B1 => n13977, B2 => n2462, C1 => n13974, C2 => 
                           n2441, A => n4974, ZN => n4967);
   U7828 : AOI221_X1 port map( B1 => n14006, B2 => n1947, C1 => n14001, C2 => 
                           n1971, A => n4972, ZN => n4969);
   U7829 : NAND4_X1 port map( A1 => n5004, A2 => n5005, A3 => n5006, A4 => 
                           n5007, ZN => n4994);
   U7830 : AOI221_X1 port map( B1 => n13992, B2 => n8169, C1 => n13989, C2 => 
                           n8137, A => n5010, ZN => n5005);
   U7831 : AOI221_X1 port map( B1 => n13977, B2 => n2461, C1 => n13974, C2 => 
                           n2440, A => n5011, ZN => n5004);
   U7832 : AOI221_X1 port map( B1 => n14006, B2 => n1946, C1 => n14001, C2 => 
                           n1970, A => n5009, ZN => n5006);
   U7833 : NAND4_X1 port map( A1 => n5041, A2 => n5042, A3 => n5043, A4 => 
                           n5044, ZN => n5031);
   U7834 : AOI221_X1 port map( B1 => n13992, B2 => n8168, C1 => n13989, C2 => 
                           n8136, A => n5047, ZN => n5042);
   U7835 : AOI221_X1 port map( B1 => n13977, B2 => n2460, C1 => n13974, C2 => 
                           n2439, A => n5048, ZN => n5041);
   U7836 : AOI221_X1 port map( B1 => n14006, B2 => n1945, C1 => n14001, C2 => 
                           n1969, A => n5046, ZN => n5043);
   U7837 : NAND4_X1 port map( A1 => n5078, A2 => n5079, A3 => n5080, A4 => 
                           n5081, ZN => n5068);
   U7838 : AOI221_X1 port map( B1 => n13992, B2 => n8167, C1 => n13989, C2 => 
                           n8135, A => n5084, ZN => n5079);
   U7839 : AOI221_X1 port map( B1 => n13977, B2 => n2486, C1 => n13974, C2 => 
                           n2485, A => n5085, ZN => n5078);
   U7840 : AOI221_X1 port map( B1 => n14006, B2 => n1944, C1 => n14001, C2 => 
                           n1968, A => n5083, ZN => n5080);
   U7841 : NAND4_X1 port map( A1 => n5115, A2 => n5116, A3 => n5117, A4 => 
                           n5118, ZN => n5105);
   U7842 : AOI221_X1 port map( B1 => n13992, B2 => n8166, C1 => n13989, C2 => 
                           n8134, A => n5121, ZN => n5116);
   U7843 : AOI221_X1 port map( B1 => n13977, B2 => n2410, C1 => n13974, C2 => 
                           n2408, A => n5122, ZN => n5115);
   U7844 : AOI221_X1 port map( B1 => n14006, B2 => n1943, C1 => n14001, C2 => 
                           n1967, A => n5120, ZN => n5117);
   U7845 : NAND4_X1 port map( A1 => n5152, A2 => n5153, A3 => n5154, A4 => 
                           n5155, ZN => n5142);
   U7846 : AOI221_X1 port map( B1 => n13992, B2 => n8165, C1 => n13989, C2 => 
                           n8133, A => n5158, ZN => n5153);
   U7847 : AOI221_X1 port map( B1 => n13977, B2 => n2409, C1 => n13974, C2 => 
                           n2407, A => n5159, ZN => n5152);
   U7848 : AOI221_X1 port map( B1 => n14006, B2 => n1942, C1 => n14001, C2 => 
                           n1966, A => n5157, ZN => n5154);
   U7849 : NAND4_X1 port map( A1 => n3988, A2 => n3989, A3 => n3990, A4 => 
                           n3991, ZN => n3960);
   U7850 : AOI221_X1 port map( B1 => n13994, B2 => n8195, C1 => n13991, C2 => 
                           n8163, A => n4005, ZN => n3989);
   U7851 : AOI221_X1 port map( B1 => n13979, B2 => n1846, C1 => n13976, C2 => 
                           n1838, A => n4011, ZN => n3988);
   U7852 : AOI221_X1 port map( B1 => n896, B2 => n14006, C1 => n14003, C2 => 
                           n1806, A => n4000, ZN => n3990);
   U7853 : NAND4_X1 port map( A1 => n5309, A2 => n5310, A3 => n5311, A4 => 
                           n5312, ZN => n5281);
   U7854 : AOI221_X1 port map( B1 => n13774, B2 => n8195, C1 => n13771, C2 => 
                           n8163, A => n5326, ZN => n5310);
   U7855 : AOI221_X1 port map( B1 => n13759, B2 => n1846, C1 => n13756, C2 => 
                           n1838, A => n5332, ZN => n5309);
   U7856 : AOI221_X1 port map( B1 => n13786, B2 => n1806, C1 => n13783, C2 => 
                           n896, A => n5321, ZN => n5311);
   U7857 : NAND4_X1 port map( A1 => n6577, A2 => n6578, A3 => n6579, A4 => 
                           n6580, ZN => n6562);
   U7858 : AOI221_X1 port map( B1 => n8639, B2 => n14174, C1 => n8607, C2 => 
                           n14171, A => n6585, ZN => n6577);
   U7859 : AOI221_X1 port map( B1 => n8449, B2 => n14201, C1 => n8417, C2 => 
                           n14198, A => n6583, ZN => n6579);
   U7860 : AOI221_X1 port map( B1 => n14189, B2 => n1750, C1 => n8481, C2 => 
                           n14186, A => n6584, ZN => n6578);
   U7861 : NAND4_X1 port map( A1 => n4077, A2 => n4078, A3 => n4079, A4 => 
                           n4080, ZN => n4067);
   U7862 : AOI221_X1 port map( B1 => n13994, B2 => n8194, C1 => n13991, C2 => 
                           n8162, A => n4083, ZN => n4078);
   U7863 : AOI221_X1 port map( B1 => n13979, B2 => n1845, C1 => n13976, C2 => 
                           n1837, A => n4084, ZN => n4077);
   U7864 : AOI221_X1 port map( B1 => n14004, B2 => n1798, C1 => n14003, C2 => 
                           n1805, A => n4082, ZN => n4079);
   U7865 : NAND4_X1 port map( A1 => n4116, A2 => n4117, A3 => n4118, A4 => 
                           n4119, ZN => n4106);
   U7866 : AOI221_X1 port map( B1 => n13994, B2 => n8193, C1 => n13991, C2 => 
                           n8161, A => n4122, ZN => n4117);
   U7867 : AOI221_X1 port map( B1 => n13979, B2 => n1844, C1 => n13976, C2 => 
                           n1836, A => n4123, ZN => n4116);
   U7868 : AOI221_X1 port map( B1 => n14004, B2 => n1797, C1 => n14003, C2 => 
                           n1804, A => n4121, ZN => n4118);
   U7869 : NAND4_X1 port map( A1 => n5437, A2 => n5438, A3 => n5439, A4 => 
                           n5440, ZN => n5427);
   U7870 : AOI221_X1 port map( B1 => n13774, B2 => n8193, C1 => n13771, C2 => 
                           n8161, A => n5443, ZN => n5438);
   U7871 : AOI221_X1 port map( B1 => n13759, B2 => n1844, C1 => n13756, C2 => 
                           n1836, A => n5444, ZN => n5437);
   U7872 : AOI221_X1 port map( B1 => n13786, B2 => n1804, C1 => n13783, C2 => 
                           n1797, A => n5442, ZN => n5439);
   U7873 : NAND4_X1 port map( A1 => n4153, A2 => n4154, A3 => n4155, A4 => 
                           n4156, ZN => n4143);
   U7874 : AOI221_X1 port map( B1 => n13994, B2 => n8192, C1 => n13991, C2 => 
                           n8160, A => n4159, ZN => n4154);
   U7875 : AOI221_X1 port map( B1 => n13979, B2 => n1843, C1 => n13976, C2 => 
                           n1835, A => n4160, ZN => n4153);
   U7876 : AOI221_X1 port map( B1 => n14004, B2 => n1796, C1 => n14003, C2 => 
                           n1803, A => n4158, ZN => n4155);
   U7877 : NAND4_X1 port map( A1 => n4190, A2 => n4191, A3 => n4192, A4 => 
                           n4193, ZN => n4180);
   U7878 : AOI221_X1 port map( B1 => n13994, B2 => n8191, C1 => n13991, C2 => 
                           n8159, A => n4196, ZN => n4191);
   U7879 : AOI221_X1 port map( B1 => n13979, B2 => n1842, C1 => n13976, C2 => 
                           n1834, A => n4197, ZN => n4190);
   U7880 : AOI221_X1 port map( B1 => n14004, B2 => n1795, C1 => n14003, C2 => 
                           n1802, A => n4195, ZN => n4192);
   U7881 : NAND4_X1 port map( A1 => n4227, A2 => n4228, A3 => n4229, A4 => 
                           n4230, ZN => n4217);
   U7882 : AOI221_X1 port map( B1 => n13994, B2 => n8190, C1 => n13991, C2 => 
                           n8158, A => n4233, ZN => n4228);
   U7883 : AOI221_X1 port map( B1 => n13979, B2 => n1841, C1 => n13976, C2 => 
                           n1833, A => n4234, ZN => n4227);
   U7884 : AOI221_X1 port map( B1 => n14004, B2 => n1794, C1 => n14003, C2 => 
                           n1801, A => n4232, ZN => n4229);
   U7885 : NAND4_X1 port map( A1 => n4301, A2 => n4302, A3 => n4303, A4 => 
                           n4304, ZN => n4291);
   U7886 : AOI221_X1 port map( B1 => n13994, B2 => n8188, C1 => n13991, C2 => 
                           n8156, A => n4307, ZN => n4302);
   U7887 : AOI221_X1 port map( B1 => n13979, B2 => n1839, C1 => n13976, C2 => 
                           n1831, A => n4308, ZN => n4301);
   U7888 : AOI221_X1 port map( B1 => n14004, B2 => n1792, C1 => n14003, C2 => 
                           n1799, A => n4306, ZN => n4303);
   U7889 : NAND4_X1 port map( A1 => n5622, A2 => n5623, A3 => n5624, A4 => 
                           n5625, ZN => n5612);
   U7890 : AOI221_X1 port map( B1 => n13774, B2 => n8188, C1 => n13771, C2 => 
                           n8156, A => n5628, ZN => n5623);
   U7891 : AOI221_X1 port map( B1 => n13759, B2 => n1839, C1 => n13756, C2 => 
                           n1831, A => n5629, ZN => n5622);
   U7892 : AOI221_X1 port map( B1 => n13786, B2 => n1799, C1 => n13783, C2 => 
                           n1792, A => n5627, ZN => n5624);
   U7893 : NAND4_X1 port map( A1 => n4338, A2 => n4339, A3 => n4340, A4 => 
                           n4341, ZN => n4328);
   U7894 : AOI221_X1 port map( B1 => n13993, B2 => n8187, C1 => n13990, C2 => 
                           n8155, A => n4344, ZN => n4339);
   U7895 : AOI221_X1 port map( B1 => n13978, B2 => n2479, C1 => n13975, C2 => 
                           n2458, A => n4345, ZN => n4338);
   U7896 : AOI221_X1 port map( B1 => n14005, B2 => n1964, C1 => n14002, C2 => 
                           n1988, A => n4343, ZN => n4340);
   U7897 : NAND4_X1 port map( A1 => n5659, A2 => n5660, A3 => n5661, A4 => 
                           n5662, ZN => n5649);
   U7898 : AOI221_X1 port map( B1 => n13773, B2 => n8187, C1 => n13770, C2 => 
                           n8155, A => n5665, ZN => n5660);
   U7899 : AOI221_X1 port map( B1 => n13758, B2 => n2479, C1 => n13755, C2 => 
                           n2458, A => n5666, ZN => n5659);
   U7900 : AOI221_X1 port map( B1 => n13785, B2 => n1988, C1 => n13782, C2 => 
                           n1964, A => n5664, ZN => n5661);
   U7901 : NAND4_X1 port map( A1 => n4375, A2 => n4376, A3 => n4377, A4 => 
                           n4378, ZN => n4365);
   U7902 : AOI221_X1 port map( B1 => n13993, B2 => n8186, C1 => n13990, C2 => 
                           n8154, A => n4381, ZN => n4376);
   U7903 : AOI221_X1 port map( B1 => n13978, B2 => n2478, C1 => n13975, C2 => 
                           n2457, A => n4382, ZN => n4375);
   U7904 : AOI221_X1 port map( B1 => n14004, B2 => n1963, C1 => n14002, C2 => 
                           n1987, A => n4380, ZN => n4377);
   U7905 : NAND4_X1 port map( A1 => n5696, A2 => n5697, A3 => n5698, A4 => 
                           n5699, ZN => n5686);
   U7906 : AOI221_X1 port map( B1 => n13773, B2 => n8186, C1 => n13770, C2 => 
                           n8154, A => n5702, ZN => n5697);
   U7907 : AOI221_X1 port map( B1 => n13758, B2 => n2478, C1 => n13755, C2 => 
                           n2457, A => n5703, ZN => n5696);
   U7908 : AOI221_X1 port map( B1 => n13785, B2 => n1987, C1 => n13782, C2 => 
                           n1963, A => n5701, ZN => n5698);
   U7909 : NAND4_X1 port map( A1 => n3150, A2 => n3151, A3 => n3152, A4 => 
                           n3153, ZN => n3140);
   U7910 : AOI221_X1 port map( B1 => n8630, B2 => n14175, C1 => n8598, C2 => 
                           n14172, A => n3157, ZN => n3150);
   U7911 : AOI221_X1 port map( B1 => n8440, B2 => n14202, C1 => n8408, C2 => 
                           n14199, A => n3155, ZN => n3152);
   U7912 : AOI221_X1 port map( B1 => n14189, B2 => n2117, C1 => n8472, C2 => 
                           n14187, A => n3156, ZN => n3151);
   U7913 : NAND4_X1 port map( A1 => n4412, A2 => n4413, A3 => n4414, A4 => 
                           n4415, ZN => n4402);
   U7914 : AOI221_X1 port map( B1 => n13993, B2 => n8185, C1 => n13990, C2 => 
                           n8153, A => n4418, ZN => n4413);
   U7915 : AOI221_X1 port map( B1 => n13978, B2 => n2477, C1 => n13975, C2 => 
                           n2456, A => n4419, ZN => n4412);
   U7916 : AOI221_X1 port map( B1 => n14004, B2 => n1962, C1 => n14002, C2 => 
                           n1986, A => n4417, ZN => n4414);
   U7917 : NAND4_X1 port map( A1 => n5733, A2 => n5734, A3 => n5735, A4 => 
                           n5736, ZN => n5723);
   U7918 : AOI221_X1 port map( B1 => n13773, B2 => n8185, C1 => n13770, C2 => 
                           n8153, A => n5739, ZN => n5734);
   U7919 : AOI221_X1 port map( B1 => n13758, B2 => n2477, C1 => n13755, C2 => 
                           n2456, A => n5740, ZN => n5733);
   U7920 : AOI221_X1 port map( B1 => n13785, B2 => n1986, C1 => n13782, C2 => 
                           n1962, A => n5738, ZN => n5735);
   U7921 : NAND4_X1 port map( A1 => n3187, A2 => n3188, A3 => n3189, A4 => 
                           n3190, ZN => n3177);
   U7922 : AOI221_X1 port map( B1 => n8629, B2 => n14175, C1 => n8597, C2 => 
                           n14172, A => n3194, ZN => n3187);
   U7923 : AOI221_X1 port map( B1 => n8439, B2 => n14202, C1 => n8407, C2 => 
                           n14199, A => n3192, ZN => n3189);
   U7924 : AOI221_X1 port map( B1 => n14189, B2 => n2116, C1 => n8471, C2 => 
                           n14187, A => n3193, ZN => n3188);
   U7925 : NAND4_X1 port map( A1 => n4449, A2 => n4450, A3 => n4451, A4 => 
                           n4452, ZN => n4439);
   U7926 : AOI221_X1 port map( B1 => n13993, B2 => n8184, C1 => n13990, C2 => 
                           n8152, A => n4455, ZN => n4450);
   U7927 : AOI221_X1 port map( B1 => n13978, B2 => n2476, C1 => n13975, C2 => 
                           n2455, A => n4456, ZN => n4449);
   U7928 : AOI221_X1 port map( B1 => n14004, B2 => n1961, C1 => n14002, C2 => 
                           n1985, A => n4454, ZN => n4451);
   U7929 : NAND4_X1 port map( A1 => n5770, A2 => n5771, A3 => n5772, A4 => 
                           n5773, ZN => n5760);
   U7930 : AOI221_X1 port map( B1 => n13773, B2 => n8184, C1 => n13770, C2 => 
                           n8152, A => n5776, ZN => n5771);
   U7931 : AOI221_X1 port map( B1 => n13758, B2 => n2476, C1 => n13755, C2 => 
                           n2455, A => n5777, ZN => n5770);
   U7932 : AOI221_X1 port map( B1 => n13785, B2 => n1985, C1 => n13782, C2 => 
                           n1961, A => n5775, ZN => n5772);
   U7933 : NAND4_X1 port map( A1 => n3224, A2 => n3225, A3 => n3226, A4 => 
                           n3227, ZN => n3214);
   U7934 : AOI221_X1 port map( B1 => n8628, B2 => n14175, C1 => n8596, C2 => 
                           n14172, A => n3231, ZN => n3224);
   U7935 : AOI221_X1 port map( B1 => n8438, B2 => n14202, C1 => n8406, C2 => 
                           n14199, A => n3229, ZN => n3226);
   U7936 : AOI221_X1 port map( B1 => n14189, B2 => n2115, C1 => n8470, C2 => 
                           n14187, A => n3230, ZN => n3225);
   U7937 : NAND4_X1 port map( A1 => n4486, A2 => n4487, A3 => n4488, A4 => 
                           n4489, ZN => n4476);
   U7938 : AOI221_X1 port map( B1 => n13993, B2 => n8183, C1 => n13990, C2 => 
                           n8151, A => n4492, ZN => n4487);
   U7939 : AOI221_X1 port map( B1 => n13978, B2 => n2475, C1 => n13975, C2 => 
                           n2454, A => n4493, ZN => n4486);
   U7940 : AOI221_X1 port map( B1 => n14004, B2 => n1960, C1 => n14002, C2 => 
                           n1984, A => n4491, ZN => n4488);
   U7941 : NAND4_X1 port map( A1 => n5807, A2 => n5808, A3 => n5809, A4 => 
                           n5810, ZN => n5797);
   U7942 : AOI221_X1 port map( B1 => n13773, B2 => n8183, C1 => n13770, C2 => 
                           n8151, A => n5813, ZN => n5808);
   U7943 : AOI221_X1 port map( B1 => n13758, B2 => n2475, C1 => n13755, C2 => 
                           n2454, A => n5814, ZN => n5807);
   U7944 : AOI221_X1 port map( B1 => n13785, B2 => n1984, C1 => n13782, C2 => 
                           n1960, A => n5812, ZN => n5809);
   U7945 : NAND4_X1 port map( A1 => n3261, A2 => n3262, A3 => n3263, A4 => 
                           n3264, ZN => n3251);
   U7946 : AOI221_X1 port map( B1 => n8627, B2 => n14175, C1 => n8595, C2 => 
                           n14172, A => n3268, ZN => n3261);
   U7947 : AOI221_X1 port map( B1 => n8437, B2 => n14202, C1 => n8405, C2 => 
                           n14199, A => n3266, ZN => n3263);
   U7948 : AOI221_X1 port map( B1 => n14189, B2 => n2114, C1 => n8469, C2 => 
                           n14187, A => n3267, ZN => n3262);
   U7949 : NAND4_X1 port map( A1 => n4523, A2 => n4524, A3 => n4525, A4 => 
                           n4526, ZN => n4513);
   U7950 : AOI221_X1 port map( B1 => n13978, B2 => n2474, C1 => n13975, C2 => 
                           n2453, A => n4530, ZN => n4523);
   U7951 : AOI221_X1 port map( B1 => n14004, B2 => n1959, C1 => n14002, C2 => 
                           n1983, A => n4528, ZN => n4525);
   U7952 : AOI221_X1 port map( B1 => n13993, B2 => n8182, C1 => n13990, C2 => 
                           n8150, A => n4529, ZN => n4524);
   U7953 : NAND4_X1 port map( A1 => n5844, A2 => n5845, A3 => n5846, A4 => 
                           n5847, ZN => n5834);
   U7954 : AOI221_X1 port map( B1 => n13758, B2 => n2474, C1 => n13755, C2 => 
                           n2453, A => n5851, ZN => n5844);
   U7955 : AOI221_X1 port map( B1 => n13785, B2 => n1983, C1 => n13782, C2 => 
                           n1959, A => n5849, ZN => n5846);
   U7956 : AOI221_X1 port map( B1 => n13773, B2 => n8182, C1 => n13770, C2 => 
                           n8150, A => n5850, ZN => n5845);
   U7957 : NAND4_X1 port map( A1 => n3298, A2 => n3299, A3 => n3300, A4 => 
                           n3301, ZN => n3288);
   U7958 : AOI221_X1 port map( B1 => n8626, B2 => n14175, C1 => n8594, C2 => 
                           n14172, A => n3305, ZN => n3298);
   U7959 : AOI221_X1 port map( B1 => n8436, B2 => n14202, C1 => n8404, C2 => 
                           n14199, A => n3303, ZN => n3300);
   U7960 : AOI221_X1 port map( B1 => n14190, B2 => n2113, C1 => n8468, C2 => 
                           n14187, A => n3304, ZN => n3299);
   U7961 : NAND4_X1 port map( A1 => n4560, A2 => n4561, A3 => n4562, A4 => 
                           n4563, ZN => n4550);
   U7962 : AOI221_X1 port map( B1 => n13978, B2 => n2473, C1 => n13975, C2 => 
                           n2452, A => n4567, ZN => n4560);
   U7963 : AOI221_X1 port map( B1 => n14005, B2 => n1958, C1 => n14002, C2 => 
                           n1982, A => n4565, ZN => n4562);
   U7964 : AOI221_X1 port map( B1 => n13993, B2 => n8181, C1 => n13990, C2 => 
                           n8149, A => n4566, ZN => n4561);
   U7965 : NAND4_X1 port map( A1 => n5881, A2 => n5882, A3 => n5883, A4 => 
                           n5884, ZN => n5871);
   U7966 : AOI221_X1 port map( B1 => n13758, B2 => n2473, C1 => n13755, C2 => 
                           n2452, A => n5888, ZN => n5881);
   U7967 : AOI221_X1 port map( B1 => n13785, B2 => n1982, C1 => n13782, C2 => 
                           n1958, A => n5886, ZN => n5883);
   U7968 : AOI221_X1 port map( B1 => n13773, B2 => n8181, C1 => n13770, C2 => 
                           n8149, A => n5887, ZN => n5882);
   U7969 : NAND4_X1 port map( A1 => n3337, A2 => n3338, A3 => n3339, A4 => 
                           n3340, ZN => n3327);
   U7970 : AOI221_X1 port map( B1 => n8625, B2 => n14175, C1 => n8593, C2 => 
                           n14172, A => n3344, ZN => n3337);
   U7971 : AOI221_X1 port map( B1 => n8435, B2 => n14202, C1 => n8403, C2 => 
                           n14199, A => n3342, ZN => n3339);
   U7972 : AOI221_X1 port map( B1 => n14190, B2 => n2112, C1 => n8467, C2 => 
                           n14187, A => n3343, ZN => n3338);
   U7973 : NAND4_X1 port map( A1 => n4597, A2 => n4598, A3 => n4599, A4 => 
                           n4600, ZN => n4587);
   U7974 : AOI221_X1 port map( B1 => n13978, B2 => n2472, C1 => n13975, C2 => 
                           n2451, A => n4604, ZN => n4597);
   U7975 : AOI221_X1 port map( B1 => n14005, B2 => n1957, C1 => n14002, C2 => 
                           n1981, A => n4602, ZN => n4599);
   U7976 : AOI221_X1 port map( B1 => n13993, B2 => n8180, C1 => n13990, C2 => 
                           n8148, A => n4603, ZN => n4598);
   U7977 : NAND4_X1 port map( A1 => n5918, A2 => n5919, A3 => n5920, A4 => 
                           n5921, ZN => n5908);
   U7978 : AOI221_X1 port map( B1 => n13758, B2 => n2472, C1 => n13755, C2 => 
                           n2451, A => n5925, ZN => n5918);
   U7979 : AOI221_X1 port map( B1 => n13785, B2 => n1981, C1 => n13782, C2 => 
                           n1957, A => n5923, ZN => n5920);
   U7980 : AOI221_X1 port map( B1 => n13773, B2 => n8180, C1 => n13770, C2 => 
                           n8148, A => n5924, ZN => n5919);
   U7981 : NAND4_X1 port map( A1 => n3374, A2 => n3375, A3 => n3376, A4 => 
                           n3377, ZN => n3364);
   U7982 : AOI221_X1 port map( B1 => n8624, B2 => n14175, C1 => n8592, C2 => 
                           n14172, A => n3381, ZN => n3374);
   U7983 : AOI221_X1 port map( B1 => n8434, B2 => n14202, C1 => n8402, C2 => 
                           n14199, A => n3379, ZN => n3376);
   U7984 : AOI221_X1 port map( B1 => n14190, B2 => n2111, C1 => n8466, C2 => 
                           n14187, A => n3380, ZN => n3375);
   U7985 : NAND4_X1 port map( A1 => n4634, A2 => n4635, A3 => n4636, A4 => 
                           n4637, ZN => n4624);
   U7986 : AOI221_X1 port map( B1 => n13978, B2 => n2471, C1 => n13975, C2 => 
                           n2450, A => n4641, ZN => n4634);
   U7987 : AOI221_X1 port map( B1 => n14005, B2 => n1956, C1 => n14002, C2 => 
                           n1980, A => n4639, ZN => n4636);
   U7988 : AOI221_X1 port map( B1 => n13993, B2 => n8179, C1 => n13990, C2 => 
                           n8147, A => n4640, ZN => n4635);
   U7989 : NAND4_X1 port map( A1 => n5955, A2 => n5956, A3 => n5957, A4 => 
                           n5958, ZN => n5945);
   U7990 : AOI221_X1 port map( B1 => n13758, B2 => n2471, C1 => n13755, C2 => 
                           n2450, A => n5962, ZN => n5955);
   U7991 : AOI221_X1 port map( B1 => n13785, B2 => n1980, C1 => n13782, C2 => 
                           n1956, A => n5960, ZN => n5957);
   U7992 : AOI221_X1 port map( B1 => n13773, B2 => n8179, C1 => n13770, C2 => 
                           n8147, A => n5961, ZN => n5956);
   U7993 : NAND4_X1 port map( A1 => n3411, A2 => n3412, A3 => n3413, A4 => 
                           n3414, ZN => n3401);
   U7994 : AOI221_X1 port map( B1 => n8623, B2 => n14175, C1 => n8591, C2 => 
                           n14172, A => n3418, ZN => n3411);
   U7995 : AOI221_X1 port map( B1 => n8433, B2 => n14202, C1 => n8401, C2 => 
                           n14199, A => n3416, ZN => n3413);
   U7996 : AOI221_X1 port map( B1 => n14190, B2 => n2110, C1 => n8465, C2 => 
                           n14187, A => n3417, ZN => n3412);
   U7997 : NAND4_X1 port map( A1 => n4671, A2 => n4672, A3 => n4673, A4 => 
                           n4674, ZN => n4661);
   U7998 : AOI221_X1 port map( B1 => n13993, B2 => n8178, C1 => n13990, C2 => 
                           n8146, A => n4677, ZN => n4672);
   U7999 : AOI221_X1 port map( B1 => n13978, B2 => n2470, C1 => n13975, C2 => 
                           n2449, A => n4678, ZN => n4671);
   U8000 : AOI221_X1 port map( B1 => n14005, B2 => n1955, C1 => n14002, C2 => 
                           n1979, A => n4676, ZN => n4673);
   U8001 : NAND4_X1 port map( A1 => n5992, A2 => n5993, A3 => n5994, A4 => 
                           n5995, ZN => n5982);
   U8002 : AOI221_X1 port map( B1 => n13773, B2 => n8178, C1 => n13770, C2 => 
                           n8146, A => n5998, ZN => n5993);
   U8003 : AOI221_X1 port map( B1 => n13758, B2 => n2470, C1 => n13755, C2 => 
                           n2449, A => n5999, ZN => n5992);
   U8004 : AOI221_X1 port map( B1 => n13785, B2 => n1979, C1 => n13782, C2 => 
                           n1955, A => n5997, ZN => n5994);
   U8005 : NAND4_X1 port map( A1 => n3448, A2 => n3449, A3 => n3450, A4 => 
                           n3451, ZN => n3438);
   U8006 : AOI221_X1 port map( B1 => n8622, B2 => n14175, C1 => n8590, C2 => 
                           n14172, A => n3455, ZN => n3448);
   U8007 : AOI221_X1 port map( B1 => n8432, B2 => n14202, C1 => n8400, C2 => 
                           n14199, A => n3453, ZN => n3450);
   U8008 : AOI221_X1 port map( B1 => n14190, B2 => n2109, C1 => n8464, C2 => 
                           n14187, A => n3454, ZN => n3449);
   U8009 : NAND4_X1 port map( A1 => n3485, A2 => n3486, A3 => n3487, A4 => 
                           n3488, ZN => n3475);
   U8010 : AOI221_X1 port map( B1 => n8621, B2 => n14175, C1 => n8589, C2 => 
                           n14172, A => n3492, ZN => n3485);
   U8011 : AOI221_X1 port map( B1 => n8431, B2 => n14202, C1 => n8399, C2 => 
                           n14199, A => n3490, ZN => n3487);
   U8012 : AOI221_X1 port map( B1 => n14190, B2 => n2108, C1 => n8463, C2 => 
                           n14187, A => n3491, ZN => n3486);
   U8013 : NAND4_X1 port map( A1 => n3522, A2 => n3523, A3 => n3524, A4 => 
                           n3525, ZN => n3512);
   U8014 : AOI221_X1 port map( B1 => n8620, B2 => n14175, C1 => n8588, C2 => 
                           n14172, A => n3529, ZN => n3522);
   U8015 : AOI221_X1 port map( B1 => n8430, B2 => n14202, C1 => n8398, C2 => 
                           n14199, A => n3527, ZN => n3524);
   U8016 : AOI221_X1 port map( B1 => n14190, B2 => n2107, C1 => n8462, C2 => 
                           n14187, A => n3528, ZN => n3523);
   U8017 : NAND4_X1 port map( A1 => n3559, A2 => n3560, A3 => n3561, A4 => 
                           n3562, ZN => n3549);
   U8018 : AOI221_X1 port map( B1 => n8619, B2 => n14175, C1 => n8587, C2 => 
                           n14172, A => n3566, ZN => n3559);
   U8019 : AOI221_X1 port map( B1 => n8429, B2 => n14202, C1 => n8397, C2 => 
                           n14199, A => n3564, ZN => n3561);
   U8020 : AOI221_X1 port map( B1 => n784, B2 => n14191, C1 => n8461, C2 => 
                           n14187, A => n3565, ZN => n3560);
   U8021 : NAND4_X1 port map( A1 => n3596, A2 => n3597, A3 => n3598, A4 => 
                           n3599, ZN => n3586);
   U8022 : AOI221_X1 port map( B1 => n8618, B2 => n14174, C1 => n8586, C2 => 
                           n14171, A => n3603, ZN => n3596);
   U8023 : AOI221_X1 port map( B1 => n8428, B2 => n14201, C1 => n8396, C2 => 
                           n14198, A => n3601, ZN => n3598);
   U8024 : AOI221_X1 port map( B1 => n14190, B2 => n2105, C1 => n8460, C2 => 
                           n14186, A => n3602, ZN => n3597);
   U8025 : NAND4_X1 port map( A1 => n3633, A2 => n3634, A3 => n3635, A4 => 
                           n3636, ZN => n3623);
   U8026 : AOI221_X1 port map( B1 => n8617, B2 => n14174, C1 => n8585, C2 => 
                           n14171, A => n3640, ZN => n3633);
   U8027 : AOI221_X1 port map( B1 => n8427, B2 => n14201, C1 => n8395, C2 => 
                           n14198, A => n3638, ZN => n3635);
   U8028 : AOI221_X1 port map( B1 => n14190, B2 => n2104, C1 => n8459, C2 => 
                           n14186, A => n3639, ZN => n3634);
   U8029 : NAND4_X1 port map( A1 => n3670, A2 => n3671, A3 => n3672, A4 => 
                           n3673, ZN => n3660);
   U8030 : AOI221_X1 port map( B1 => n8616, B2 => n14174, C1 => n8584, C2 => 
                           n14171, A => n3677, ZN => n3670);
   U8031 : AOI221_X1 port map( B1 => n8426, B2 => n14201, C1 => n8394, C2 => 
                           n14198, A => n3675, ZN => n3672);
   U8032 : AOI221_X1 port map( B1 => n14190, B2 => n2103, C1 => n8458, C2 => 
                           n14186, A => n3676, ZN => n3671);
   U8033 : NAND4_X1 port map( A1 => n3707, A2 => n3708, A3 => n3709, A4 => 
                           n3710, ZN => n3697);
   U8034 : AOI221_X1 port map( B1 => n8615, B2 => n14174, C1 => n8583, C2 => 
                           n14171, A => n3714, ZN => n3707);
   U8035 : AOI221_X1 port map( B1 => n8425, B2 => n14201, C1 => n8393, C2 => 
                           n14198, A => n3712, ZN => n3709);
   U8036 : AOI221_X1 port map( B1 => n14190, B2 => n2102, C1 => n8457, C2 => 
                           n14186, A => n3713, ZN => n3708);
   U8037 : NAND4_X1 port map( A1 => n3744, A2 => n3745, A3 => n3746, A4 => 
                           n3747, ZN => n3734);
   U8038 : AOI221_X1 port map( B1 => n8614, B2 => n14174, C1 => n8582, C2 => 
                           n14171, A => n3751, ZN => n3744);
   U8039 : AOI221_X1 port map( B1 => n8424, B2 => n14201, C1 => n8392, C2 => 
                           n14198, A => n3749, ZN => n3746);
   U8040 : AOI221_X1 port map( B1 => n14191, B2 => n2101, C1 => n8456, C2 => 
                           n14186, A => n3750, ZN => n3745);
   U8041 : NAND4_X1 port map( A1 => n3781, A2 => n3782, A3 => n3783, A4 => 
                           n3784, ZN => n3771);
   U8042 : AOI221_X1 port map( B1 => n8613, B2 => n14174, C1 => n8581, C2 => 
                           n14171, A => n3788, ZN => n3781);
   U8043 : AOI221_X1 port map( B1 => n8423, B2 => n14201, C1 => n8391, C2 => 
                           n14198, A => n3786, ZN => n3783);
   U8044 : AOI221_X1 port map( B1 => n14191, B2 => n2100, C1 => n8455, C2 => 
                           n14186, A => n3787, ZN => n3782);
   U8045 : NAND4_X1 port map( A1 => n3818, A2 => n3819, A3 => n3820, A4 => 
                           n3821, ZN => n3808);
   U8046 : AOI221_X1 port map( B1 => n8612, B2 => n14174, C1 => n8580, C2 => 
                           n14171, A => n3825, ZN => n3818);
   U8047 : AOI221_X1 port map( B1 => n8422, B2 => n14201, C1 => n8390, C2 => 
                           n14198, A => n3823, ZN => n3820);
   U8048 : AOI221_X1 port map( B1 => n14191, B2 => n2099, C1 => n8454, C2 => 
                           n14186, A => n3824, ZN => n3819);
   U8049 : NAND4_X1 port map( A1 => n3855, A2 => n3856, A3 => n3857, A4 => 
                           n3858, ZN => n3845);
   U8050 : AOI221_X1 port map( B1 => n8611, B2 => n14174, C1 => n8579, C2 => 
                           n14171, A => n3862, ZN => n3855);
   U8051 : AOI221_X1 port map( B1 => n8421, B2 => n14201, C1 => n8389, C2 => 
                           n14198, A => n3860, ZN => n3857);
   U8052 : AOI221_X1 port map( B1 => n14191, B2 => n2098, C1 => n8453, C2 => 
                           n14186, A => n3861, ZN => n3856);
   U8053 : NAND4_X1 port map( A1 => n3892, A2 => n3893, A3 => n3894, A4 => 
                           n3895, ZN => n3882);
   U8054 : AOI221_X1 port map( B1 => n8610, B2 => n14174, C1 => n8578, C2 => 
                           n14171, A => n3899, ZN => n3892);
   U8055 : AOI221_X1 port map( B1 => n8420, B2 => n14201, C1 => n8388, C2 => 
                           n14198, A => n3897, ZN => n3894);
   U8056 : AOI221_X1 port map( B1 => n14191, B2 => n2097, C1 => n8452, C2 => 
                           n14186, A => n3898, ZN => n3893);
   U8057 : NAND4_X1 port map( A1 => n3929, A2 => n3930, A3 => n3931, A4 => 
                           n3932, ZN => n3919);
   U8058 : AOI221_X1 port map( B1 => n8609, B2 => n14174, C1 => n8577, C2 => 
                           n14171, A => n3936, ZN => n3929);
   U8059 : AOI221_X1 port map( B1 => n8419, B2 => n14201, C1 => n8387, C2 => 
                           n14198, A => n3934, ZN => n3931);
   U8060 : AOI221_X1 port map( B1 => n14191, B2 => n2096, C1 => n8451, C2 => 
                           n14186, A => n3935, ZN => n3930);
   U8061 : NAND4_X1 port map( A1 => n5251, A2 => n5252, A3 => n5253, A4 => 
                           n5254, ZN => n5241);
   U8062 : AOI221_X1 port map( B1 => n8608, B2 => n14174, C1 => n8576, C2 => 
                           n14171, A => n5258, ZN => n5251);
   U8063 : AOI221_X1 port map( B1 => n8418, B2 => n14201, C1 => n8386, C2 => 
                           n14198, A => n5256, ZN => n5253);
   U8064 : AOI221_X1 port map( B1 => n14191, B2 => n2095, C1 => n8450, C2 => 
                           n14186, A => n5257, ZN => n5252);
   U8065 : NAND4_X1 port map( A1 => n2835, A2 => n2836, A3 => n2837, A4 => 
                           n2838, ZN => n2780);
   U8066 : AOI221_X1 port map( B1 => n14722, B2 => n8162, C1 => n14719, C2 => 
                           n8194, A => n2845, ZN => n2837);
   U8067 : AOI221_X1 port map( B1 => n8320, B2 => n14130, C1 => n8288, C2 => 
                           n14127, A => n2856, ZN => n2835);
   U8068 : AOI221_X1 port map( B1 => n14164, B2 => n1813, C1 => n14161, C2 => 
                           n6760, A => n2841, ZN => n2838);
   U8069 : NAND4_X1 port map( A1 => n2899, A2 => n2900, A3 => n2901, A4 => 
                           n2902, ZN => n2880);
   U8070 : AOI221_X1 port map( B1 => n14722, B2 => n8161, C1 => n14719, C2 => 
                           n8193, A => n2904, ZN => n2901);
   U8071 : AOI221_X1 port map( B1 => n8319, B2 => n14130, C1 => n8287, C2 => 
                           n14127, A => n2906, ZN => n2899);
   U8072 : AOI221_X1 port map( B1 => n14164, B2 => n1812, C1 => n14161, C2 => 
                           n6773, A => n2903, ZN => n2902);
   U8073 : NAND4_X1 port map( A1 => n2936, A2 => n2937, A3 => n2938, A4 => 
                           n2939, ZN => n2917);
   U8074 : AOI221_X1 port map( B1 => n14722, B2 => n8160, C1 => n14719, C2 => 
                           n8192, A => n2941, ZN => n2938);
   U8075 : AOI221_X1 port map( B1 => n8318, B2 => n14130, C1 => n8286, C2 => 
                           n14127, A => n2943, ZN => n2936);
   U8076 : AOI221_X1 port map( B1 => n14164, B2 => n1811, C1 => n14161, C2 => 
                           n6781, A => n2940, ZN => n2939);
   U8077 : NAND4_X1 port map( A1 => n2973, A2 => n2974, A3 => n2975, A4 => 
                           n2976, ZN => n2954);
   U8078 : AOI221_X1 port map( B1 => n14722, B2 => n8159, C1 => n14719, C2 => 
                           n8191, A => n2978, ZN => n2975);
   U8079 : AOI221_X1 port map( B1 => n8317, B2 => n14130, C1 => n8285, C2 => 
                           n14127, A => n2980, ZN => n2973);
   U8080 : AOI221_X1 port map( B1 => n14164, B2 => n1810, C1 => n14161, C2 => 
                           n6795, A => n2977, ZN => n2976);
   U8081 : NAND4_X1 port map( A1 => n3010, A2 => n3011, A3 => n3012, A4 => 
                           n3013, ZN => n2991);
   U8082 : AOI221_X1 port map( B1 => n14722, B2 => n8158, C1 => n14719, C2 => 
                           n8190, A => n3015, ZN => n3012);
   U8083 : AOI221_X1 port map( B1 => n8316, B2 => n14130, C1 => n8284, C2 => 
                           n14127, A => n3017, ZN => n3010);
   U8084 : AOI221_X1 port map( B1 => n14164, B2 => n1809, C1 => n14161, C2 => 
                           n6805, A => n3014, ZN => n3013);
   U8085 : NAND4_X1 port map( A1 => n3047, A2 => n3048, A3 => n3049, A4 => 
                           n3050, ZN => n3028);
   U8086 : AOI221_X1 port map( B1 => n14722, B2 => n8157, C1 => n14719, C2 => 
                           n8189, A => n3052, ZN => n3049);
   U8087 : AOI221_X1 port map( B1 => n8315, B2 => n14130, C1 => n8283, C2 => 
                           n14127, A => n3054, ZN => n3047);
   U8088 : AOI221_X1 port map( B1 => n14164, B2 => n1808, C1 => n14161, C2 => 
                           n6820, A => n3051, ZN => n3050);
   U8089 : NAND4_X1 port map( A1 => n3084, A2 => n3085, A3 => n3086, A4 => 
                           n3087, ZN => n3065);
   U8090 : AOI221_X1 port map( B1 => n14722, B2 => n8156, C1 => n14719, C2 => 
                           n8188, A => n3089, ZN => n3086);
   U8091 : AOI221_X1 port map( B1 => n8314, B2 => n14130, C1 => n8282, C2 => 
                           n14127, A => n3091, ZN => n3084);
   U8092 : AOI221_X1 port map( B1 => n14164, B2 => n1807, C1 => n14161, C2 => 
                           n6832, A => n3088, ZN => n3087);
   U8093 : NAND4_X1 port map( A1 => n3121, A2 => n3122, A3 => n3123, A4 => 
                           n3124, ZN => n3102);
   U8094 : AOI221_X1 port map( B1 => n14722, B2 => n8155, C1 => n14719, C2 => 
                           n8187, A => n3126, ZN => n3123);
   U8095 : AOI221_X1 port map( B1 => n8313, B2 => n14130, C1 => n8281, C2 => 
                           n14127, A => n3128, ZN => n3121);
   U8096 : AOI221_X1 port map( B1 => n14164, B2 => n2009, C1 => n14161, C2 => 
                           n6845, A => n3125, ZN => n3124);
   U8097 : NAND4_X1 port map( A1 => n6586, A2 => n6587, A3 => n6588, A4 => 
                           n6589, ZN => n6561);
   U8098 : AOI221_X1 port map( B1 => n14724, B2 => n8163, C1 => n14721, C2 => 
                           n8195, A => n6592, ZN => n6588);
   U8099 : AOI221_X1 port map( B1 => n8321, B2 => n14128, C1 => n8289, C2 => 
                           n14125, A => n6594, ZN => n6586);
   U8100 : AOI221_X1 port map( B1 => n14162, B2 => n1814, C1 => n14159, C2 => 
                           n7107, A => n6590, ZN => n6589);
   U8101 : NAND4_X1 port map( A1 => n3158, A2 => n3159, A3 => n3160, A4 => 
                           n3161, ZN => n3139);
   U8102 : AOI221_X1 port map( B1 => n14722, B2 => n8154, C1 => n14719, C2 => 
                           n8186, A => n3163, ZN => n3160);
   U8103 : AOI221_X1 port map( B1 => n8312, B2 => n14129, C1 => n8280, C2 => 
                           n14126, A => n3165, ZN => n3158);
   U8104 : AOI221_X1 port map( B1 => n14163, B2 => n2008, C1 => n14160, C2 => 
                           n6859, A => n3162, ZN => n3161);
   U8105 : NAND4_X1 port map( A1 => n3195, A2 => n3196, A3 => n3197, A4 => 
                           n3198, ZN => n3176);
   U8106 : AOI221_X1 port map( B1 => n14722, B2 => n8153, C1 => n14719, C2 => 
                           n8185, A => n3200, ZN => n3197);
   U8107 : AOI221_X1 port map( B1 => n8311, B2 => n14129, C1 => n8279, C2 => 
                           n14126, A => n3202, ZN => n3195);
   U8108 : AOI221_X1 port map( B1 => n14163, B2 => n2007, C1 => n14160, C2 => 
                           n6871, A => n3199, ZN => n3198);
   U8109 : NAND4_X1 port map( A1 => n3232, A2 => n3233, A3 => n3234, A4 => 
                           n3235, ZN => n3213);
   U8110 : AOI221_X1 port map( B1 => n14722, B2 => n8152, C1 => n14719, C2 => 
                           n8184, A => n3237, ZN => n3234);
   U8111 : AOI221_X1 port map( B1 => n8310, B2 => n14129, C1 => n8278, C2 => 
                           n14126, A => n3239, ZN => n3232);
   U8112 : AOI221_X1 port map( B1 => n14163, B2 => n2006, C1 => n14160, C2 => 
                           n6889, A => n3236, ZN => n3235);
   U8113 : NAND4_X1 port map( A1 => n3269, A2 => n3270, A3 => n3271, A4 => 
                           n3272, ZN => n3250);
   U8114 : AOI221_X1 port map( B1 => n14722, B2 => n8151, C1 => n14719, C2 => 
                           n8183, A => n3274, ZN => n3271);
   U8115 : AOI221_X1 port map( B1 => n8309, B2 => n14129, C1 => n8277, C2 => 
                           n14126, A => n3276, ZN => n3269);
   U8116 : AOI221_X1 port map( B1 => n14163, B2 => n2005, C1 => n14160, C2 => 
                           n6898, A => n3273, ZN => n3272);
   U8117 : NAND4_X1 port map( A1 => n3306, A2 => n3307, A3 => n3308, A4 => 
                           n3309, ZN => n3287);
   U8118 : AOI221_X1 port map( B1 => n8308, B2 => n14129, C1 => n8276, C2 => 
                           n14126, A => n3315, ZN => n3306);
   U8119 : AOI221_X1 port map( B1 => n76, B2 => n14147, C1 => n14149, C2 => 
                           n2436, A => n3311, ZN => n3308);
   U8120 : AOI221_X1 port map( B1 => n14163, B2 => n2004, C1 => n14160, C2 => 
                           n6915, A => n3310, ZN => n3309);
   U8121 : NAND4_X1 port map( A1 => n3345, A2 => n3346, A3 => n3347, A4 => 
                           n3348, ZN => n3326);
   U8122 : AOI221_X1 port map( B1 => n8307, B2 => n14129, C1 => n8275, C2 => 
                           n14126, A => n3352, ZN => n3345);
   U8123 : AOI221_X1 port map( B1 => n82, B2 => n14147, C1 => n14149, C2 => 
                           n2435, A => n3350, ZN => n3347);
   U8124 : AOI221_X1 port map( B1 => n14163, B2 => n2003, C1 => n14160, C2 => 
                           n6925, A => n3349, ZN => n3348);
   U8125 : NAND4_X1 port map( A1 => n3382, A2 => n3383, A3 => n3384, A4 => 
                           n3385, ZN => n3363);
   U8126 : AOI221_X1 port map( B1 => n8306, B2 => n14129, C1 => n8274, C2 => 
                           n14126, A => n3389, ZN => n3382);
   U8127 : AOI221_X1 port map( B1 => n88, B2 => n14147, C1 => n14149, C2 => 
                           n2434, A => n3387, ZN => n3384);
   U8128 : AOI221_X1 port map( B1 => n14163, B2 => n2002, C1 => n14160, C2 => 
                           n6940, A => n3386, ZN => n3385);
   U8129 : NAND4_X1 port map( A1 => n3419, A2 => n3420, A3 => n3421, A4 => 
                           n3422, ZN => n3400);
   U8130 : AOI221_X1 port map( B1 => n8305, B2 => n14129, C1 => n8273, C2 => 
                           n14126, A => n3426, ZN => n3419);
   U8131 : AOI221_X1 port map( B1 => n94, B2 => n14147, C1 => n14149, C2 => 
                           n2433, A => n3424, ZN => n3421);
   U8132 : AOI221_X1 port map( B1 => n14163, B2 => n2001, C1 => n14160, C2 => 
                           n6952, A => n3423, ZN => n3422);
   U8133 : NAND4_X1 port map( A1 => n3456, A2 => n3457, A3 => n3458, A4 => 
                           n3459, ZN => n3437);
   U8134 : AOI221_X1 port map( B1 => n14723, B2 => n8146, C1 => n14720, C2 => 
                           n8178, A => n3461, ZN => n3458);
   U8135 : AOI221_X1 port map( B1 => n8304, B2 => n14129, C1 => n8272, C2 => 
                           n14126, A => n3463, ZN => n3456);
   U8136 : AOI221_X1 port map( B1 => n14163, B2 => n2000, C1 => n14160, C2 => 
                           n6965, A => n3460, ZN => n3459);
   U8137 : NAND4_X1 port map( A1 => n3493, A2 => n3494, A3 => n3495, A4 => 
                           n3496, ZN => n3474);
   U8138 : AOI221_X1 port map( B1 => n14723, B2 => n8145, C1 => n14720, C2 => 
                           n8177, A => n3498, ZN => n3495);
   U8139 : AOI221_X1 port map( B1 => n8303, B2 => n14129, C1 => n8271, C2 => 
                           n14126, A => n3500, ZN => n3493);
   U8140 : AOI221_X1 port map( B1 => n14163, B2 => n1999, C1 => n14160, C2 => 
                           n6979, A => n3497, ZN => n3496);
   U8141 : NAND4_X1 port map( A1 => n3530, A2 => n3531, A3 => n3532, A4 => 
                           n3533, ZN => n3511);
   U8142 : AOI221_X1 port map( B1 => n827, B2 => n14147, C1 => n826, C2 => 
                           n14149, A => n3535, ZN => n3532);
   U8143 : AOI221_X1 port map( B1 => n14144, B2 => n2391, C1 => n14141, C2 => 
                           n1977, A => n3536, ZN => n3531);
   U8144 : AOI221_X1 port map( B1 => n8302, B2 => n14129, C1 => n8270, C2 => 
                           n14126, A => n3537, ZN => n3530);
   U8145 : NAND4_X1 port map( A1 => n3567, A2 => n3568, A3 => n3569, A4 => 
                           n3570, ZN => n3548);
   U8146 : AOI221_X1 port map( B1 => n8301, B2 => n14129, C1 => n8269, C2 => 
                           n14126, A => n3574, ZN => n3567);
   U8147 : AOI221_X1 port map( B1 => n763, B2 => n14147, C1 => n762, C2 => 
                           n14149, A => n3572, ZN => n3569);
   U8148 : AOI221_X1 port map( B1 => n14163, B2 => n761, C1 => n14160, C2 => 
                           n1658, A => n3571, ZN => n3570);
   U8149 : NAND4_X1 port map( A1 => n3604, A2 => n3605, A3 => n3606, A4 => 
                           n3607, ZN => n3585);
   U8150 : AOI221_X1 port map( B1 => n14723, B2 => n8142, C1 => n14720, C2 => 
                           n8174, A => n3609, ZN => n3606);
   U8151 : AOI221_X1 port map( B1 => n8300, B2 => n14128, C1 => n8268, C2 => 
                           n14125, A => n3611, ZN => n3604);
   U8152 : AOI221_X1 port map( B1 => n14162, B2 => n1996, C1 => n14159, C2 => 
                           n7018, A => n3608, ZN => n3607);
   U8153 : NAND4_X1 port map( A1 => n3641, A2 => n3642, A3 => n3643, A4 => 
                           n3644, ZN => n3622);
   U8154 : AOI221_X1 port map( B1 => n14723, B2 => n8141, C1 => n14720, C2 => 
                           n8173, A => n3646, ZN => n3643);
   U8155 : AOI221_X1 port map( B1 => n8299, B2 => n14128, C1 => n8267, C2 => 
                           n14125, A => n3648, ZN => n3641);
   U8156 : AOI221_X1 port map( B1 => n14162, B2 => n1995, C1 => n14159, C2 => 
                           n7032, A => n3645, ZN => n3644);
   U8157 : NAND4_X1 port map( A1 => n3678, A2 => n3679, A3 => n3680, A4 => 
                           n3681, ZN => n3659);
   U8158 : AOI221_X1 port map( B1 => n14723, B2 => n8140, C1 => n14720, C2 => 
                           n8172, A => n3683, ZN => n3680);
   U8159 : AOI221_X1 port map( B1 => n8298, B2 => n14128, C1 => n8266, C2 => 
                           n14125, A => n3685, ZN => n3678);
   U8160 : AOI221_X1 port map( B1 => n14162, B2 => n1994, C1 => n14159, C2 => 
                           n7039, A => n3682, ZN => n3681);
   U8161 : NAND4_X1 port map( A1 => n3715, A2 => n3716, A3 => n3717, A4 => 
                           n3718, ZN => n3696);
   U8162 : AOI221_X1 port map( B1 => n14723, B2 => n8139, C1 => n14720, C2 => 
                           n8171, A => n3720, ZN => n3717);
   U8163 : AOI221_X1 port map( B1 => n8297, B2 => n14128, C1 => n8265, C2 => 
                           n14125, A => n3722, ZN => n3715);
   U8164 : AOI221_X1 port map( B1 => n14162, B2 => n1993, C1 => n14159, C2 => 
                           n7047, A => n3719, ZN => n3718);
   U8165 : NAND4_X1 port map( A1 => n3752, A2 => n3753, A3 => n3754, A4 => 
                           n3755, ZN => n3733);
   U8166 : AOI221_X1 port map( B1 => n14723, B2 => n8138, C1 => n14720, C2 => 
                           n8170, A => n3757, ZN => n3754);
   U8167 : AOI221_X1 port map( B1 => n8296, B2 => n14128, C1 => n8264, C2 => 
                           n14125, A => n3759, ZN => n3752);
   U8168 : AOI221_X1 port map( B1 => n14162, B2 => n1992, C1 => n14159, C2 => 
                           n7056, A => n3756, ZN => n3755);
   U8169 : NAND4_X1 port map( A1 => n3789, A2 => n3790, A3 => n3791, A4 => 
                           n3792, ZN => n3770);
   U8170 : AOI221_X1 port map( B1 => n14723, B2 => n8137, C1 => n14720, C2 => 
                           n8169, A => n3794, ZN => n3791);
   U8171 : AOI221_X1 port map( B1 => n8295, B2 => n14128, C1 => n8263, C2 => 
                           n14125, A => n3796, ZN => n3789);
   U8172 : AOI221_X1 port map( B1 => n14162, B2 => n1991, C1 => n14159, C2 => 
                           n7063, A => n3793, ZN => n3792);
   U8173 : NAND4_X1 port map( A1 => n3826, A2 => n3827, A3 => n3828, A4 => 
                           n3829, ZN => n3807);
   U8174 : AOI221_X1 port map( B1 => n14723, B2 => n8136, C1 => n14720, C2 => 
                           n8168, A => n3831, ZN => n3828);
   U8175 : AOI221_X1 port map( B1 => n8294, B2 => n14128, C1 => n8262, C2 => 
                           n14125, A => n3833, ZN => n3826);
   U8176 : AOI221_X1 port map( B1 => n14162, B2 => n1990, C1 => n14159, C2 => 
                           n7071, A => n3830, ZN => n3829);
   U8177 : NAND4_X1 port map( A1 => n3863, A2 => n3864, A3 => n3865, A4 => 
                           n3866, ZN => n3844);
   U8178 : AOI221_X1 port map( B1 => n14723, B2 => n8135, C1 => n14720, C2 => 
                           n8167, A => n3868, ZN => n3865);
   U8179 : AOI221_X1 port map( B1 => n8293, B2 => n14128, C1 => n8261, C2 => 
                           n14125, A => n3870, ZN => n3863);
   U8180 : AOI221_X1 port map( B1 => n14162, B2 => n1989, C1 => n14159, C2 => 
                           n7080, A => n3867, ZN => n3866);
   U8181 : NAND4_X1 port map( A1 => n3900, A2 => n3901, A3 => n3902, A4 => 
                           n3903, ZN => n3881);
   U8182 : AOI221_X1 port map( B1 => n14723, B2 => n8134, C1 => n14720, C2 => 
                           n8166, A => n3905, ZN => n3902);
   U8183 : AOI221_X1 port map( B1 => n8292, B2 => n14128, C1 => n8260, C2 => 
                           n14125, A => n3907, ZN => n3900);
   U8184 : AOI221_X1 port map( B1 => n14162, B2 => n2406, C1 => n14159, C2 => 
                           n7087, A => n3904, ZN => n3903);
   U8185 : NAND4_X1 port map( A1 => n3937, A2 => n3938, A3 => n3939, A4 => 
                           n3940, ZN => n3918);
   U8186 : AOI221_X1 port map( B1 => n14723, B2 => n8133, C1 => n14720, C2 => 
                           n8165, A => n3942, ZN => n3939);
   U8187 : AOI221_X1 port map( B1 => n8291, B2 => n14128, C1 => n8259, C2 => 
                           n14125, A => n3944, ZN => n3937);
   U8188 : AOI221_X1 port map( B1 => n14162, B2 => n2405, C1 => n14159, C2 => 
                           n7095, A => n3941, ZN => n3940);
   U8189 : NAND4_X1 port map( A1 => n5259, A2 => n5260, A3 => n5261, A4 => 
                           n5262, ZN => n5240);
   U8190 : AOI221_X1 port map( B1 => n14724, B2 => n8132, C1 => n14721, C2 => 
                           n8164, A => n5264, ZN => n5261);
   U8191 : AOI221_X1 port map( B1 => n8290, B2 => n14128, C1 => n8258, C2 => 
                           n14125, A => n5266, ZN => n5259);
   U8192 : AOI221_X1 port map( B1 => n14162, B2 => n2437, C1 => n14159, C2 => 
                           n7104, A => n5263, ZN => n5262);
   U8193 : OAI21_X1 port map( B1 => n13861, B2 => n2241, A => n14944, ZN => 
                           n9042);
   U8194 : OAI21_X1 port map( B1 => n13861, B2 => n2242, A => n14944, ZN => 
                           n9041);
   U8195 : OAI21_X1 port map( B1 => n14081, B2 => n2273, A => n14941, ZN => 
                           n9010);
   U8196 : OAI21_X1 port map( B1 => n14081, B2 => n2274, A => n14941, ZN => 
                           n9009);
   U8197 : OAI21_X1 port map( B1 => n13859, B2 => n2215, A => n14942, ZN => 
                           n9068);
   U8198 : OAI21_X1 port map( B1 => n13859, B2 => n2216, A => n14942, ZN => 
                           n9067);
   U8199 : OAI21_X1 port map( B1 => n13859, B2 => n2217, A => n14942, ZN => 
                           n9066);
   U8200 : OAI21_X1 port map( B1 => n13859, B2 => n2218, A => n14943, ZN => 
                           n9065);
   U8201 : OAI21_X1 port map( B1 => n13859, B2 => n2220, A => n14943, ZN => 
                           n9063);
   U8202 : OAI21_X1 port map( B1 => n13859, B2 => n2221, A => n14943, ZN => 
                           n9062);
   U8203 : OAI21_X1 port map( B1 => n13859, B2 => n2222, A => n14943, ZN => 
                           n9061);
   U8204 : OAI21_X1 port map( B1 => n13859, B2 => n2223, A => n14943, ZN => 
                           n9060);
   U8205 : OAI21_X1 port map( B1 => n13859, B2 => n2224, A => n14943, ZN => 
                           n9059);
   U8206 : OAI21_X1 port map( B1 => n13859, B2 => n2225, A => n14943, ZN => 
                           n9058);
   U8207 : OAI21_X1 port map( B1 => n13859, B2 => n2226, A => n14943, ZN => 
                           n9057);
   U8208 : OAI21_X1 port map( B1 => n13859, B2 => n2227, A => n14943, ZN => 
                           n9056);
   U8209 : OAI21_X1 port map( B1 => n13860, B2 => n2228, A => n14943, ZN => 
                           n9055);
   U8210 : OAI21_X1 port map( B1 => n13860, B2 => n2229, A => n14943, ZN => 
                           n9054);
   U8211 : OAI21_X1 port map( B1 => n13860, B2 => n2230, A => n14943, ZN => 
                           n9053);
   U8212 : OAI21_X1 port map( B1 => n13859, B2 => n2231, A => n14944, ZN => 
                           n9052);
   U8213 : OAI21_X1 port map( B1 => n13860, B2 => n2232, A => n14944, ZN => 
                           n9051);
   U8214 : OAI21_X1 port map( B1 => n13860, B2 => n2233, A => n14944, ZN => 
                           n9050);
   U8215 : OAI21_X1 port map( B1 => n13860, B2 => n2234, A => n14944, ZN => 
                           n9049);
   U8216 : OAI21_X1 port map( B1 => n13860, B2 => n2235, A => n14944, ZN => 
                           n9048);
   U8217 : OAI21_X1 port map( B1 => n13860, B2 => n2236, A => n14944, ZN => 
                           n9047);
   U8218 : OAI21_X1 port map( B1 => n13860, B2 => n2237, A => n14944, ZN => 
                           n9046);
   U8219 : OAI21_X1 port map( B1 => n13860, B2 => n2238, A => n14944, ZN => 
                           n9045);
   U8220 : OAI21_X1 port map( B1 => n13860, B2 => n2239, A => n14944, ZN => 
                           n9044);
   U8221 : OAI21_X1 port map( B1 => n13860, B2 => n2240, A => n14944, ZN => 
                           n9043);
   U8222 : OAI21_X1 port map( B1 => n13860, B2 => n2243, A => n14944, ZN => 
                           n9040);
   U8223 : OAI21_X1 port map( B1 => n14079, B2 => n2247, A => n14945, ZN => 
                           n9036);
   U8224 : OAI21_X1 port map( B1 => n14079, B2 => n2248, A => n14945, ZN => 
                           n9035);
   U8225 : OAI21_X1 port map( B1 => n14079, B2 => n2249, A => n14945, ZN => 
                           n9034);
   U8226 : OAI21_X1 port map( B1 => n14079, B2 => n2250, A => n14945, ZN => 
                           n9033);
   U8227 : OAI21_X1 port map( B1 => n14079, B2 => n2252, A => n14945, ZN => 
                           n9031);
   U8228 : OAI21_X1 port map( B1 => n14079, B2 => n2253, A => n14945, ZN => 
                           n9030);
   U8229 : OAI21_X1 port map( B1 => n14079, B2 => n2254, A => n14945, ZN => 
                           n9029);
   U8230 : OAI21_X1 port map( B1 => n14079, B2 => n2255, A => n14945, ZN => 
                           n9028);
   U8231 : OAI21_X1 port map( B1 => n14079, B2 => n2256, A => n14946, ZN => 
                           n9027);
   U8232 : OAI21_X1 port map( B1 => n14079, B2 => n2257, A => n14946, ZN => 
                           n9026);
   U8233 : OAI21_X1 port map( B1 => n14079, B2 => n2258, A => n14946, ZN => 
                           n9025);
   U8234 : OAI21_X1 port map( B1 => n14079, B2 => n2259, A => n14946, ZN => 
                           n9024);
   U8235 : OAI21_X1 port map( B1 => n14080, B2 => n2260, A => n14946, ZN => 
                           n9023);
   U8236 : OAI21_X1 port map( B1 => n14080, B2 => n2261, A => n14946, ZN => 
                           n9022);
   U8237 : OAI21_X1 port map( B1 => n14080, B2 => n2262, A => n14946, ZN => 
                           n9021);
   U8238 : OAI21_X1 port map( B1 => n14079, B2 => n2263, A => n14946, ZN => 
                           n9020);
   U8239 : OAI21_X1 port map( B1 => n14080, B2 => n2264, A => n14946, ZN => 
                           n9019);
   U8240 : OAI21_X1 port map( B1 => n14080, B2 => n2265, A => n14946, ZN => 
                           n9018);
   U8241 : OAI21_X1 port map( B1 => n14080, B2 => n2266, A => n14946, ZN => 
                           n9017);
   U8242 : OAI21_X1 port map( B1 => n14080, B2 => n2267, A => n14946, ZN => 
                           n9016);
   U8243 : OAI21_X1 port map( B1 => n14080, B2 => n2268, A => n14941, ZN => 
                           n9015);
   U8244 : OAI21_X1 port map( B1 => n14080, B2 => n2269, A => n14946, ZN => 
                           n9014);
   U8245 : OAI21_X1 port map( B1 => n14080, B2 => n2270, A => n14941, ZN => 
                           n9013);
   U8246 : OAI21_X1 port map( B1 => n14080, B2 => n2271, A => ENABLE, ZN => 
                           n9012);
   U8247 : OAI21_X1 port map( B1 => n14080, B2 => n2272, A => n14941, ZN => 
                           n9011);
   U8248 : OAI21_X1 port map( B1 => n14080, B2 => n2275, A => ENABLE, ZN => 
                           n9008);
   U8249 : OAI21_X1 port map( B1 => n13858, B2 => n2214, A => n14945, ZN => 
                           n9069);
   U8250 : OAI21_X1 port map( B1 => n13858, B2 => n2219, A => n14943, ZN => 
                           n9064);
   U8251 : OAI21_X1 port map( B1 => n13858, B2 => n2244, A => n14945, ZN => 
                           n9039);
   U8252 : OAI21_X1 port map( B1 => n13858, B2 => n2245, A => n14945, ZN => 
                           n9038);
   U8253 : OAI21_X1 port map( B1 => n14078, B2 => n2246, A => n14945, ZN => 
                           n9037);
   U8254 : OAI21_X1 port map( B1 => n14078, B2 => n2251, A => n14945, ZN => 
                           n9032);
   U8255 : OAI21_X1 port map( B1 => n14078, B2 => n2276, A => n14941, ZN => 
                           n9007);
   U8256 : OAI21_X1 port map( B1 => n14078, B2 => n2277, A => ENABLE, ZN => 
                           n9006);
   U8257 : NOR3_X2 port map( A1 => n2548, A2 => ADD_RD1(2), A3 => n2547, ZN => 
                           n5195);
   U8258 : NOR3_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n2546, 
                           ZN => n5194);
   U8259 : NOR3_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n2547, 
                           ZN => n5196);
   U8260 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n2553, 
                           ZN => n6515);
   U8261 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n2554, 
                           ZN => n6511);
   U8262 : NOR3_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n2552, 
                           ZN => n6516);
   U8263 : NOR3_X2 port map( A1 => n2554, A2 => ADD_RD2(2), A3 => n2553, ZN => 
                           n6517);
   U8264 : NOR3_X2 port map( A1 => n2547, A2 => ADD_RD1(0), A3 => n2546, ZN => 
                           n5192);
   U8265 : NOR2_X1 port map( A1 => ADD_SF(4), A2 => ADD_SF(5), ZN => n6601);
   U8266 : NOR2_X1 port map( A1 => ADD_SF(1), A2 => ADD_SF(2), ZN => n6572);
   U8267 : NOR2_X1 port map( A1 => n2588, A2 => ADD_SF(2), ZN => n6573);
   U8268 : NOR2_X1 port map( A1 => n2587, A2 => ADD_SF(1), ZN => n6574);
   U8269 : NOR4_X1 port map( A1 => n5233, A2 => n5234, A3 => n5235, A4 => n5236
                           , ZN => n5232);
   U8270 : NOR4_X1 port map( A1 => n6554, A2 => n6555, A3 => n6556, A4 => n6557
                           , ZN => n6553);
   U8271 : NAND2_X1 port map( A1 => RD_Mem, A2 => n14943, ZN => n2748);
   U8272 : NOR2_X1 port map( A1 => n2586, A2 => ADD_SF(0), ZN => n6709);
   U8273 : NOR2_X1 port map( A1 => n2589, A2 => ADD_SF(3), ZN => n6715);
   U8274 : NOR2_X1 port map( A1 => n2532, A2 => ADD_WR(6), ZN => n3953);
   U8275 : NOR2_X1 port map( A1 => ADD_SF(3), A2 => ADD_SF(0), ZN => n6720);
   U8276 : AND3_X1 port map( A1 => n3953, A2 => n2534, A3 => ADD_WR(5), ZN => 
                           n6685);
   U8277 : AND3_X1 port map( A1 => ADD_WR(4), A2 => n3953, A3 => ADD_WR(5), ZN 
                           => n6634);
   U8278 : NOR2_X1 port map( A1 => n2748, A2 => ADD_SF(6), ZN => n6680);
   U8279 : INV_X1 port map( A => ADD_RD1(0), ZN => n2548);
   U8280 : INV_X1 port map( A => ADD_RD1(1), ZN => n2547);
   U8281 : INV_X1 port map( A => ADD_RD2(0), ZN => n2554);
   U8282 : INV_X1 port map( A => ADD_RD1(2), ZN => n2546);
   U8283 : AND2_X1 port map( A1 => ADD_SF(5), A2 => ADD_SF(4), ZN => n6569);
   U8284 : AND2_X1 port map( A1 => ADD_SF(5), A2 => n2569, ZN => n6582);
   U8285 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n14944, ZN => n2649);
   U8286 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n14945, ZN => n2650);
   U8287 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n14946, ZN => n2651);
   U8288 : NAND2_X1 port map( A1 => DATAIN(21), A2 => ENABLE, ZN => n2652);
   U8289 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n14941, ZN => n2653);
   U8290 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n14942, ZN => n2654);
   U8291 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n14943, ZN => n2655);
   U8292 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n14944, ZN => n2656);
   U8293 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n14945, ZN => n2657);
   U8294 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n14946, ZN => n2658);
   U8295 : NAND2_X1 port map( A1 => DATAIN(28), A2 => ENABLE, ZN => n2659);
   U8296 : NAND2_X1 port map( A1 => DATAIN(8), A2 => ENABLE, ZN => n2639);
   U8297 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n14941, ZN => n2640);
   U8298 : NAND2_X1 port map( A1 => DATAIN(10), A2 => ENABLE, ZN => n2641);
   U8299 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n14941, ZN => n2642);
   U8300 : NAND2_X1 port map( A1 => DATAIN(12), A2 => ENABLE, ZN => n2643);
   U8301 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n14941, ZN => n2644);
   U8302 : NAND2_X1 port map( A1 => DATAIN(14), A2 => ENABLE, ZN => n2645);
   U8303 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n14941, ZN => n2646);
   U8304 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n14942, ZN => n2647);
   U8305 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n14942, ZN => n2648);
   U8306 : NAND2_X1 port map( A1 => DATAIN(6), A2 => ENABLE, ZN => n2637);
   U8307 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n14941, ZN => n2638);
   U8308 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n14942, ZN => n2626);
   U8309 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n14942, ZN => n2627);
   U8310 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n14942, ZN => n2631);
   U8311 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n14942, ZN => n2632);
   U8312 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n14942, ZN => n2633);
   U8313 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n14942, ZN => n2634);
   U8314 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n14942, ZN => n2635);
   U8315 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n14942, ZN => n2636);
   U8316 : NAND2_X1 port map( A1 => n14941, A2 => DATAIN(29), ZN => n2623);
   U8317 : INV_X1 port map( A => ADD_RD2(1), ZN => n2553);
   U8318 : INV_X1 port map( A => ADD_RD2(2), ZN => n2552);
   U8319 : NAND2_X1 port map( A1 => n6513, A2 => ADD_RD2(6), ZN => n5370);
   U8320 : INV_X1 port map( A => RESET, ZN => n2521);
   U8321 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n6707);
   U8322 : NAND4_X1 port map( A1 => n5229, A2 => n5230, A3 => n5231, A4 => 
                           n5232, ZN => n3954);
   U8323 : NOR3_X1 port map( A1 => n5237, A2 => n2532, A3 => n2530, ZN => n5231
                           );
   U8324 : NAND4_X1 port map( A1 => n6550, A2 => n6551, A3 => n6552, A4 => 
                           n6553, ZN => n5275);
   U8325 : NOR3_X1 port map( A1 => n6558, A2 => n2532, A3 => n2531, ZN => n6552
                           );
   U8326 : NOR2_X1 port map( A1 => n2538, A2 => ADD_WR(1), ZN => n6724);
   U8327 : NOR2_X1 port map( A1 => n2537, A2 => ADD_WR(0), ZN => n6719);
   U8328 : NOR2_X1 port map( A1 => n2535, A2 => ADD_WR(2), ZN => n6708);
   U8329 : NOR2_X1 port map( A1 => n2536, A2 => ADD_WR(3), ZN => n6713);
   U8330 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(3), ZN => n6736);
   U8331 : NAND2_X1 port map( A1 => n5196, A2 => ADD_RD1(6), ZN => n4052);
   U8332 : NAND2_X1 port map( A1 => n6511, A2 => ADD_RD2(6), ZN => n5374);
   U8333 : NAND2_X1 port map( A1 => n6515, A2 => ADD_RD2(6), ZN => n5375);
   U8334 : NAND2_X1 port map( A1 => n5189, A2 => ADD_RD1(6), ZN => n4045);
   U8335 : AND4_X1 port map( A1 => ADD_WR(6), A2 => WR, A3 => n2534, A4 => 
                           n2533, ZN => n6608);
   U8336 : NAND2_X1 port map( A1 => n5192, A2 => ADD_RD1(6), ZN => n4047);
   U8337 : NAND2_X1 port map( A1 => n6510, A2 => ADD_RD2(6), ZN => n5368);
   U8338 : NAND2_X1 port map( A1 => n5191, A2 => ADD_RD1(6), ZN => n4046);
   U8339 : NAND2_X1 port map( A1 => n5190, A2 => ADD_RD1(6), ZN => n4051);
   U8340 : NAND2_X1 port map( A1 => n6512, A2 => ADD_RD2(6), ZN => n5369);
   U8341 : INV_X1 port map( A => ADD_SF(0), ZN => n2589);
   U8342 : INV_X1 port map( A => ADD_RD1(5), ZN => n2543);
   U8343 : INV_X1 port map( A => ADD_RD2(5), ZN => n2549);
   U8344 : INV_X1 port map( A => ADD_RD1(4), ZN => n2544);
   U8345 : INV_X1 port map( A => ADD_RD2(4), ZN => n2550);
   U8346 : INV_X1 port map( A => ADD_RD1(3), ZN => n2545);
   U8347 : INV_X1 port map( A => ADD_RD2(3), ZN => n2551);
   U8348 : INV_X1 port map( A => ADD_WR(5), ZN => n2533);
   U8349 : INV_X1 port map( A => ADD_WR(1), ZN => n2537);
   U8350 : INV_X1 port map( A => ADD_WR(2), ZN => n2536);
   U8351 : INV_X1 port map( A => ADD_WR(4), ZN => n2534);
   U8352 : AND2_X1 port map( A1 => n6508, A2 => ADD_RD2(6), ZN => n5371);
   U8353 : AND2_X1 port map( A1 => n5187, A2 => ADD_RD1(6), ZN => n4048);
   U8354 : AND3_X1 port map( A1 => n6576, A2 => ADD_SF(0), A3 => ADD_SF(6), ZN 
                           => n2804);
   U8355 : AND3_X1 port map( A1 => n6576, A2 => n2589, A3 => ADD_SF(6), ZN => 
                           n2805);
   U8356 : AND3_X1 port map( A1 => n6573, A2 => n2589, A3 => ADD_SF(6), ZN => 
                           n2799);
   U8357 : AND3_X1 port map( A1 => n6574, A2 => ADD_SF(0), A3 => ADD_SF(6), ZN 
                           => n2798);
   U8358 : INV_X1 port map( A => ADD_SF(4), ZN => n2569);
   U8359 : AND2_X1 port map( A1 => n5195, A2 => ADD_RD1(6), ZN => n4043);
   U8360 : AND2_X1 port map( A1 => n5194, A2 => ADD_RD1(6), ZN => n4042);
   U8361 : AND2_X1 port map( A1 => n6516, A2 => ADD_RD2(6), ZN => n5365);
   U8362 : AND2_X1 port map( A1 => n6517, A2 => ADD_RD2(6), ZN => n5366);
   U8363 : INV_X1 port map( A => WR, ZN => n2532);
   U8364 : NAND2_X1 port map( A1 => WR_Mem, A2 => n14942, ZN => n2778);
   U8365 : INV_X1 port map( A => ADD_WR(3), ZN => n2535);
   U8366 : INV_X1 port map( A => ADD_WR(0), ZN => n2538);
   U8367 : BUF_X1 port map( A => ENABLE, Z => n14941);
   U8368 : INV_X1 port map( A => ADD_SF(1), ZN => n2588);
   U8369 : INV_X1 port map( A => ADD_SF(2), ZN => n2587);
   U8370 : INV_X1 port map( A => ADD_SF(3), ZN => n2586);
   U8371 : INV_X1 port map( A => RD1, ZN => n2530);
   U8372 : INV_X1 port map( A => RD2, ZN => n2531);
   U8373 : INV_X1 port map( A => DATAIN(6), ZN => n2615);
   U8374 : INV_X1 port map( A => DATAIN(20), ZN => n2601);
   U8375 : INV_X1 port map( A => DATAIN(21), ZN => n2600);
   U8376 : INV_X1 port map( A => DATAIN(22), ZN => n2599);
   U8377 : INV_X1 port map( A => DATAIN(23), ZN => n2598);
   U8378 : INV_X1 port map( A => DATAIN(24), ZN => n2597);
   U8379 : INV_X1 port map( A => DATAIN(18), ZN => n2603);
   U8380 : INV_X1 port map( A => DATAIN(19), ZN => n2602);
   U8381 : INV_X1 port map( A => DATAIN(31), ZN => n2590);
   U8382 : INV_X1 port map( A => DATAIN(25), ZN => n2596);
   U8383 : INV_X1 port map( A => DATAIN(26), ZN => n2595);
   U8384 : INV_X1 port map( A => DATAIN(27), ZN => n2594);
   U8385 : INV_X1 port map( A => DATAIN(28), ZN => n2593);
   U8386 : INV_X1 port map( A => DATAIN(29), ZN => n2592);
   U8387 : INV_X1 port map( A => DATAIN(30), ZN => n2591);
   U8388 : INV_X1 port map( A => DATAIN(0), ZN => n2621);
   U8389 : INV_X1 port map( A => DATAIN(1), ZN => n2620);
   U8390 : INV_X1 port map( A => DATAIN(2), ZN => n2619);
   U8391 : INV_X1 port map( A => DATAIN(3), ZN => n2618);
   U8392 : INV_X1 port map( A => DATAIN(4), ZN => n2617);
   U8393 : INV_X1 port map( A => DATAIN(5), ZN => n2616);
   U8394 : INV_X1 port map( A => DATAIN(7), ZN => n2614);
   U8395 : INV_X1 port map( A => DATAIN(8), ZN => n2613);
   U8396 : INV_X1 port map( A => DATAIN(9), ZN => n2612);
   U8397 : INV_X1 port map( A => DATAIN(10), ZN => n2611);
   U8398 : INV_X1 port map( A => DATAIN(11), ZN => n2610);
   U8399 : INV_X1 port map( A => DATAIN(12), ZN => n2609);
   U8400 : INV_X1 port map( A => DATAIN(13), ZN => n2608);
   U8401 : INV_X1 port map( A => DATAIN(14), ZN => n2607);
   U8402 : INV_X1 port map( A => DATAIN(15), ZN => n2606);
   U8403 : INV_X1 port map( A => DATAIN(16), ZN => n2605);
   U8404 : INV_X1 port map( A => DATAIN(17), ZN => n2604);
   U8405 : CLKBUF_X1 port map( A => n5278, Z => n13861);
   U8406 : INV_X1 port map( A => n4093, ZN => n13871);
   U8407 : CLKBUF_X1 port map( A => n3957, Z => n14081);
   U8408 : INV_X1 port map( A => n2847, ZN => n14147);
   U8409 : INV_X1 port map( A => n2846, ZN => n14149);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   port( clk, reset, enable, rd1, rd2, wr, fill, spill : in std_logic;  add_wr,
         add_rd1, add_rd2, add_SF : in std_logic_vector (4 downto 0);  cwp : in
         std_logic_vector (3 downto 0);  add_wr_out, add_rd1_out, add_rd2_out, 
         add_SF_out : out std_logic_vector (6 downto 0));

end translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7;

architecture SYN_beh of 
   translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N52, N53, N76, N77, N164, N165, N221, N222, N239, N240, N241, N242, 
      N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, 
      N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, 
      N267, N268, N269, N270, r239_B_AS_4_port, r239_carry_4_port, 
      r239_carry_5_port, r39_B_AS_4_port, r39_carry_4_port, r39_carry_5_port, 
      r237_B_AS_4_port, r237_carry_4_port, r237_carry_5_port, r238_B_AS_4_port,
      r238_carry_4_port, r238_carry_5_port, n2, n3, n4, n5, n6, n7, n8, n9, n10
      , n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43 : std_logic;

begin
   
   add_SF_outVar_reg_6_inst : DLH_X1 port map( G => N263, D => N270, Q => 
                           add_SF_out(6));
   add_SF_outVar_reg_5_inst : DLH_X1 port map( G => N263, D => N269, Q => 
                           add_SF_out(5));
   add_SF_outVar_reg_4_inst : DLH_X1 port map( G => N263, D => N268, Q => 
                           add_SF_out(4));
   add_SF_outVar_reg_3_inst : DLH_X1 port map( G => N263, D => N267, Q => 
                           add_SF_out(3));
   add_SF_outVar_reg_2_inst : DLH_X1 port map( G => N263, D => N266, Q => 
                           add_SF_out(2));
   add_SF_outVar_reg_1_inst : DLH_X1 port map( G => N263, D => N265, Q => 
                           add_SF_out(1));
   add_SF_outVar_reg_0_inst : DLH_X1 port map( G => N263, D => N264, Q => 
                           add_SF_out(0));
   add_wr_outVar_reg_6_inst : DLH_X1 port map( G => N239, D => N246, Q => 
                           add_wr_out(6));
   add_wr_outVar_reg_5_inst : DLH_X1 port map( G => N239, D => N245, Q => 
                           add_wr_out(5));
   add_wr_outVar_reg_4_inst : DLH_X1 port map( G => N239, D => N244, Q => 
                           add_wr_out(4));
   add_wr_outVar_reg_3_inst : DLH_X1 port map( G => N239, D => N243, Q => 
                           add_wr_out(3));
   add_wr_outVar_reg_2_inst : DLH_X1 port map( G => N239, D => N242, Q => 
                           add_wr_out(2));
   add_wr_outVar_reg_1_inst : DLH_X1 port map( G => N239, D => N241, Q => 
                           add_wr_out(1));
   add_wr_outVar_reg_0_inst : DLH_X1 port map( G => N239, D => N240, Q => 
                           add_wr_out(0));
   add_rd1_outVar_reg_6_inst : DLH_X1 port map( G => N247, D => N254, Q => 
                           add_rd1_out(6));
   add_rd1_outVar_reg_5_inst : DLH_X1 port map( G => N247, D => N253, Q => 
                           add_rd1_out(5));
   add_rd1_outVar_reg_4_inst : DLH_X1 port map( G => N247, D => N252, Q => 
                           add_rd1_out(4));
   add_rd1_outVar_reg_3_inst : DLH_X1 port map( G => N247, D => N251, Q => 
                           add_rd1_out(3));
   add_rd1_outVar_reg_2_inst : DLH_X1 port map( G => N247, D => N250, Q => 
                           add_rd1_out(2));
   add_rd1_outVar_reg_1_inst : DLH_X1 port map( G => N247, D => N249, Q => 
                           add_rd1_out(1));
   add_rd1_outVar_reg_0_inst : DLH_X1 port map( G => N247, D => N248, Q => 
                           add_rd1_out(0));
   add_rd2_outVar_reg_6_inst : DLH_X1 port map( G => N255, D => N262, Q => 
                           add_rd2_out(6));
   add_rd2_outVar_reg_5_inst : DLH_X1 port map( G => N255, D => N261, Q => 
                           add_rd2_out(5));
   add_rd2_outVar_reg_4_inst : DLH_X1 port map( G => N255, D => N260, Q => 
                           add_rd2_out(4));
   add_rd2_outVar_reg_3_inst : DLH_X1 port map( G => N255, D => N259, Q => 
                           add_rd2_out(3));
   add_rd2_outVar_reg_2_inst : DLH_X1 port map( G => N255, D => N258, Q => 
                           add_rd2_out(2));
   add_rd2_outVar_reg_1_inst : DLH_X1 port map( G => N255, D => N257, Q => 
                           add_rd2_out(1));
   add_rd2_outVar_reg_0_inst : DLH_X1 port map( G => N255, D => N256, Q => 
                           add_rd2_out(0));
   r239_U1_3 : FA_X1 port map( A => add_wr(3), B => n2, CI => n36, CO => 
                           r239_carry_4_port, S => N52);
   r239_U1_4 : FA_X1 port map( A => add_wr(4), B => r239_B_AS_4_port, CI => 
                           r239_carry_4_port, CO => r239_carry_5_port, S => N53
                           );
   r39_U1_3 : FA_X1 port map( A => add_SF(3), B => n11, CI => n39, CO => 
                           r39_carry_4_port, S => N221);
   r39_U1_4 : FA_X1 port map( A => add_SF(4), B => r39_B_AS_4_port, CI => 
                           r39_carry_4_port, CO => r39_carry_5_port, S => N222)
                           ;
   r237_U1_3 : FA_X1 port map( A => add_rd1(3), B => n5, CI => n37, CO => 
                           r237_carry_4_port, S => N76);
   r237_U1_4 : FA_X1 port map( A => add_rd1(4), B => r237_B_AS_4_port, CI => 
                           r237_carry_4_port, CO => r237_carry_5_port, S => N77
                           );
   r238_U1_3 : FA_X1 port map( A => add_rd2(3), B => n8, CI => n38, CO => 
                           r238_carry_4_port, S => N164);
   r238_U1_4 : FA_X1 port map( A => add_rd2(4), B => r238_B_AS_4_port, CI => 
                           r238_carry_4_port, CO => r238_carry_5_port, S => 
                           N165);
   U74 : XOR2_X1 port map( A => n20, B => n39, Z => n19);
   U75 : XOR2_X1 port map( A => n25, B => n38, Z => n24);
   U76 : XOR2_X1 port map( A => n29, B => n37, Z => n28);
   U77 : XOR2_X1 port map( A => n33, B => n36, Z => n32);
   U3 : INV_X1 port map( A => n42, ZN => n43);
   U4 : NOR2_X1 port map( A1 => n43, A2 => n26, ZN => N261);
   U5 : XNOR2_X1 port map( A => r238_carry_5_port, B => n9, ZN => n26);
   U6 : NOR2_X1 port map( A1 => n43, A2 => n30, ZN => N253);
   U7 : XNOR2_X1 port map( A => r237_carry_5_port, B => n6, ZN => n30);
   U8 : NOR2_X1 port map( A1 => n43, A2 => n34, ZN => N245);
   U9 : XNOR2_X1 port map( A => r239_carry_5_port, B => n3, ZN => n34);
   U10 : NOR2_X1 port map( A1 => n43, A2 => n22, ZN => N269);
   U11 : XNOR2_X1 port map( A => r39_carry_5_port, B => n12, ZN => n22);
   U12 : NOR2_X1 port map( A1 => n24, A2 => n43, ZN => N262);
   U13 : NAND2_X1 port map( A1 => r238_carry_5_port, A2 => n9, ZN => n25);
   U14 : NOR2_X1 port map( A1 => n28, A2 => n43, ZN => N254);
   U15 : NAND2_X1 port map( A1 => r237_carry_5_port, A2 => n6, ZN => n29);
   U16 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => N246);
   U17 : NAND2_X1 port map( A1 => r239_carry_5_port, A2 => n3, ZN => n33);
   U18 : NOR2_X1 port map( A1 => n19, A2 => n43, ZN => N270);
   U19 : NAND2_X1 port map( A1 => r39_carry_5_port, A2 => n12, ZN => n20);
   U20 : AND2_X1 port map( A1 => N52, A2 => n42, ZN => N243);
   U21 : AND2_X1 port map( A1 => N53, A2 => n42, ZN => N244);
   U22 : AND2_X1 port map( A1 => N164, A2 => n40, ZN => N259);
   U23 : AND2_X1 port map( A1 => N165, A2 => n40, ZN => N260);
   U24 : AND2_X1 port map( A1 => N76, A2 => n41, ZN => N251);
   U25 : AND2_X1 port map( A1 => N77, A2 => n41, ZN => N252);
   U26 : AND2_X1 port map( A1 => N221, A2 => n40, ZN => N267);
   U27 : AND2_X1 port map( A1 => N222, A2 => n40, ZN => N268);
   U28 : NOR2_X1 port map( A1 => n11, A2 => n14, ZN => r39_B_AS_4_port);
   U29 : NOR2_X1 port map( A1 => n8, A2 => n14, ZN => r238_B_AS_4_port);
   U30 : NOR2_X1 port map( A1 => n5, A2 => n14, ZN => r237_B_AS_4_port);
   U31 : NOR2_X1 port map( A1 => n2, A2 => n14, ZN => r239_B_AS_4_port);
   U32 : INV_X1 port map( A => cwp(0), ZN => n14);
   U33 : AND3_X1 port map( A1 => add_SF(4), A2 => n13, A3 => n21, ZN => n39);
   U34 : INV_X1 port map( A => add_SF(3), ZN => n13);
   U35 : BUF_X1 port map( A => enable, Z => n42);
   U36 : AND3_X1 port map( A1 => n21, A2 => n10, A3 => add_rd2(4), ZN => n38);
   U37 : INV_X1 port map( A => add_rd2(3), ZN => n10);
   U38 : AND3_X1 port map( A1 => n21, A2 => n7, A3 => add_rd1(4), ZN => n37);
   U39 : INV_X1 port map( A => add_rd1(3), ZN => n7);
   U40 : AND3_X1 port map( A1 => n21, A2 => n4, A3 => add_wr(4), ZN => n36);
   U41 : INV_X1 port map( A => add_wr(3), ZN => n4);
   U42 : BUF_X1 port map( A => enable, Z => n41);
   U43 : BUF_X1 port map( A => enable, Z => n40);
   U44 : OR2_X1 port map( A1 => rd2, A2 => n43, ZN => N255);
   U45 : OR2_X1 port map( A1 => rd1, A2 => n43, ZN => N247);
   U46 : OR2_X1 port map( A1 => wr, A2 => n43, ZN => N239);
   U47 : AND2_X1 port map( A1 => cwp(1), A2 => cwp(0), ZN => n21);
   U48 : INV_X1 port map( A => n27, ZN => n9);
   U49 : AOI21_X1 port map( B1 => add_rd2(4), B2 => add_rd2(3), A => cwp(1), ZN
                           => n27);
   U50 : INV_X1 port map( A => n31, ZN => n6);
   U51 : AOI21_X1 port map( B1 => add_rd1(3), B2 => add_rd1(4), A => cwp(1), ZN
                           => n31);
   U52 : INV_X1 port map( A => n35, ZN => n3);
   U53 : AOI21_X1 port map( B1 => add_wr(4), B2 => add_wr(3), A => cwp(1), ZN 
                           => n35);
   U54 : INV_X1 port map( A => n23, ZN => n12);
   U55 : AOI21_X1 port map( B1 => add_SF(4), B2 => add_SF(3), A => cwp(1), ZN 
                           => n23);
   U56 : OR3_X1 port map( A1 => spill, A2 => fill, A3 => n43, ZN => N263);
   U57 : INV_X1 port map( A => n15, ZN => n11);
   U58 : AOI21_X1 port map( B1 => add_SF(4), B2 => add_SF(3), A => n39, ZN => 
                           n15);
   U59 : INV_X1 port map( A => n17, ZN => n8);
   U60 : AOI21_X1 port map( B1 => add_rd2(4), B2 => add_rd2(3), A => n38, ZN =>
                           n17);
   U61 : INV_X1 port map( A => n18, ZN => n5);
   U62 : AOI21_X1 port map( B1 => add_rd1(3), B2 => add_rd1(4), A => n37, ZN =>
                           n18);
   U63 : INV_X1 port map( A => n16, ZN => n2);
   U64 : AOI21_X1 port map( B1 => add_wr(4), B2 => add_wr(3), A => n36, ZN => 
                           n16);
   U65 : AND2_X1 port map( A1 => add_rd1(0), A2 => n42, ZN => N248);
   U66 : AND2_X1 port map( A1 => add_wr(0), A2 => n42, ZN => N240);
   U67 : AND2_X1 port map( A1 => add_wr(1), A2 => n42, ZN => N241);
   U68 : AND2_X1 port map( A1 => add_wr(2), A2 => n42, ZN => N242);
   U69 : AND2_X1 port map( A1 => add_rd2(0), A2 => n41, ZN => N256);
   U70 : AND2_X1 port map( A1 => add_rd2(1), A2 => n41, ZN => N257);
   U71 : AND2_X1 port map( A1 => add_rd2(2), A2 => n41, ZN => N258);
   U72 : AND2_X1 port map( A1 => add_rd1(1), A2 => n41, ZN => N249);
   U73 : AND2_X1 port map( A1 => add_rd1(2), A2 => n41, ZN => N250);
   U78 : AND2_X1 port map( A1 => add_SF(0), A2 => n40, ZN => N264);
   U79 : AND2_X1 port map( A1 => add_SF(1), A2 => n40, ZN => N265);
   U80 : AND2_X1 port map( A1 => add_SF(2), A2 => n40, ZN => N266);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
         std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, spill
         , RD_Mem, WR_Mem : out std_logic;  add_SF : out std_logic_vector (4 
         downto 0);  MMUStrobe : in std_logic;  dataACK : out std_logic);

end controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5;

architecture SYN_beh of 
   controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port, 
      swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port, 
      need_to_fill_0_port, need_to_spill_0_port, nextState_2_port, 
      nextState_1_port, nextState_0_port, cansaveNext_3_port, 
      cansaveNext_2_port, cansaveNext_1_port, cansaveNext_0_port, 
      canrestoreNext_3_port, canrestoreNext_2_port, canrestoreNext_1_port, 
      canrestoreNext_0_port, oldCWP_3_port, oldCWP_2_port, oldCWP_1_port, 
      oldCWP_0_port, regCntNext_4_port, regCntNext_3_port, regCntNext_2_port, 
      regCntNext_1_port, regCntNext_0_port, regCnt_4_port, regCnt_3_port, 
      regCnt_2_port, regCnt_1_port, regCnt_0_port, N418, N420, N422, N424, N426
      , N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
      N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, 
      N451, N452, N453, N454, N455, N456, N457, N463, N464, N465, N466, N467, 
      n227, n234, n235, n6, n7, n29, n49, n53, n56, n58, n60, n65, n223, n224, 
      n1, n2, n3, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n50, n51, n52, n54, n55, n57, n59, n61, n62, n63, n64, n66, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n225, n226, n_1782, n_1783, n_1784 : std_logic;

begin
   cwpOut <= ( cwpOut_3_port, cwpOut_2_port, cwpOut_1_port, cwpOut_0_port );
   swpOut <= ( swpOut_3_port, swpOut_2_port, swpOut_1_port, swpOut_0_port );
   
   cansaveNext_reg_3_inst : DLH_X1 port map( G => N428, D => N432, Q => 
                           cansaveNext_3_port);
   cwp_reg_3_inst : DLH_X1 port map( G => N441, D => N445, Q => cwpOut_3_port);
   canrestoreNext_reg_3_inst : DLH_X1 port map( G => N428, D => N440, Q => 
                           canrestoreNext_3_port);
   nextState_reg_2_inst : DLH_X1 port map( G => N433, D => N436, Q => 
                           nextState_2_port);
   nextState_reg_1_inst : DLH_X1 port map( G => N433, D => N435, Q => 
                           nextState_1_port);
   oldCWP_reg_0_inst : DLH_X1 port map( G => N451, D => N452, Q => 
                           oldCWP_0_port);
   cansaveNext_reg_2_inst : DLH_X1 port map( G => N428, D => N431, Q => 
                           cansaveNext_2_port);
   nextState_reg_0_inst : DLH_X1 port map( G => N433, D => N434, Q => 
                           nextState_0_port);
   need_to_fill_reg_0_inst : DLH_X1 port map( G => N418, D => n43, Q => 
                           need_to_fill_0_port);
   need_to_spill_reg_0_inst : DLH_X1 port map( G => N420, D => n221, Q => 
                           need_to_spill_0_port);
   WR_Mem_reg : DLH_X1 port map( G => N427, D => n225, Q => WR_Mem);
   swp_reg_3_inst : DLH_X1 port map( G => N446, D => N450, Q => swpOut_3_port);
   swp_reg_2_inst : DLH_X1 port map( G => N446, D => N449, Q => swpOut_2_port);
   swp_reg_0_inst : DLH_X1 port map( G => N446, D => N447, Q => swpOut_0_port);
   add_SF_reg_0_inst : DLH_X1 port map( G => N456, D => N457, Q => add_SF(0));
   RD_Mem_reg : DLH_X1 port map( G => N426, D => n226, Q => RD_Mem);
   cansaveNext_reg_0_inst : DLH_X1 port map( G => N428, D => N429, Q => 
                           cansaveNext_0_port);
   canrestoreNext_reg_0_inst : DLH_X1 port map( G => N428, D => N437, Q => 
                           canrestoreNext_0_port);
   cwp_reg_0_inst : DLH_X1 port map( G => N441, D => N442, Q => cwpOut_0_port);
   oldCWP_reg_1_inst : DLH_X1 port map( G => N451, D => N453, Q => 
                           oldCWP_1_port);
   cansaveNext_reg_1_inst : DLH_X1 port map( G => N428, D => N430, Q => 
                           cansaveNext_1_port);
   swp_reg_1_inst : DLH_X1 port map( G => N446, D => N448, Q => swpOut_1_port);
   canrestoreNext_reg_1_inst : DLH_X1 port map( G => N428, D => N438, Q => 
                           canrestoreNext_1_port);
   cwp_reg_1_inst : DLH_X1 port map( G => N441, D => N443, Q => cwpOut_1_port);
   canrestoreNext_reg_2_inst : DLH_X1 port map( G => N428, D => N439, Q => 
                           canrestoreNext_2_port);
   cwp_reg_2_inst : DLH_X1 port map( G => N441, D => N444, Q => cwpOut_2_port);
   oldCWP_reg_2_inst : DLH_X1 port map( G => N451, D => N454, Q => 
                           oldCWP_2_port);
   oldCWP_reg_3_inst : DLH_X1 port map( G => N451, D => N455, Q => 
                           oldCWP_3_port);
   regCntNext_reg_4_inst : DLH_X1 port map( G => n224, D => N467, Q => 
                           regCntNext_4_port);
   regCntNext_reg_0_inst : DLH_X1 port map( G => n224, D => N463, Q => 
                           regCntNext_0_port);
   regCntNext_reg_1_inst : DLH_X1 port map( G => n224, D => N464, Q => 
                           regCntNext_1_port);
   add_SF_reg_1_inst : DLH_X1 port map( G => N456, D => n222, Q => add_SF(1));
   regCntNext_reg_2_inst : DLH_X1 port map( G => n224, D => N465, Q => 
                           regCntNext_2_port);
   add_SF_reg_2_inst : DLH_X1 port map( G => N456, D => n219, Q => add_SF(2));
   regCntNext_reg_3_inst : DLH_X1 port map( G => n224, D => N466, Q => 
                           regCntNext_3_port);
   add_SF_reg_3_inst : DLH_X1 port map( G => N456, D => n220, Q => add_SF(3));
   add_SF_reg_4_inst : DLH_X1 port map( G => N456, D => n218, Q => add_SF(4));
   fill_reg : DLH_X1 port map( G => N422, D => N424, Q => fill);
   spill_reg : DLH_X1 port map( G => N422, D => n223, Q => spill);
   dataACK <= '0';
   U159 : NOR2_X2 port map( A1 => n226, A2 => n225, ZN => n112);
   U171 : NOR4_X2 port map( A1 => n46, A2 => n29, A3 => n58, A4 => n7, ZN => 
                           n99);
   U250 : XOR2_X1 port map( A => n142, B => n143, Z => n124);
   U251 : XOR2_X1 port map( A => n155, B => n148, Z => n127);
   U252 : XOR2_X1 port map( A => n156, B => n160, Z => n130);
   U253 : NAND3_X1 port map( A1 => n176, A2 => n85, A3 => call, ZN => n175);
   U254 : NAND3_X1 port map( A1 => n98, A2 => call, A3 => n17, ZN => n173);
   U255 : NAND3_X1 port map( A1 => n57, A2 => n18, A3 => need_to_fill_0_port, 
                           ZN => n172);
   U256 : NAND3_X1 port map( A1 => n118, A2 => n42, A3 => n11, ZN => N428);
   U257 : OAI33_X1 port map( A1 => n167, A2 => n69, A3 => n85, B1 => n206, B2 
                           => n179, B3 => n163, ZN => n137);
   U258 : NAND3_X1 port map( A1 => n171, A2 => n18, A3 => need_to_fill_0_port, 
                           ZN => n208);
   U259 : NAND3_X1 port map( A1 => n70, A2 => n64, A3 => n118, ZN => N427);
   U260 : NAND3_X1 port map( A1 => n79, A2 => n81, A3 => n49, ZN => n163);
   U261 : NAND3_X1 port map( A1 => n70, A2 => n68, A3 => n118, ZN => N426);
   regCnt_reg_4_inst : DFF_X1 port map( D => n30, CK => clk, Q => regCnt_4_port
                           , QN => n40);
   regCnt_reg_2_inst : DFF_X1 port map( D => n33, CK => clk, Q => regCnt_2_port
                           , QN => n50);
   regCnt_reg_1_inst : DFF_X1 port map( D => n32, CK => clk, Q => regCnt_1_port
                           , QN => n72);
   regCnt_reg_3_inst : DFF_X1 port map( D => n34, CK => clk, Q => regCnt_3_port
                           , QN => n52);
   cansave_reg_0_inst : DFF_X1 port map( D => n235, CK => clk, Q => n56, QN => 
                           n78);
   cansave_reg_1_inst : DFF_X1 port map( D => n234, CK => clk, Q => n60, QN => 
                           n77);
   canrestore_reg_3_inst : DFF_X1 port map( D => n3, CK => clk, Q => n29, QN =>
                           n_1782);
   canrestore_reg_0_inst : DFF_X1 port map( D => n19, CK => clk, Q => n58, QN 
                           => n_1783);
   canrestore_reg_1_inst : DFF_X1 port map( D => n24, CK => clk, Q => n7, QN =>
                           n_1784);
   regCnt_reg_0_inst : DFF_X1 port map( D => n31, CK => clk, Q => regCnt_0_port
                           , QN => n76);
   currentState_reg_0_inst : DFF_X1 port map( D => n227, CK => clk, Q => n53, 
                           QN => n79);
   cansave_reg_2_inst : DFF_X1 port map( D => n216, CK => clk, Q => n73, QN => 
                           n213);
   canrestore_reg_2_inst : DFF_X1 port map( D => n217, CK => clk, Q => n46, QN 
                           => n65);
   currentState_reg_1_inst : DFF_X1 port map( D => n215, CK => clk, Q => n81, 
                           QN => n6);
   currentState_reg_2_inst : DFF_X1 port map( D => n214, CK => clk, Q => n71, 
                           QN => n49);
   cansave_reg_3_inst : DFF_X1 port map( D => n1, CK => clk, Q => n80, QN => 
                           n212);
   U3 : NOR4_X1 port map( A1 => call, A2 => regCnt_0_port, A3 => n40, A4 => 
                           n209, ZN => n104);
   U4 : NOR3_X1 port map( A1 => n79, A2 => n6, A3 => n71, ZN => n98);
   U5 : INV_X1 port map( A => n191, ZN => n37);
   U6 : NAND2_X1 port map( A1 => n44, A2 => n59, ZN => N441);
   U7 : NOR2_X1 port map( A1 => n68, A2 => n38, ZN => n191);
   U8 : INV_X1 port map( A => n145, ZN => n42);
   U9 : INV_X1 port map( A => n137, ZN => n16);
   U10 : OAI222_X1 port map( A1 => n123, A2 => n127, B1 => n128, B2 => n103, C1
                           => n122, C2 => n129, ZN => N444);
   U11 : OAI222_X1 port map( A1 => n123, A2 => n130, B1 => n103, B2 => n131, C1
                           => n122, C2 => n132, ZN => N443);
   U12 : OAI222_X1 port map( A1 => n123, A2 => n21, B1 => n14, B2 => n103, C1 
                           => n122, C2 => n8, ZN => N442);
   U13 : INV_X1 port map( A => n122, ZN => n35);
   U14 : INV_X1 port map( A => n112, ZN => n61);
   U15 : NAND2_X1 port map( A1 => n61, A2 => n38, ZN => n103);
   U16 : OAI22_X1 port map( A1 => n42, A2 => n130, B1 => n133, B2 => n131, ZN 
                           => N438);
   U17 : OAI22_X1 port map( A1 => n42, A2 => n127, B1 => n133, B2 => n128, ZN 
                           => N439);
   U18 : OAI22_X1 port map( A1 => n42, A2 => n21, B1 => n133, B2 => n14, ZN => 
                           N437);
   U19 : OAI22_X1 port map( A1 => n129, A2 => n42, B1 => n133, B2 => n120, ZN 
                           => N431);
   U20 : NAND4_X1 port map( A1 => n123, A2 => n55, A3 => n70, A4 => n59, ZN => 
                           N422);
   U21 : INV_X1 port map( A => n147, ZN => n41);
   U22 : INV_X1 port map( A => N456, ZN => n59);
   U23 : INV_X1 port map( A => n183, ZN => n36);
   U24 : INV_X1 port map( A => n144, ZN => n44);
   U25 : INV_X1 port map( A => n111, ZN => n48);
   U26 : AND2_X1 port map( A1 => n190, A2 => n28, ZN => n192);
   U27 : NAND2_X1 port map( A1 => n164, A2 => n18, ZN => n206);
   U28 : NOR3_X2 port map( A1 => n70, A2 => n99, A3 => n179, ZN => n145);
   U29 : AOI21_X1 port map( B1 => n225, B2 => n104, A => n191, ZN => n122);
   U30 : NOR3_X1 port map( A1 => n72, A2 => n50, A3 => n76, ZN => n111);
   U31 : NOR3_X1 port map( A1 => n45, A2 => n70, A3 => n179, ZN => n100);
   U32 : NOR2_X1 port map( A1 => n98, A2 => n66, ZN => n123);
   U33 : NOR2_X1 port map( A1 => n168, A2 => n98, ZN => n117);
   U34 : OAI21_X1 port map( B1 => n204, B2 => n162, A => n37, ZN => n183);
   U35 : INV_X1 port map( A => n87, ZN => n82);
   U36 : OAI21_X1 port map( B1 => n204, B2 => n162, A => n16, ZN => n138);
   U37 : XNOR2_X1 port map( A => n149, B => n147, ZN => n155);
   U38 : XNOR2_X1 port map( A => n41, B => n21, ZN => n160);
   U39 : OAI21_X1 port map( B1 => n162, B2 => n163, A => n161, ZN => n144);
   U40 : OAI222_X1 port map( A1 => n123, A2 => n124, B1 => n125, B2 => n103, C1
                           => n122, C2 => n126, ZN => N445);
   U41 : XNOR2_X1 port map( A => n137, B => n159, ZN => n131);
   U42 : XNOR2_X1 port map( A => n14, B => n153, ZN => n159);
   U43 : INV_X1 port map( A => n138, ZN => n11);
   U44 : NAND2_X1 port map( A1 => n112, A2 => n118, ZN => N456);
   U45 : INV_X1 port map( A => n89, ZN => n83);
   U46 : AND2_X1 port map( A1 => n123, A2 => n205, ZN => n133);
   U47 : OAI21_X1 port map( B1 => n99, B2 => n179, A => n176, ZN => n205);
   U48 : AOI21_X1 port map( B1 => n85, B2 => n176, A => n66, ZN => n204);
   U49 : OAI21_X1 port map( B1 => n183, B2 => n13, A => n195, ZN => n185);
   U50 : INV_X1 port map( A => n196, ZN => n13);
   U51 : OAI21_X1 port map( B1 => n196, B2 => n36, A => n197, ZN => n195);
   U52 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n152, ZN => n140);
   U53 : INV_X1 port map( A => n153, ZN => n15);
   U54 : OAI21_X1 port map( B1 => n153, B2 => n154, A => n16, ZN => n152);
   U55 : OAI21_X1 port map( B1 => n199, B2 => n200, A => n201, ZN => n190);
   U56 : OAI21_X1 port map( B1 => n23, B2 => n8, A => n191, ZN => n201);
   U57 : NOR3_X1 port map( A1 => n163, A2 => n74, A3 => n18, ZN => n169);
   U58 : OAI221_X1 port map( B1 => n133, B2 => n121, C1 => n132, C2 => n42, A 
                           => n118, ZN => N430);
   U59 : OAI221_X1 port map( B1 => n133, B2 => n12, C1 => n42, C2 => n8, A => 
                           n118, ZN => N429);
   U60 : OAI21_X1 port map( B1 => n41, B2 => n156, A => n22, ZN => n148);
   U61 : INV_X1 port map( A => n157, ZN => n22);
   U62 : AOI21_X1 port map( B1 => n156, B2 => n41, A => n158, ZN => n157);
   U63 : INV_X1 port map( A => n99, ZN => n45);
   U64 : XNOR2_X1 port map( A => n134, B => n135, ZN => n125);
   U65 : OAI22_X1 port map( A1 => n139, A2 => n140, B1 => n16, B2 => n141, ZN 
                           => n134);
   U66 : XNOR2_X1 port map( A => n136, B => n137, ZN => n135);
   U67 : AND2_X1 port map( A1 => n140, A2 => n139, ZN => n141);
   U68 : OAI211_X1 port map( C1 => n17, C2 => n69, A => n118, B => n55, ZN => 
                           N451);
   U69 : XNOR2_X1 port map( A => n194, B => n185, ZN => n120);
   U70 : XNOR2_X1 port map( A => n36, B => n184, ZN => n194);
   U71 : XNOR2_X1 port map( A => n183, B => n203, ZN => n121);
   U72 : XNOR2_X1 port map( A => n12, B => n196, ZN => n203);
   U73 : XNOR2_X1 port map( A => n151, B => n140, ZN => n128);
   U74 : XNOR2_X1 port map( A => n16, B => n139, ZN => n151);
   U75 : NAND2_X1 port map( A1 => n42, A2 => n161, ZN => n147);
   U76 : XNOR2_X1 port map( A => n198, B => n190, ZN => n129);
   U77 : XNOR2_X1 port map( A => n193, B => n191, ZN => n198);
   U78 : INV_X1 port map( A => n104, ZN => n38);
   U79 : OAI21_X1 port map( B1 => n101, B2 => n102, A => n103, ZN => n224);
   U80 : OAI21_X1 port map( B1 => n112, B2 => n121, A => n118, ZN => N448);
   U81 : OAI21_X1 port map( B1 => n112, B2 => n12, A => n118, ZN => N447);
   U82 : OAI21_X1 port map( B1 => n112, B2 => n120, A => n118, ZN => N449);
   U83 : OAI21_X1 port map( B1 => n112, B2 => n119, A => n118, ZN => N450);
   U84 : XNOR2_X1 port map( A => n191, B => n202, ZN => n132);
   U85 : XNOR2_X1 port map( A => n199, B => n23, ZN => n202);
   U86 : NOR2_X1 port map( A1 => n40, A2 => n112, ZN => n218);
   U87 : NOR2_X1 port map( A1 => n52, A2 => n112, ZN => n220);
   U88 : NOR2_X1 port map( A1 => n50, A2 => n112, ZN => n219);
   U89 : NOR2_X1 port map( A1 => n72, A2 => n112, ZN => n222);
   U90 : OAI22_X1 port map( A1 => n124, A2 => n42, B1 => n133, B2 => n125, ZN 
                           => N440);
   U91 : OAI22_X1 port map( A1 => n42, A2 => n126, B1 => n133, B2 => n119, ZN 
                           => N432);
   U92 : OAI22_X1 port map( A1 => n114, A2 => n47, B1 => n62, B2 => n115, ZN =>
                           N465);
   U93 : INV_X1 port map( A => n222, ZN => n62);
   U94 : INV_X1 port map( A => n219, ZN => n47);
   U95 : NOR2_X1 port map( A1 => n72, A2 => n76, ZN => n114);
   U96 : OAI22_X1 port map( A1 => n109, A2 => n39, B1 => n51, B2 => n110, ZN =>
                           N467);
   U97 : INV_X1 port map( A => n220, ZN => n51);
   U98 : INV_X1 port map( A => n218, ZN => n39);
   U99 : NOR2_X1 port map( A1 => n52, A2 => n48, ZN => n109);
   U100 : OAI22_X1 port map( A1 => n104, A2 => n64, B1 => n54, B2 => n18, ZN =>
                           n223);
   U101 : INV_X1 port map( A => n176, ZN => n70);
   U102 : INV_X1 port map( A => n98, ZN => n69);
   U103 : INV_X1 port map( A => n163, ZN => n66);
   U104 : NOR2_X1 port map( A1 => n112, A2 => n76, ZN => N457);
   U105 : NAND2_X1 port map( A1 => n122, A2 => n118, ZN => N446);
   U106 : INV_X1 port map( A => n154, ZN => n14);
   U107 : NAND2_X1 port map( A1 => n89, A2 => n82, ZN => n94);
   U108 : OAI21_X1 port map( B1 => n210, B2 => n163, A => n63, ZN => N420);
   U109 : INV_X1 port map( A => N427, ZN => n63);
   U110 : NOR2_X1 port map( A1 => n74, A2 => n75, ZN => n210);
   U111 : INV_X1 port map( A => n164, ZN => n75);
   U112 : INV_X1 port map( A => n168, ZN => n55);
   U113 : INV_X1 port map( A => n158, ZN => n21);
   U114 : INV_X1 port map( A => n199, ZN => n8);
   U115 : INV_X1 port map( A => n197, ZN => n12);
   U116 : INV_X1 port map( A => n226, ZN => n68);
   U117 : INV_X1 port map( A => n225, ZN => n64);
   U118 : INV_X1 port map( A => n162, ZN => n74);
   U119 : NAND2_X1 port map( A1 => n111, A2 => n40, ZN => n110);
   U120 : NAND4_X1 port map( A1 => n103, A2 => n54, A3 => n165, A4 => n166, ZN 
                           => N436);
   U121 : NOR2_X1 port map( A1 => n221, A2 => n100, ZN => n165);
   U122 : AOI221_X1 port map( B1 => n98, B2 => n167, C1 => n168, C2 => n10, A 
                           => n169, ZN => n166);
   U123 : INV_X1 port map( A => n101, ZN => n10);
   U124 : INV_X1 port map( A => n200, ZN => n23);
   U125 : NOR2_X1 port map( A1 => n117, A2 => n27, ZN => N454);
   U126 : INV_X1 port map( A => n193, ZN => n28);
   U127 : INV_X1 port map( A => n171, ZN => n54);
   U128 : INV_X1 port map( A => n102, ZN => n57);
   U129 : AND2_X1 port map( A1 => n75, A2 => n170, ZN => n221);
   U130 : INV_X1 port map( A => n167, ZN => n17);
   U131 : AND2_X1 port map( A1 => n185, A2 => n184, ZN => n186);
   U132 : AND2_X1 port map( A1 => n148, A2 => n149, ZN => n150);
   U133 : INV_X1 port map( A => n97, ZN => n43);
   U134 : AOI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n97);
   U135 : OAI22_X1 port map( A1 => n89, A2 => n4, B1 => n49, B2 => n82, ZN => 
                           n214);
   U136 : INV_X1 port map( A => nextState_2_port, ZN => n4);
   U137 : OAI22_X1 port map( A1 => n89, A2 => n5, B1 => n6, B2 => n82, ZN => 
                           n215);
   U138 : INV_X1 port map( A => nextState_1_port, ZN => n5);
   U139 : OAI22_X1 port map( A1 => n89, A2 => n9, B1 => n213, B2 => n82, ZN => 
                           n216);
   U140 : INV_X1 port map( A => cansaveNext_2_port, ZN => n9);
   U141 : OAI22_X1 port map( A1 => n89, A2 => n26, B1 => n65, B2 => n82, ZN => 
                           n217);
   U142 : INV_X1 port map( A => canrestoreNext_2_port, ZN => n26);
   U143 : INV_X1 port map( A => n91, ZN => n24);
   U144 : AOI22_X1 port map( A1 => n83, A2 => canrestoreNext_1_port, B1 => n87,
                           B2 => n7, ZN => n91);
   U145 : OAI211_X1 port map( C1 => n82, C2 => n79, A => n96, B => n94, ZN => 
                           n227);
   U146 : NAND2_X1 port map( A1 => nextState_0_port, A2 => n82, ZN => n96);
   U147 : OAI211_X1 port map( C1 => n82, C2 => n78, A => n93, B => n94, ZN => 
                           n235);
   U148 : NAND2_X1 port map( A1 => cansaveNext_0_port, A2 => n82, ZN => n93);
   U149 : OAI211_X1 port map( C1 => n82, C2 => n77, A => n95, B => n94, ZN => 
                           n234);
   U150 : NAND2_X1 port map( A1 => cansaveNext_1_port, A2 => n82, ZN => n95);
   U151 : INV_X1 port map( A => n90, ZN => n19);
   U152 : AOI22_X1 port map( A1 => n83, A2 => canrestoreNext_0_port, B1 => n87,
                           B2 => n58, ZN => n90);
   U153 : INV_X1 port map( A => n88, ZN => n3);
   U154 : AOI22_X1 port map( A1 => n83, A2 => canrestoreNext_3_port, B1 => n87,
                           B2 => n29, ZN => n88);
   U155 : INV_X1 port map( A => n105, ZN => n31);
   U156 : AOI22_X1 port map( A1 => n89, A2 => regCnt_0_port, B1 => n83, B2 => 
                           regCntNext_0_port, ZN => n105);
   U157 : INV_X1 port map( A => n107, ZN => n32);
   U158 : AOI22_X1 port map( A1 => n89, A2 => regCnt_1_port, B1 => n83, B2 => 
                           regCntNext_1_port, ZN => n107);
   U160 : INV_X1 port map( A => n92, ZN => n34);
   U161 : AOI22_X1 port map( A1 => n89, A2 => regCnt_3_port, B1 => n83, B2 => 
                           regCntNext_3_port, ZN => n92);
   U162 : INV_X1 port map( A => n106, ZN => n33);
   U163 : AOI22_X1 port map( A1 => n89, A2 => regCnt_2_port, B1 => n83, B2 => 
                           regCntNext_2_port, ZN => n106);
   U164 : INV_X1 port map( A => n108, ZN => n30);
   U165 : AOI22_X1 port map( A1 => n89, A2 => regCnt_4_port, B1 => n83, B2 => 
                           regCntNext_4_port, ZN => n108);
   U166 : INV_X1 port map( A => n86, ZN => n1);
   U167 : AOI22_X1 port map( A1 => n83, A2 => cansaveNext_3_port, B1 => n80, B2
                           => n87, ZN => n86);
   U168 : NAND4_X1 port map( A1 => n85, A2 => n52, A3 => n50, A4 => n72, ZN => 
                           n209);
   U169 : NOR3_X1 port map( A1 => n79, A2 => n49, A3 => n81, ZN => n225);
   U170 : NOR3_X1 port map( A1 => n49, A2 => n53, A3 => n81, ZN => n168);
   U172 : NAND3_X1 port map( A1 => n6, A2 => n53, A3 => n49, ZN => n118);
   U173 : NOR3_X1 port map( A1 => n81, A2 => n53, A3 => n71, ZN => n176);
   U174 : NOR3_X1 port map( A1 => n53, A2 => n6, A3 => n49, ZN => n226);
   U175 : NAND2_X1 port map( A1 => enable, A2 => n84, ZN => n89);
   U176 : NOR2_X1 port map( A1 => enable, A2 => reset, ZN => n87);
   U177 : OAI22_X1 port map( A1 => n65, A2 => n42, B1 => n44, B2 => n27, ZN => 
                           n149);
   U178 : AOI22_X1 port map( A1 => n61, A2 => swpOut_1_port, B1 => n138, B2 => 
                           n7, ZN => n153);
   U179 : AOI22_X1 port map( A1 => n35, A2 => swpOut_1_port, B1 => n138, B2 => 
                           n60, ZN => n196);
   U180 : XNOR2_X1 port map( A => n146, B => n147, ZN => n142);
   U181 : AOI22_X1 port map( A1 => cwpOut_3_port, A2 => n144, B1 => n145, B2 =>
                           n29, ZN => n143);
   U182 : OAI22_X1 port map( A1 => n148, A2 => n149, B1 => n150, B2 => n147, ZN
                           => n146);
   U183 : AOI22_X1 port map( A1 => n35, A2 => oldCWP_0_port, B1 => n56, B2 => 
                           n145, ZN => n199);
   U184 : NAND4_X1 port map( A1 => n212, A2 => n213, A3 => n78, A4 => n77, ZN 
                           => n164);
   U185 : AOI22_X1 port map( A1 => n61, A2 => swpOut_2_port, B1 => n138, B2 => 
                           n46, ZN => n139);
   U186 : AOI22_X1 port map( A1 => n35, A2 => swpOut_2_port, B1 => n138, B2 => 
                           n73, ZN => n184);
   U187 : AOI22_X1 port map( A1 => n7, A2 => n145, B1 => n144, B2 => 
                           cwpOut_1_port, ZN => n156);
   U188 : AOI22_X1 port map( A1 => n35, A2 => oldCWP_2_port, B1 => n73, B2 => 
                           n145, ZN => n193);
   U189 : AOI22_X1 port map( A1 => n35, A2 => oldCWP_1_port, B1 => n60, B2 => 
                           n145, ZN => n200);
   U190 : NAND4_X1 port map( A1 => ret, A2 => n98, A3 => n45, A4 => n164, ZN =>
                           n161);
   U191 : AOI22_X1 port map( A1 => n61, A2 => swpOut_0_port, B1 => n138, B2 => 
                           n58, ZN => n154);
   U192 : AOI22_X1 port map( A1 => n58, A2 => n145, B1 => n144, B2 => 
                           cwpOut_0_port, ZN => n158);
   U193 : AOI22_X1 port map( A1 => n35, A2 => swpOut_0_port, B1 => n138, B2 => 
                           n56, ZN => n197);
   U194 : NAND2_X1 port map( A1 => call, A2 => n164, ZN => n162);
   U195 : XNOR2_X1 port map( A => n180, B => n181, ZN => n119);
   U196 : XNOR2_X1 port map( A => n182, B => n183, ZN => n181);
   U197 : OAI22_X1 port map( A1 => n184, A2 => n185, B1 => n36, B2 => n186, ZN 
                           => n180);
   U198 : AOI22_X1 port map( A1 => n80, A2 => n138, B1 => swpOut_3_port, B2 => 
                           n35, ZN => n182);
   U199 : XNOR2_X1 port map( A => n187, B => n188, ZN => n126);
   U200 : XNOR2_X1 port map( A => n189, B => n37, ZN => n188);
   U201 : OAI22_X1 port map( A1 => n190, A2 => n28, B1 => n191, B2 => n192, ZN 
                           => n187);
   U202 : AOI22_X1 port map( A1 => n145, A2 => n80, B1 => oldCWP_3_port, B2 => 
                           n35, ZN => n189);
   U203 : AOI22_X1 port map( A1 => n29, A2 => n138, B1 => swpOut_3_port, B2 => 
                           n61, ZN => n136);
   U204 : OAI211_X1 port map( C1 => n118, C2 => n84, A => n16, B => n177, ZN =>
                           N434);
   U205 : AOI221_X1 port map( B1 => n225, B2 => n38, C1 => need_to_spill_0_port
                           , C2 => n57, A => n145, ZN => n177);
   U206 : NAND4_X1 port map( A1 => ret, A2 => n163, A3 => n117, A4 => n178, ZN 
                           => N433);
   U207 : NOR4_X1 port map( A1 => n53, A2 => N456, A3 => n145, A4 => n100, ZN 
                           => n178);
   U208 : NOR2_X1 port map( A1 => need_to_spill_0_port, A2 => 
                           need_to_fill_0_port, ZN => n101);
   U209 : NAND2_X1 port map( A1 => n163, A2 => n175, ZN => n170);
   U210 : NOR2_X1 port map( A1 => regCnt_0_port, A2 => n112, ZN => N463);
   U211 : NOR2_X1 port map( A1 => n112, A2 => n113, ZN => N466);
   U212 : XNOR2_X1 port map( A => n111, B => regCnt_3_port, ZN => n113);
   U213 : NOR2_X1 port map( A1 => n112, A2 => n116, ZN => N464);
   U214 : XNOR2_X1 port map( A => regCnt_1_port, B => regCnt_0_port, ZN => n116
                           );
   U215 : INV_X1 port map( A => ret, ZN => n85);
   U216 : OR2_X1 port map( A1 => n85, A2 => call, ZN => n179);
   U217 : OAI21_X1 port map( B1 => n104, B2 => n68, A => n208, ZN => N424);
   U218 : NOR2_X1 port map( A1 => n55, A2 => MMUStrobe, ZN => n171);
   U219 : INV_X1 port map( A => need_to_spill_0_port, ZN => n18);
   U220 : NAND2_X1 port map( A1 => n207, A2 => n45, ZN => n167);
   U221 : OAI21_X1 port map( B1 => n75, B2 => n85, A => need_to_fill_0_port, ZN
                           => n207);
   U222 : NAND4_X1 port map( A1 => n172, A2 => n42, A3 => n173, A4 => n174, ZN 
                           => N435);
   U223 : AOI221_X1 port map( B1 => n74, B2 => n170, C1 => n226, C2 => n38, A 
                           => n137, ZN => n174);
   U224 : NAND2_X1 port map( A1 => MMUStrobe, A2 => n168, ZN => n102);
   U225 : OAI21_X1 port map( B1 => n211, B2 => n69, A => n67, ZN => N418);
   U226 : INV_X1 port map( A => N426, ZN => n67);
   U227 : AOI21_X1 port map( B1 => ret, B2 => n164, A => n99, ZN => n211);
   U228 : NAND2_X1 port map( A1 => regCnt_0_port, A2 => n50, ZN => n115);
   U229 : NOR2_X1 port map( A1 => n117, A2 => n2, ZN => N455);
   U230 : INV_X1 port map( A => cwpOut_3_port, ZN => n2);
   U231 : NOR2_X1 port map( A1 => n117, A2 => n25, ZN => N453);
   U232 : INV_X1 port map( A => cwpOut_1_port, ZN => n25);
   U233 : NOR2_X1 port map( A1 => n117, A2 => n20, ZN => N452);
   U234 : INV_X1 port map( A => cwpOut_0_port, ZN => n20);
   U235 : INV_X1 port map( A => cwpOut_2_port, ZN => n27);
   U236 : INV_X1 port map( A => reset, ZN => n84);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerFile_TLE.all;

entity registerFile_TLE is

   port( clk, reset, enable, rd1, rd2, wr1 : in std_logic;  add_wr, add_rd1, 
         add_rd2 : in std_logic_vector (4 downto 0);  dataIn : in 
         std_logic_vector (31 downto 0);  dataOut1, dataOut2, RFtoMEM_BUS : out
         std_logic_vector (31 downto 0);  fill, spill : out std_logic;  call, 
         ret : in std_logic;  dataACK : out std_logic;  MMUStrobe : in 
         std_logic);

end registerFile_TLE;

architecture SYN_struct of registerFile_TLE is

   component physical_RF_NData32_NRegs72_NAddr7
      port( CLK, RESET, ENABLE, RD1, RD2, WR, RD_Mem, WR_Mem : in std_logic;  
            ADD_WR, ADD_RD1, ADD_RD2, ADD_SF : in std_logic_vector (6 downto 0)
            ;  DATAIN : in std_logic_vector (31 downto 0);  OUT1, OUT2, 
            RFtoMEM_BUS : out std_logic_vector (31 downto 0));
   end component;
   
   component 
      translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7
      port( clk, reset, enable, rd1, rd2, wr, fill, spill : in std_logic;  
            add_wr, add_rd1, add_rd2, add_SF : in std_logic_vector (4 downto 0)
            ;  cwp : in std_logic_vector (3 downto 0);  add_wr_out, add_rd1_out
            , add_rd2_out, add_SF_out : out std_logic_vector (6 downto 0));
   end component;
   
   component controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5
      port( clk, reset, enable : in std_logic;  cwpOut, swpOut : out 
            std_logic_vector (3 downto 0);  call, ret : in std_logic;  fill, 
            spill, RD_Mem, WR_Mem : out std_logic;  add_SF : out 
            std_logic_vector (4 downto 0);  MMUStrobe : in std_logic;  dataACK 
            : out std_logic);
   end component;
   
   signal fill_port, spill_port, cwp_s_3_port, cwp_s_2_port, cwp_s_1_port, 
      cwp_s_0_port, RD_Mem_s, WR_Mem_s, add_SF_s_4_port, add_SF_s_3_port, 
      add_SF_s_2_port, add_SF_s_1_port, add_SF_s_0_port, add_wr_out_s_6_port, 
      add_wr_out_s_5_port, add_wr_out_s_4_port, add_wr_out_s_3_port, 
      add_wr_out_s_2_port, add_wr_out_s_1_port, add_wr_out_s_0_port, 
      add_rd1_out_s_6_port, add_rd1_out_s_5_port, add_rd1_out_s_4_port, 
      add_rd1_out_s_3_port, add_rd1_out_s_2_port, add_rd1_out_s_1_port, 
      add_rd1_out_s_0_port, add_rd2_out_s_6_port, add_rd2_out_s_5_port, 
      add_rd2_out_s_4_port, add_rd2_out_s_3_port, add_rd2_out_s_2_port, 
      add_rd2_out_s_1_port, add_rd2_out_s_0_port, add_SF_out_6_port, 
      add_SF_out_5_port, add_SF_out_4_port, add_SF_out_3_port, 
      add_SF_out_2_port, add_SF_out_1_port, add_SF_out_0_port, n_1785, n_1786, 
      n_1787, n_1788, n_1789 : std_logic;

begin
   fill <= fill_port;
   spill <= spill_port;
   
   contrU : controlUnit_RF_N8_M8_F4_windowBlocks3_NData32_NAddr_Windowed5 port 
                           map( clk => clk, reset => reset, enable => enable, 
                           cwpOut(3) => cwp_s_3_port, cwpOut(2) => cwp_s_2_port
                           , cwpOut(1) => cwp_s_1_port, cwpOut(0) => 
                           cwp_s_0_port, swpOut(3) => n_1785, swpOut(2) => 
                           n_1786, swpOut(1) => n_1787, swpOut(0) => n_1788, 
                           call => call, ret => ret, fill => fill_port, spill 
                           => spill_port, RD_Mem => RD_Mem_s, WR_Mem => 
                           WR_Mem_s, add_SF(4) => add_SF_s_4_port, add_SF(3) =>
                           add_SF_s_3_port, add_SF(2) => add_SF_s_2_port, 
                           add_SF(1) => add_SF_s_1_port, add_SF(0) => 
                           add_SF_s_0_port, MMUStrobe => MMUStrobe, dataACK => 
                           n_1789);
   translU : 
                           translationUnit_RF_N8_M8_windowBlocks3_F4_NAddr_Windowed5_NAddr_Physical7 
                           port map( clk => clk, reset => reset, enable => 
                           enable, rd1 => rd1, rd2 => rd2, wr => wr1, fill => 
                           fill_port, spill => spill_port, add_wr(4) => 
                           add_wr(4), add_wr(3) => add_wr(3), add_wr(2) => 
                           add_wr(2), add_wr(1) => add_wr(1), add_wr(0) => 
                           add_wr(0), add_rd1(4) => add_rd1(4), add_rd1(3) => 
                           add_rd1(3), add_rd1(2) => add_rd1(2), add_rd1(1) => 
                           add_rd1(1), add_rd1(0) => add_rd1(0), add_rd2(4) => 
                           add_rd2(4), add_rd2(3) => add_rd2(3), add_rd2(2) => 
                           add_rd2(2), add_rd2(1) => add_rd2(1), add_rd2(0) => 
                           add_rd2(0), add_SF(4) => add_SF_s_4_port, add_SF(3) 
                           => add_SF_s_3_port, add_SF(2) => add_SF_s_2_port, 
                           add_SF(1) => add_SF_s_1_port, add_SF(0) => 
                           add_SF_s_0_port, cwp(3) => cwp_s_3_port, cwp(2) => 
                           cwp_s_2_port, cwp(1) => cwp_s_1_port, cwp(0) => 
                           cwp_s_0_port, add_wr_out(6) => add_wr_out_s_6_port, 
                           add_wr_out(5) => add_wr_out_s_5_port, add_wr_out(4) 
                           => add_wr_out_s_4_port, add_wr_out(3) => 
                           add_wr_out_s_3_port, add_wr_out(2) => 
                           add_wr_out_s_2_port, add_wr_out(1) => 
                           add_wr_out_s_1_port, add_wr_out(0) => 
                           add_wr_out_s_0_port, add_rd1_out(6) => 
                           add_rd1_out_s_6_port, add_rd1_out(5) => 
                           add_rd1_out_s_5_port, add_rd1_out(4) => 
                           add_rd1_out_s_4_port, add_rd1_out(3) => 
                           add_rd1_out_s_3_port, add_rd1_out(2) => 
                           add_rd1_out_s_2_port, add_rd1_out(1) => 
                           add_rd1_out_s_1_port, add_rd1_out(0) => 
                           add_rd1_out_s_0_port, add_rd2_out(6) => 
                           add_rd2_out_s_6_port, add_rd2_out(5) => 
                           add_rd2_out_s_5_port, add_rd2_out(4) => 
                           add_rd2_out_s_4_port, add_rd2_out(3) => 
                           add_rd2_out_s_3_port, add_rd2_out(2) => 
                           add_rd2_out_s_2_port, add_rd2_out(1) => 
                           add_rd2_out_s_1_port, add_rd2_out(0) => 
                           add_rd2_out_s_0_port, add_SF_out(6) => 
                           add_SF_out_6_port, add_SF_out(5) => 
                           add_SF_out_5_port, add_SF_out(4) => 
                           add_SF_out_4_port, add_SF_out(3) => 
                           add_SF_out_3_port, add_SF_out(2) => 
                           add_SF_out_2_port, add_SF_out(1) => 
                           add_SF_out_1_port, add_SF_out(0) => 
                           add_SF_out_0_port);
   physRF : physical_RF_NData32_NRegs72_NAddr7 port map( CLK => clk, RESET => 
                           reset, ENABLE => enable, RD1 => rd1, RD2 => rd2, WR 
                           => wr1, RD_Mem => RD_Mem_s, WR_Mem => WR_Mem_s, 
                           ADD_WR(6) => add_wr_out_s_6_port, ADD_WR(5) => 
                           add_wr_out_s_5_port, ADD_WR(4) => 
                           add_wr_out_s_4_port, ADD_WR(3) => 
                           add_wr_out_s_3_port, ADD_WR(2) => 
                           add_wr_out_s_2_port, ADD_WR(1) => 
                           add_wr_out_s_1_port, ADD_WR(0) => 
                           add_wr_out_s_0_port, ADD_RD1(6) => 
                           add_rd1_out_s_6_port, ADD_RD1(5) => 
                           add_rd1_out_s_5_port, ADD_RD1(4) => 
                           add_rd1_out_s_4_port, ADD_RD1(3) => 
                           add_rd1_out_s_3_port, ADD_RD1(2) => 
                           add_rd1_out_s_2_port, ADD_RD1(1) => 
                           add_rd1_out_s_1_port, ADD_RD1(0) => 
                           add_rd1_out_s_0_port, ADD_RD2(6) => 
                           add_rd2_out_s_6_port, ADD_RD2(5) => 
                           add_rd2_out_s_5_port, ADD_RD2(4) => 
                           add_rd2_out_s_4_port, ADD_RD2(3) => 
                           add_rd2_out_s_3_port, ADD_RD2(2) => 
                           add_rd2_out_s_2_port, ADD_RD2(1) => 
                           add_rd2_out_s_1_port, ADD_RD2(0) => 
                           add_rd2_out_s_0_port, ADD_SF(6) => add_SF_out_6_port
                           , ADD_SF(5) => add_SF_out_5_port, ADD_SF(4) => 
                           add_SF_out_4_port, ADD_SF(3) => add_SF_out_3_port, 
                           ADD_SF(2) => add_SF_out_2_port, ADD_SF(1) => 
                           add_SF_out_1_port, ADD_SF(0) => add_SF_out_0_port, 
                           DATAIN(31) => dataIn(31), DATAIN(30) => dataIn(30), 
                           DATAIN(29) => dataIn(29), DATAIN(28) => dataIn(28), 
                           DATAIN(27) => dataIn(27), DATAIN(26) => dataIn(26), 
                           DATAIN(25) => dataIn(25), DATAIN(24) => dataIn(24), 
                           DATAIN(23) => dataIn(23), DATAIN(22) => dataIn(22), 
                           DATAIN(21) => dataIn(21), DATAIN(20) => dataIn(20), 
                           DATAIN(19) => dataIn(19), DATAIN(18) => dataIn(18), 
                           DATAIN(17) => dataIn(17), DATAIN(16) => dataIn(16), 
                           DATAIN(15) => dataIn(15), DATAIN(14) => dataIn(14), 
                           DATAIN(13) => dataIn(13), DATAIN(12) => dataIn(12), 
                           DATAIN(11) => dataIn(11), DATAIN(10) => dataIn(10), 
                           DATAIN(9) => dataIn(9), DATAIN(8) => dataIn(8), 
                           DATAIN(7) => dataIn(7), DATAIN(6) => dataIn(6), 
                           DATAIN(5) => dataIn(5), DATAIN(4) => dataIn(4), 
                           DATAIN(3) => dataIn(3), DATAIN(2) => dataIn(2), 
                           DATAIN(1) => dataIn(1), DATAIN(0) => dataIn(0), 
                           OUT1(31) => dataOut1(31), OUT1(30) => dataOut1(30), 
                           OUT1(29) => dataOut1(29), OUT1(28) => dataOut1(28), 
                           OUT1(27) => dataOut1(27), OUT1(26) => dataOut1(26), 
                           OUT1(25) => dataOut1(25), OUT1(24) => dataOut1(24), 
                           OUT1(23) => dataOut1(23), OUT1(22) => dataOut1(22), 
                           OUT1(21) => dataOut1(21), OUT1(20) => dataOut1(20), 
                           OUT1(19) => dataOut1(19), OUT1(18) => dataOut1(18), 
                           OUT1(17) => dataOut1(17), OUT1(16) => dataOut1(16), 
                           OUT1(15) => dataOut1(15), OUT1(14) => dataOut1(14), 
                           OUT1(13) => dataOut1(13), OUT1(12) => dataOut1(12), 
                           OUT1(11) => dataOut1(11), OUT1(10) => dataOut1(10), 
                           OUT1(9) => dataOut1(9), OUT1(8) => dataOut1(8), 
                           OUT1(7) => dataOut1(7), OUT1(6) => dataOut1(6), 
                           OUT1(5) => dataOut1(5), OUT1(4) => dataOut1(4), 
                           OUT1(3) => dataOut1(3), OUT1(2) => dataOut1(2), 
                           OUT1(1) => dataOut1(1), OUT1(0) => dataOut1(0), 
                           OUT2(31) => dataOut2(31), OUT2(30) => dataOut2(30), 
                           OUT2(29) => dataOut2(29), OUT2(28) => dataOut2(28), 
                           OUT2(27) => dataOut2(27), OUT2(26) => dataOut2(26), 
                           OUT2(25) => dataOut2(25), OUT2(24) => dataOut2(24), 
                           OUT2(23) => dataOut2(23), OUT2(22) => dataOut2(22), 
                           OUT2(21) => dataOut2(21), OUT2(20) => dataOut2(20), 
                           OUT2(19) => dataOut2(19), OUT2(18) => dataOut2(18), 
                           OUT2(17) => dataOut2(17), OUT2(16) => dataOut2(16), 
                           OUT2(15) => dataOut2(15), OUT2(14) => dataOut2(14), 
                           OUT2(13) => dataOut2(13), OUT2(12) => dataOut2(12), 
                           OUT2(11) => dataOut2(11), OUT2(10) => dataOut2(10), 
                           OUT2(9) => dataOut2(9), OUT2(8) => dataOut2(8), 
                           OUT2(7) => dataOut2(7), OUT2(6) => dataOut2(6), 
                           OUT2(5) => dataOut2(5), OUT2(4) => dataOut2(4), 
                           OUT2(3) => dataOut2(3), OUT2(2) => dataOut2(2), 
                           OUT2(1) => dataOut2(1), OUT2(0) => dataOut2(0), 
                           RFtoMEM_BUS(31) => RFtoMEM_BUS(31), RFtoMEM_BUS(30) 
                           => RFtoMEM_BUS(30), RFtoMEM_BUS(29) => 
                           RFtoMEM_BUS(29), RFtoMEM_BUS(28) => RFtoMEM_BUS(28),
                           RFtoMEM_BUS(27) => RFtoMEM_BUS(27), RFtoMEM_BUS(26) 
                           => RFtoMEM_BUS(26), RFtoMEM_BUS(25) => 
                           RFtoMEM_BUS(25), RFtoMEM_BUS(24) => RFtoMEM_BUS(24),
                           RFtoMEM_BUS(23) => RFtoMEM_BUS(23), RFtoMEM_BUS(22) 
                           => RFtoMEM_BUS(22), RFtoMEM_BUS(21) => 
                           RFtoMEM_BUS(21), RFtoMEM_BUS(20) => RFtoMEM_BUS(20),
                           RFtoMEM_BUS(19) => RFtoMEM_BUS(19), RFtoMEM_BUS(18) 
                           => RFtoMEM_BUS(18), RFtoMEM_BUS(17) => 
                           RFtoMEM_BUS(17), RFtoMEM_BUS(16) => RFtoMEM_BUS(16),
                           RFtoMEM_BUS(15) => RFtoMEM_BUS(15), RFtoMEM_BUS(14) 
                           => RFtoMEM_BUS(14), RFtoMEM_BUS(13) => 
                           RFtoMEM_BUS(13), RFtoMEM_BUS(12) => RFtoMEM_BUS(12),
                           RFtoMEM_BUS(11) => RFtoMEM_BUS(11), RFtoMEM_BUS(10) 
                           => RFtoMEM_BUS(10), RFtoMEM_BUS(9) => RFtoMEM_BUS(9)
                           , RFtoMEM_BUS(8) => RFtoMEM_BUS(8), RFtoMEM_BUS(7) 
                           => RFtoMEM_BUS(7), RFtoMEM_BUS(6) => RFtoMEM_BUS(6),
                           RFtoMEM_BUS(5) => RFtoMEM_BUS(5), RFtoMEM_BUS(4) => 
                           RFtoMEM_BUS(4), RFtoMEM_BUS(3) => RFtoMEM_BUS(3), 
                           RFtoMEM_BUS(2) => RFtoMEM_BUS(2), RFtoMEM_BUS(1) => 
                           RFtoMEM_BUS(1), RFtoMEM_BUS(0) => RFtoMEM_BUS(0));
   dataACK <= '0';

end SYN_struct;
