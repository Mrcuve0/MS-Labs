
package constants is

  constant numBitData : integer := 64;
--  constant numRegs    : integer := 32;

  constant numM : integer;    -- Constant for the number of global registers
  constant numN : integer;    -- Constant for the number of registers in each window 
  constant numF : integer:    -- Constant for the number of windows

end package constants;
