package constants is
  
  constant radixN : integer := 4;
  constant numBit : integer := 32;

end package constants;
